* NGSPICE file created from tt_um_ohmy90_flat_adders.ext - technology: sky130A

.subckt tt_um_ohmy90_flat_adders clk ena rst_n ua[0] ua[1] VPWR Y ua[4] ua[5] ua[6]
+ ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0]
+ uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0]
+ uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0]
+ uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0]
+ uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7] VGND
X0 a_4183_1787# a_4129_2043# a_3790_1761# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X1 a_15255_4841# a_14325_4589# a_15672_4585# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X2 a_24234_14385# ui_in[1] a_24152_14385# VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.10855 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X3 VGND a_14888_5433# a_14836_5459# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X4 a_15113_5825# VPWR a_15017_5825# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X5 a_13732_1769# VGND VPWR w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X6 a_4711_15373# VGND a_4625_15373# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X7 a_11202_5441# a_10611_5471# a_11427_5467# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X8 VPWR VGND a_2313_1791# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X9 VGND a_5636_5017# a_5584_5043# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X10 a_9865_15329# a_9587_15357# VPWR w_9490_15543# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X11 a_1950_5025# Y a_2175_5051# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X12 VPWR VPWR a_15644_5459# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X13 a_5999_1783# a_5873_1757# VPWR w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X14 VPWR VPWR a_9587_15357# w_9490_15543# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X15 a_4513_14775# VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X16 a_6129_12927# a_4913_13781# a_6057_12927# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=1764,126
X17 VPWR VPWR a_6392_5043# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X18 a_11623_4959# a_11569_4849# a_11230_4567# VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X19 VPWR VPWR a_11595_5467# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X20 A a_17125_4938# VPWR sky130_fd_sc_hd__mux2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=6334,279 d=10400,504
X21 a_13802_4955# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X22 a_7113_13395# a_6862_13645# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4010,197 d=6760,364
X23 VPWR VGND a_15239_1765# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X24 a_3820_5021# a_3229_5051# a_4045_5413# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X25 VPWR VGND a_4587_13107# w_4432_13071# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X26 a_13439_4955# a_13313_4563# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X27 a_15045_4951# a_14946_4905# a_14946_4905# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.07384 ps=0.80236 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X28 a_2175_5417# VPWR a_2079_5417# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X29 a_6089_11935# a_4849_11293# a_6003_11935# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X30 VPWR VGND a_4597_11543# w_4442_11507# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X31 VPWR a_9867_12097# a_10965_11919# w_10868_12105# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X32 a_14946_4905# a_14946_4905# a_15309_4951# VNB sky130_fd_pr__nfet_01v8 ad=0.07384 pd=0.80236 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X33 a_17346_5265# sky130_fd_sc_hd__mux2_1_0.A1 a_17125_4938# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
**devattr s=3990,179 d=2772,150
X34 VGND VGND a_9467_13091# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X35 a_15936_2131# VPWR a_15185_2021# VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X36 VGND VPWR a_4213_5413# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X37 a_9671_5727# VGND a_10088_5471# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X38 a_11553_1773# a_11499_2029# a_11160_1747# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X39 a_13774_5463# VGND VPWR w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X40 a_3949_5047# VGND VPWR w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X41 VGND VGND a_8566_2145# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X42 a_9715_16323# VGND VPWR w_9392_16287# sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X43 a_9725_14509# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X44 VGND a_1920_1765# a_1868_1791# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X45 VPWR a_12075_13379# a_12881_13987# w_12566_13951# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=5930,268
X46 a_10422_5837# VPWR a_9671_5727# VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X47 VPWR sky130_fd_sc_hd__inv_1_2.A sky130_fd_sc_hd__inv_1_2.Y sky130_fd_sc_hd__inv_1_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X48 VPWR VPWR a_4753_16339# w_4430_16303# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X49 a_9332_5445# VGND a_9557_5837# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X50 VPWR a_5606_1757# a_5554_1783# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X51 VPWR a_12976_1743# a_12924_1769# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X52 a_4880_1787# VPWR a_4129_2043# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X53 a_5945_2039# a_5873_1757# a_6362_2149# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X54 a_12509_4593# a_11569_4849# VPWR w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X55 a_11359_4959# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X56 VGND VPWR a_4546_2153# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X57 a_4903_15345# a_4625_15373# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X58 a_11541_5723# a_10611_5471# a_11958_5833# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X59 a_11230_4567# a_10639_4597# a_11455_4593# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X60 a_15644_5825# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X61 a_7476_1753# a_6885_1783# a_7701_2145# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X62 VPWR VPWR a_4763_14775# w_4440_14739# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X63 a_11291_12911# a_10937_12911# VPWR w_10872_13125# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5689,267 d=10400,504
X64 a_8232_2145# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X65 a_7869_1779# a_7815_2035# a_7476_1753# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X66 a_5831_2149# VPWR a_5735_2149# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X67 a_4913_13781# a_4635_13809# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X68 a_10813_13753# a_9799_16073# VPWR w_10748_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X69 a_5735_1783# VGND VPWR w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X70 VGND VPWR a_9725_5837# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X71 VPWR a_11202_5441# a_11150_5467# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X72 a_11499_2029# a_10569_1777# a_11916_2139# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X73 a_11986_4593# VGND VPWR w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X74 VPWR VPWR a_9727_11527# w_9404_11491# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X75 a_9753_4597# VPWR VPWR w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X76 a_4723_10577# VGND a_4637_10577# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X77 VPWR VPWR a_11623_4593# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X78 a_4587_13107# VPWR a_4505_13107# w_4432_13071# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X79 a_2079_5051# VGND VPWR w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X80 VGND a_9360_4571# a_9308_4597# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X81 VPWR VPWR a_9599_10561# w_9502_10747# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X82 a_11331_5467# VGND VPWR w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X83 a_4597_11543# VPWR a_4515_11543# w_4442_11507# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X84 a_6944_13645# a_6329_12927# a_6862_13645# w_6756_13609# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X85 a_7669_14003# a_7173_15235# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X86 a_9467_13091# VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X87 sky130_fd_sc_hd__mux2_1_0.A1 a_15255_4841# a_14946_4905# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11427 ps=1.24175 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X88 VPWR VGND a_11595_5467# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X89 a_4635_13809# VGND VPWR w_4538_13995# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X90 a_2706_5417# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X91 VPWR VGND a_2343_5051# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X92 a_15281_5459# a_14297_5463# VPWR w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X93 VGND a_4513_14775# a_4847_14525# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X94 a_5975_5299# a_5903_5017# a_6392_5409# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X95 VGND a_4503_16339# a_4837_16089# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X96 VGND a_9475_14759# a_9809_14509# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X97 a_13315_2025# a_13243_1743# a_13732_2135# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X98 VGND VPWR a_4576_5413# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X99 VGND VGND a_10422_5837# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X100 a_6029_5043# a_5975_5299# a_5636_5017# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X101 a_12135_15219# a_11597_15219# VPWR w_11532_15433# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X102 a_15602_2131# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X103 VPWR VGND a_4880_1787# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X104 VGND sky130_fd_sc_hd__mux2_1_0.S a_16871_4938# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=5796,222
X105 a_11385_1773# VPWR a_11289_1773# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X106 VGND sky130_fd_sc_hd__inv_1_2.A a_23511_14335# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X107 VGND VGND a_4213_5413# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X108 VPWR VGND a_14136_4589# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X109 VGND VGND a_15978_5825# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X110 a_6805_15235# a_4847_14525# a_6717_15235# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X111 a_7899_5405# a_6915_5043# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X112 VPWR VPWR a_13411_5463# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X113 a_15239_2131# a_14255_1769# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X114 a_9727_11527# VGND VPWR w_9404_11491# sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X115 a_1920_1765# sky130_fd_sc_hd__inv_1_0.Y a_2145_2157# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X116 a_14325_4589# a_13385_4845# VPWR w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X117 VPWR a_11230_4567# a_11178_4593# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X118 VGND VPWR a_9753_4963# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X119 sky130_fd_sc_hd__inv_1_4.A sky130_fd_sc_hd__inv_1_5.Y VPWR sky130_fd_sc_hd__inv_1_3.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X120 a_4546_1787# VGND VPWR w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X121 a_23677_14701# ui_in[1] ui_in[0] sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.36 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=4316,272
X122 a_4905_12113# a_4627_12141# VPWR w_4530_12327# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X123 a_4915_10549# a_4637_10577# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X124 a_9461_5837# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X125 a_14888_5433# a_14297_5463# a_15113_5825# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X126 a_7815_2035# a_6885_1783# a_8232_1779# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X127 a_7605_2145# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X128 VPWR a_9809_14509# a_11597_15219# w_11532_15433# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X129 a_6087_14735# a_5809_14763# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X130 VGND a_6281_11907# a_7669_14003# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2772,150 d=2268,138
X131 VGND VPWR a_2313_2157# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X132 VGND VPWR a_11958_5833# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X133 a_13243_5829# VPWR a_13147_5829# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X134 a_9683_2143# a_9629_2033# a_9290_1751# VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X135 VGND VGND a_9725_5837# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X136 a_15672_4585# a_14946_4905# VPWR w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X137 a_13411_5463# a_13357_5719# a_13018_5437# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X138 VPWR VGND a_3010_1791# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X139 a_4183_2153# a_3199_1791# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X140 a_5099_5047# a_4159_5303# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X141 a_11553_2139# a_10569_1777# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X142 VPWR VGND a_11623_4593# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X143 a_4763_14525# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X144 a_15309_4585# a_14325_4589# VPWR w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X145 a_24962_14701# ui_in[0] a_24234_14385# VNB sky130_fd_pr__nfet_01v8 ad=0.15102 pd=1.285 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=6041,257
X146 a_4045_5047# VPWR a_3949_5047# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X147 a_2259_2047# sky130_fd_sc_hd__inv_1_0.Y a_2676_1791# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X148 VPWR VGND a_13369_1769# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X149 a_6696_1783# VPWR a_5945_2039# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X150 VPWR a_9290_1751# a_9238_1777# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X151 a_1950_5025# Y a_2175_5417# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X152 a_12631_13987# a_9877_10533# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=4368,272 d=2772,150
X153 a_9589_12125# VGND VPWR w_9492_12311# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X154 a_11906_13629# a_11291_12911# a_11824_13629# w_11718_13593# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X155 VGND VPWR a_6392_5409# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X156 sky130_fd_sc_hd__inv_1_0.A a_15185_2021# VPWR w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X157 a_9753_4597# a_9699_4853# a_9360_4571# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X158 VPWR a_13018_5437# a_12966_5463# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X159 VGND VPWR a_13732_2135# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X160 a_6915_5043# a_5975_5299# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X161 a_7635_5405# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X162 a_12292_5467# VPWR a_11541_5723# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X163 a_14946_4905# a_14946_4905# a_16006_4951# VNB sky130_fd_pr__nfet_01v8 ad=0.07384 pd=0.80236 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X164 a_14975_2131# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X165 a_15185_2021# a_14255_1769# a_15602_1765# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X166 VPWR VGND a_9547_16323# w_9392_16287# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X167 a_3040_5051# VPWR a_2289_5307# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X168 a_13201_1769# VPWR a_13105_1769# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X169 a_8755_1779# a_7815_2035# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X170 a_5895_14763# a_4849_11293# a_5809_14763# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X171 VGND VGND a_9475_14759# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X172 VGND VGND a_7899_5405# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X173 VPWR a_3790_1761# a_3738_1787# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X174 VGND VPWR a_4711_15373# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X175 VPWR a_9801_12841# a_10771_14747# w_10674_14933# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X176 a_5861_5043# VPWR a_5765_5043# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X177 a_13147_5463# VGND VPWR w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X178 VPWR a_9799_16073# a_11597_15219# w_11532_15433# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X179 a_14916_4559# a_14325_4589# a_15141_4951# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X180 a_5069_1787# a_4129_2043# VPWR w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X181 a_10639_4597# a_9699_4853# VPWR w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X182 VGND VPWR a_2676_2157# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X183 a_13271_4955# VPWR a_13175_4955# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X184 VGND VGND a_4513_14775# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X185 a_9671_5727# VGND a_10088_5837# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X186 VPWR a_14916_4559# a_14864_4585# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X187 a_11051_11919# a_9811_11277# a_10965_11919# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X188 a_13774_5829# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X189 a_3790_1761# a_3199_1791# a_4015_1787# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X190 VPWR VPWR a_13802_4589# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X191 VPWR VPWR a_8232_1779# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X192 a_11351_13753# a_10813_13753# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X193 VGND VGND a_2313_2157# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X194 VPWR a_11351_13753# a_11906_13629# w_11718_13593# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5830,267
X195 a_9515_2143# VPWR a_9419_2143# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X196 ua[0] a_24962_14701# VPWR sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X197 a_4755_13107# VGND VPWR w_4432_13071# sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X198 VPWR VGND a_6696_1783# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X199 a_5999_2149# a_5873_1757# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X200 VPWR VPWR a_4183_1787# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X201 a_5933_13769# a_4849_11293# a_5851_13769# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
X202 a_9673_15357# VGND a_9587_15357# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X203 a_4576_5047# VGND VPWR w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X204 VGND VGND a_15281_5825# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X205 VGND a_11160_1747# a_11108_1773# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X206 a_11230_4567# a_10639_4597# a_11455_4959# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X207 a_11597_15219# a_8113_13753# VPWR w_11532_15433# sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X208 a_4765_11543# VGND VPWR w_4442_11507# sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X209 a_6885_1783# a_5945_2039# VPWR w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X210 a_9683_13793# VGND a_9597_13793# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X211 VPWR VGND a_12292_5467# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X212 a_9547_16323# VPWR a_9465_16323# w_9392_16287# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X213 a_4503_16339# VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X214 a_5606_1757# a_5873_1757# a_5831_1783# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X215 a_11986_4959# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X216 a_9475_14759# VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X217 a_4015_2153# VPWR a_3919_2153# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X218 a_17339_4938# sky130_fd_sc_hd__mux2_1_0.A0 a_17125_4938# sky130_fd_sc_hd__mux2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
**devattr s=7728,268 d=3066,157
X219 VPWR VGND a_3040_5051# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X220 a_11595_5833# a_11541_5723# a_11202_5441# VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X221 a_6362_1783# VGND VPWR w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X222 a_12320_4593# VPWR a_11569_4849# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X223 VGND VPWR a_11623_4959# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X224 VPWR VPWR a_9715_16323# w_9392_16287# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X225 a_10771_14747# a_9811_11277# VPWR w_10674_14933# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X226 a_9809_14509# VPWR a_9725_14509# VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X227 a_2079_5417# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X228 a_3229_5051# a_2289_5307# VPWR w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X229 a_9629_2033# a_8755_1779# a_10046_1777# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X230 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X231 a_12481_5467# a_11541_5723# VPWR w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X232 a_12439_1773# a_11499_2029# VPWR w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X233 a_15309_4585# a_15255_4841# a_14916_4559# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X234 a_9585_4597# VPWR a_9489_4597# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X235 a_11553_2139# a_11499_2029# a_11160_1747# VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X236 a_11160_1747# a_10569_1777# a_11385_1773# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X237 a_14066_1769# VPWR a_13315_2025# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X238 VGND a_7476_1753# a_7424_1779# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X239 a_2289_5307# Y a_2706_5051# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X240 a_15978_5459# VPWR a_15227_5715# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X241 ui_in[0] a_23731_14309# a_23677_14335# VNB sky130_fd_pr__nfet_01v8 ad=0.09322 pd=1.07 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3409,185
X242 a_6389_13769# a_5851_13769# VPWR w_5786_13983# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X243 a_11958_5467# VGND VPWR w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X244 VPWR a_4903_15345# a_5851_13769# w_5786_13983# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X245 VGND VGND a_2343_5417# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X246 VPWR VPWR a_15602_1765# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X247 a_7751_14003# a_4915_10549# a_7669_14003# w_7604_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2772,150
X248 VPWR VGND a_9559_11527# w_9404_11491# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X249 sky130_fd_sc_hd__mux2_1_0.A0 a_15227_5715# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X250 VPWR VPWR a_2343_5051# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X251 a_9683_1777# a_8755_1779# VPWR w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X252 a_9699_4853# VPWR a_10116_4963# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X253 VGND VPWR a_4723_10577# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X254 a_13369_2135# a_13243_1743# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X255 a_4625_15373# VGND VPWR w_4528_15559# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X256 a_14136_4955# VPWR a_13385_4845# VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X257 a_11049_14719# a_10771_14747# VPWR w_10674_14933# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X258 a_4159_5303# a_3229_5051# a_4576_5413# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X259 a_6029_5409# a_5975_5299# a_5636_5017# VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X260 a_14946_4905# VPWR a_15672_4951# VNB sky130_fd_pr__nfet_01v8 ad=0.07384 pd=0.80236 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X261 a_8596_5405# VPWR a_7845_5295# VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X262 a_5735_2149# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X263 a_24774_14701# ui_in[0] VPWR sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X264 VPWR a_3820_5021# a_3768_5047# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X265 a_9865_15329# a_9587_15357# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X266 VPWR VPWR a_4635_13809# w_4538_13995# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X267 VGND VPWR a_13411_5829# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X268 a_14108_5463# VPWR a_13357_5719# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X269 a_9875_13765# a_9597_13793# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X270 a_10569_1777# a_9629_2033# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X271 VPWR VGND a_4183_1787# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X272 a_17125_4938# sky130_fd_sc_hd__mux2_1_0.A1 a_17053_4938# sky130_fd_sc_hd__mux2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=7728,268
X273 VPWR VGND a_12320_4593# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X274 a_11291_12911# a_10937_12911# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=5266,228 d=6760,364
X275 VGND a_7506_5013# a_7454_5039# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X276 VPWR sky130_fd_sc_hd__inv_1_2.A a_23511_14701# sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X277 a_8113_13753# a_7669_14003# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4075,198 d=7020,368
X278 VGND a_14846_1739# a_14794_1765# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X279 a_15071_2131# VPWR a_14975_2131# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X280 VPWR sky130_fd_sc_hd__inv_1_0.A sky130_fd_sc_hd__inv_1_0.Y sky130_fd_sc_hd__inv_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X281 VGND a_13046_4563# a_12994_4589# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X282 ui_in[0] a_24774_14701# a_24962_14701# VNB sky130_fd_pr__nfet_01v8 ad=0.09322 pd=1.07 as=0.15102 ps=1.285 w=0.42 l=0.15
**devattr s=6041,257 d=4368,272
X283 a_6057_12927# a_4849_11293# a_5975_12927# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X284 a_9725_5471# VGND VPWR w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X285 a_7869_1779# a_6885_1783# VPWR w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X286 a_3199_1791# a_2259_2047# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X287 VPWR VPWR a_8262_5039# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X288 a_23677_14335# sky130_fd_sc_hd__inv_1_5.Y VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X289 VPWR VGND a_14066_1769# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X290 a_13411_5829# a_13357_5719# a_13018_5437# VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X291 VGND a_6389_13769# a_6862_13645# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4010,197
X292 a_9559_11527# VPWR a_9477_11527# w_9404_11491# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X293 a_11427_5833# VPWR a_11331_5833# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X294 a_16006_4585# VPWR a_15255_4841# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X295 VGND VGND a_11623_4959# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X296 a_7919_14003# a_7173_15235# a_7847_14003# w_7604_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X297 a_14255_1769# a_13315_2025# VPWR w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X298 a_11243_11891# a_10965_11919# VPWR w_10868_12105# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X299 VPWR VPWR a_10046_1777# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X300 a_12976_1743# a_13243_1743# a_13201_1769# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X301 a_2313_1791# sky130_fd_sc_hd__inv_1_0.Y VPWR w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X302 a_5975_12927# a_4913_13781# VPWR w_5910_13141# sky130_fd_pr__pfet_01v8_hvt ad=0.0805 pd=0.94333 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2646,147
X303 a_11385_2139# VPWR a_11289_2139# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X304 VPWR VPWR a_2706_5051# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X305 a_11289_1773# VGND VPWR w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X306 a_4213_5047# a_4159_5303# a_3820_5021# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X307 a_5636_5017# a_5903_5017# a_5861_5043# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X308 VPWR VPWR a_5999_1783# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X309 VPWR VPWR a_13369_1769# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X310 a_15141_4585# VPWR a_15045_4585# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X311 VGND VGND a_8596_5405# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X312 a_6392_5043# VGND VPWR w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X313 VGND a_4837_16089# a_6911_15235# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X314 VGND VGND a_15936_2131# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X315 VGND VPWR a_10116_4963# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X316 a_13046_4563# a_13313_4563# a_13271_4955# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X317 VPWR VGND a_11553_1773# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X318 VPWR VGND a_14108_5463# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X319 a_4847_14525# VPWR a_4763_14525# VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X320 a_6029_5043# a_5903_5017# VPWR w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X321 VGND VPWR a_13439_4955# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X322 a_3040_5417# VPWR a_2289_5307# VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X323 a_7506_5013# a_6915_5043# a_7731_5405# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X324 a_8262_5405# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X325 a_10380_2143# VPWR a_9629_2033# VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X326 a_13147_5829# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X327 a_9290_1751# a_8755_1779# a_9515_2143# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X328 a_4713_12141# VGND a_4627_12141# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X329 a_5861_5409# VPWR a_5765_5409# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X330 a_14297_5463# a_13357_5719# VPWR w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X331 a_10983_13753# a_9865_15329# a_10895_13753# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X332 a_11089_13753# a_9799_16073# a_10983_13753# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X333 a_13018_5437# a_13285_5437# a_13243_5463# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X334 a_13369_2135# a_13315_2025# a_12976_1743# VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X335 VGND VGND a_3010_2157# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X336 a_9867_12097# a_9589_12125# VPWR w_9492_12311# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X337 a_6717_15235# sky130_fd_sc_hd__inv_1_2.Y a_6635_15235# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
X338 a_4837_16089# a_4503_16339# a_4753_16339# w_4430_16303# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X339 VPWR VPWR a_9589_12125# w_9492_12311# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X340 VPWR VPWR a_10088_5471# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X341 a_9877_10533# a_9599_10561# VPWR w_9502_10747# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X342 VPWR VGND a_7869_1779# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X343 VGND VPWR a_9683_2143# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X344 a_2259_2047# sky130_fd_sc_hd__inv_1_0.Y a_2676_2157# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X345 a_4753_16089# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X346 VPWR a_4849_11293# a_5975_12927# w_5910_13141# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0805 ps=0.94333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X347 VGND a_4839_12857# a_5895_14763# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X348 a_6696_2149# VPWR a_5945_2039# VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X349 a_15227_5715# a_14297_5463# a_15644_5825# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X350 a_10450_4597# VPWR a_9699_4853# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X351 VPWR a_14888_5433# a_14836_5459# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X352 a_9360_4571# VPWR a_9585_4597# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X353 sky130_fd_sc_hd__inv_1_5.Y sky130_fd_sc_hd__inv_1_5.A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X354 VPWR a_5636_5017# a_5584_5043# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X355 a_7701_1779# VPWR a_7605_1779# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X356 a_12135_15219# a_11597_15219# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X357 a_4910_5047# VPWR a_4159_5303# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X358 a_13439_4589# a_13385_4845# a_13046_4563# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X359 a_11569_4849# a_10639_4597# a_11986_4593# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X360 VGND a_9867_12097# a_11051_11919# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X361 a_13105_1769# VGND VPWR w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X362 VGND VPWR a_7869_2145# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X363 a_17125_4938# sky130_fd_sc_hd__mux2_1_0.A0 a_17125_5265# VNB sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=3990,179
X364 a_15017_5459# VGND VPWR w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X365 VGND sky130_fd_sc_hd__inv_1_2.A sky130_fd_sc_hd__inv_1_2.Y VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X366 VGND VGND a_3040_5417# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X367 VPWR VGND a_5999_1783# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X368 a_7899_5039# a_7845_5295# a_7506_5013# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X369 a_11873_15219# a_11049_14719# a_11767_15219# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X370 VPWR a_9801_12841# a_10813_13753# w_10748_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X371 a_5765_5043# VGND VPWR w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X372 a_12509_4593# a_11569_4849# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X373 a_12320_4959# VPWR a_11569_4849# VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X374 VGND VGND a_10380_2143# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X375 VGND a_4505_13107# a_4839_12857# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X376 VPWR VPWR a_4755_13107# w_4432_13071# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X377 A a_17125_4938# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4514,209 d=6760,364
X378 a_10937_12911# a_9875_13765# VPWR w_10872_13125# sky130_fd_pr__pfet_01v8_hvt ad=0.0805 pd=0.94333 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2646,147
X379 a_11595_5467# a_10611_5471# VPWR w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X380 a_13175_4955# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X381 a_4905_12113# a_4627_12141# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X382 a_2289_5307# Y a_2706_5417# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X383 VPWR VPWR a_15281_5459# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X384 VGND VPWR a_9673_15357# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X385 VPWR A a_24407_14651# sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.09013 ps=0.995 w=0.42 l=0.15
**devattr s=3605,199 d=2268,138
X386 VPWR VPWR a_4765_11543# w_4442_11507# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X387 VPWR a_7113_13395# a_7919_14003# w_7604_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=5930,268
X388 VGND VGND a_13439_4955# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X389 VGND VPWR a_9683_13793# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X390 a_10046_2143# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X391 VGND VGND a_4503_16339# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X392 VGND VPWR a_2343_5417# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X393 a_9419_2143# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X394 a_12075_13379# a_11824_13629# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4010,197 d=6760,364
X395 VGND VGND a_6696_2149# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X396 sky130_fd_sc_hd__inv_1_2.A a_12631_13987# VPWR w_12566_13951# sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5930,268 d=10800,508
X397 a_12250_1773# VPWR a_11499_2029# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X398 a_4213_5413# a_3229_5051# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X399 a_14846_1739# a_14255_1769# a_15071_2131# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X400 VPWR VGND a_10450_4597# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X401 VPWR VPWR a_13774_5463# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X402 a_15239_1765# a_15185_2021# a_14846_1739# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X403 a_15281_5459# a_15227_5715# a_14888_5433# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X404 VGND VPWR a_7899_5405# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X405 VGND VPWR a_15239_2131# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X406 VGND VGND a_9683_2143# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X407 a_15255_4841# a_14325_4589# a_15672_4951# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X408 sky130_fd_sc_hd__inv_1_5.A sky130_fd_sc_hd__inv_1_4.A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X409 a_6862_13645# a_6329_12927# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X410 VPWR VGND a_4910_5047# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X411 VPWR VGND a_13411_5463# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X412 a_5606_1757# a_5873_1757# a_5831_2149# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X413 a_11202_5441# a_10611_5471# a_11427_5833# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X414 a_14108_5829# VPWR a_13357_5719# VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X415 a_6362_2149# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X416 VGND a_5606_1757# a_5554_1783# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X417 a_3919_2153# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X418 a_4129_2043# a_3199_1791# a_4546_1787# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X419 a_5851_13769# a_4849_11293# VPWR w_5786_13983# sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X420 a_4721_13809# VGND a_4635_13809# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X421 VPWR a_9865_15329# a_10813_13753# w_10748_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X422 VPWR a_4847_14525# a_6635_15235# w_6570_15449# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X423 VGND VPWR a_15644_5825# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X424 a_8566_1779# VPWR a_7815_2035# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X425 a_10116_4597# VGND VPWR w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X426 VGND VGND a_12320_4959# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X427 VGND a_9801_12841# a_11089_13753# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X428 a_9489_4597# VGND VPWR w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X429 VPWR VPWR a_4625_15373# w_4528_15559# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X430 a_12631_13987# a_12135_15219# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X431 a_9725_5837# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X432 a_11160_1747# a_10569_1777# a_11385_2139# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X433 a_13385_4845# a_13313_4563# a_13802_4589# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X434 VGND VPWR a_11595_5833# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X435 VPWR VPWR a_11986_4593# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X436 a_7113_13395# a_6862_13645# VPWR w_6756_13609# sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5830,267 d=13600,536
X437 a_11091_12911# a_9875_13765# a_11019_12911# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=1764,126
X438 sky130_fd_sc_hd__mux2_1_0.S a_7845_5295# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X439 a_11623_4593# a_10639_4597# VPWR w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X440 a_7845_5295# a_6915_5043# a_8262_5039# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X441 a_14325_4589# a_13385_4845# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X442 a_9557_5471# VPWR a_9461_5471# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X443 VPWR VPWR a_15309_4585# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X444 VPWR VGND a_9753_4597# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X445 VPWR sky130_fd_sc_hd__mux2_1_0.S a_17339_4938# sky130_fd_sc_hd__mux2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=6334,279
X446 VGND a_11230_4567# a_11178_4593# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X447 a_7731_5039# VPWR a_7635_5039# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X448 a_24774_14701# ui_in[0] VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X449 VPWR VGND a_12250_1773# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X450 a_23677_14701# sky130_fd_sc_hd__inv_1_5.Y VPWR sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.36 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X451 VGND VGND a_4505_13107# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X452 VGND VPWR a_2706_5417# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X453 a_5636_5017# a_5903_5017# a_5861_5409# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X454 a_4183_2153# a_4129_2043# a_3790_1761# VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X455 a_3949_5413# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X456 a_6392_5409# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X457 ua[0] a_24962_14701# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X458 a_9801_12841# a_9467_13091# a_9717_13091# w_9394_13055# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X459 a_13732_2135# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X460 a_2145_1791# VPWR a_2049_1791# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X461 a_6726_5043# VPWR a_5975_5299# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X462 a_15936_1765# VPWR a_15185_2021# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X463 a_5809_14763# a_4849_11293# VPWR w_5712_14949# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X464 a_6029_5409# a_5903_5017# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X465 VGND VGND a_14108_5829# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X466 a_11916_1773# VGND VPWR w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X467 VGND a_9801_12841# a_11091_12911# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5266,228
X468 VPWR VPWR a_11553_1773# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X469 VPWR VGND a_8566_1779# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X470 a_15113_5459# VPWR a_15017_5459# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X471 VGND a_11243_11891# a_12631_13987# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2772,150 d=2268,138
X472 VPWR a_4837_16089# a_6635_15235# w_6570_15449# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X473 VGND VGND a_15239_2131# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X474 a_13018_5437# a_13285_5437# a_13243_5829# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X475 a_8755_1779# a_7815_2035# VPWR w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X476 a_9753_4963# VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X477 VPWR VPWR a_4546_1787# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X478 VGND VPWR a_10088_5837# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X479 a_7476_1753# a_6885_1783# a_7701_1779# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X480 a_13802_4589# VGND VPWR w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X481 a_12713_13987# a_9877_10533# a_12631_13987# w_12566_13951# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2772,150
X482 a_8232_1779# VGND VPWR w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X483 a_10611_5471# a_9671_5727# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X484 a_11331_5833# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X485 a_2313_2157# sky130_fd_sc_hd__inv_1_0.Y VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X486 a_11767_15219# a_9809_14509# a_11679_15219# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X487 a_11824_13629# a_11291_12911# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X488 a_5099_5047# a_4159_5303# VPWR w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X489 a_11289_2139# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X490 VGND a_9332_5445# a_9280_5471# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X491 a_3820_5021# a_3229_5051# a_4045_5047# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X492 VGND VPWR a_5999_2149# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X493 a_10813_13753# a_9811_11277# VPWR w_10748_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X494 a_4505_13107# VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X495 VGND VGND a_11595_5833# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X496 a_13439_4589# a_13313_4563# VPWR w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X497 a_15045_4585# a_14946_4905# VPWR w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X498 a_6635_15235# sky130_fd_sc_hd__inv_1_2.Y VPWR w_6570_15449# sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X499 VGND VPWR a_4713_12141# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X500 a_15281_5825# a_14297_5463# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X501 VGND VGND a_4515_11543# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X502 a_10639_4597# a_9699_4853# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X503 VGND a_9801_12841# a_10857_14747# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X504 VPWR a_14946_4905# a_15309_4585# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X505 a_14946_4905# a_14916_4559# a_14864_4585# VNB sky130_fd_pr__nfet_01v8 ad=0.11427 pd=1.24175 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X506 a_11049_14719# a_10771_14747# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X507 a_9597_13793# VGND VPWR w_9500_13979# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X508 VGND VGND a_11553_2139# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X509 VPWR VPWR a_4213_5047# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X510 VPWR VGND a_6726_5043# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X511 a_4880_2153# VPWR a_4129_2043# VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X512 a_11569_4849# a_10639_4597# a_11986_4959# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X513 a_9715_16073# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X514 a_2676_1791# VGND VPWR w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X515 VPWR a_11160_1747# a_11108_1773# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X516 a_7869_2145# a_7815_2035# a_7476_1753# VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X517 a_5765_5409# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X518 VGND VGND a_14136_4955# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X519 a_4837_16089# VPWR a_4753_16089# VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X520 a_6915_5043# a_5975_5299# VPWR w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X521 a_4913_13781# a_4635_13809# VPWR w_4538_13995# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X522 VPWR a_4839_12857# a_5975_12927# w_5910_13141# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0805 ps=0.94333 w=0.42 l=0.15
**devattr s=2646,147 d=5689,267
X523 a_6329_12927# a_5975_12927# VPWR w_5910_13141# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5689,267 d=10400,504
X524 VGND a_1950_5025# a_1898_5051# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X525 a_13315_2025# a_13243_1743# a_13732_1769# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X526 VPWR a_9811_11277# a_10937_12911# w_10872_13125# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0805 ps=0.94333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X527 VPWR VPWR a_11916_1773# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X528 a_11541_5723# a_10611_5471# a_11958_5467# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X529 a_15644_5459# VGND VPWR w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X530 a_9675_12125# VGND a_9589_12125# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X531 a_15602_1765# VGND VPWR w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X532 a_11597_15219# a_11049_14719# VPWR w_11532_15433# sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X533 a_24234_14385# ui_in[1] a_24241_14651# sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1274 pd=1.16667 as=0.10855 ps=1.36 w=0.42 l=0.15
**devattr s=4316,272 d=2268,138
X534 VPWR VPWR a_9717_13091# w_9394_13055# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X535 a_6281_11907# a_6003_11935# VPWR w_5906_12121# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X536 a_9811_11277# VPWR a_9727_11277# VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X537 VGND a_3790_1761# a_3738_1787# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X538 VPWR a_4905_12113# a_6003_11935# w_5906_12121# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X539 a_9685_10561# VGND a_9599_10561# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X540 a_15239_1765# a_14255_1769# VPWR w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X541 VPWR a_7476_1753# a_7424_1779# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X542 a_4847_14525# a_4513_14775# a_4763_14775# w_4440_14739# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X543 a_5069_1787# a_4129_2043# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X544 a_15672_4951# a_14946_4905# a_14946_4905# VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.07384 ps=0.80236 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X545 a_9809_14509# a_9475_14759# a_9725_14759# w_9402_14723# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X546 a_10895_13753# a_9811_11277# a_10813_13753# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
X547 a_4515_11543# VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X548 VGND VPWR a_13774_5829# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X549 a_10857_14747# a_9811_11277# a_10771_14747# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X550 a_7605_1779# VGND VPWR w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X551 a_7847_14003# a_6281_11907# a_7751_14003# w_7604_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X552 a_15309_4951# a_14325_4589# a_14946_4905# VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.07384 ps=0.80236 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X553 a_13357_5719# a_13285_5437# a_13774_5463# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X554 a_9683_1777# a_9629_2033# a_9290_1751# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X555 a_17125_5265# a_16871_4938# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=5796,222 d=2772,150
X556 a_24241_14651# sky130_fd_sc_hd__inv_1_0.A VPWR sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.36 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X557 a_4045_5413# VPWR a_3949_5413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X558 VGND VGND a_13411_5829# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X559 VGND VGND a_4880_2153# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X560 VGND a_9465_16323# a_9799_16073# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X561 VGND VGND a_5999_2149# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X562 a_4183_1787# a_3199_1791# VPWR w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X563 VPWR VPWR a_4576_5047# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X564 a_6021_13769# a_4903_15345# a_5933_13769# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X565 VPWR a_1920_1765# a_1868_1791# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X566 VGND A a_24152_14385# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.10855 ps=1.36 w=0.42 l=0.15
**devattr s=4316,272 d=2268,138
X567 a_6127_13769# a_4837_16089# a_6021_13769# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X568 a_4627_12141# VGND VPWR w_4530_12327# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X569 a_6885_1783# a_5945_2039# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X570 a_9753_4963# a_9699_4853# a_9360_4571# VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X571 VPWR VGND a_4213_5047# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X572 a_12292_5833# VPWR a_11541_5723# VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X573 a_4546_2153# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X574 VGND VPWR a_11986_4959# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X575 a_4637_10577# VGND VPWR w_4540_10763# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X576 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X577 a_10569_1777# a_9629_2033# VPWR w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X578 a_11623_4959# a_10639_4597# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X579 VPWR VGND a_15978_5459# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X580 a_9717_13091# VGND VPWR w_9394_13055# sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X581 a_9727_11277# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X582 a_7815_2035# a_6885_1783# a_8232_2145# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X583 a_7899_5039# a_6915_5043# VPWR w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X584 VGND ui_in[1] a_23731_14309# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X585 VPWR a_14846_1739# a_14794_1765# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X586 a_6003_11935# a_4849_11293# VPWR w_5906_12121# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X587 a_9557_5837# VPWR a_9461_5837# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X588 VPWR VPWR a_6362_1783# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X589 a_12250_2139# VPWR a_11499_2029# VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X590 VPWR VPWR a_13732_1769# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X591 sky130_fd_sc_hd__inv_1_4.A sky130_fd_sc_hd__inv_1_5.Y VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X592 VGND VPWR a_4721_13809# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X593 a_9725_5471# a_9671_5727# a_9332_5445# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X594 VPWR VPWR a_9753_4597# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X595 a_11455_4593# VPWR a_11359_4593# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X596 sky130_fd_sc_hd__mux2_1_0.A0 a_15227_5715# VPWR w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X597 a_9877_10533# a_9599_10561# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X598 VGND a_11202_5441# a_11150_5467# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X599 a_14975_1765# VGND VPWR w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X600 a_14888_5433# a_14297_5463# a_15113_5459# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X601 VGND a_12075_13379# a_12631_13987# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2268,138 d=4075,198
X602 VPWR a_9801_12841# a_10937_12911# w_10872_13125# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0805 ps=0.94333 w=0.42 l=0.15
**devattr s=2646,147 d=5689,267
X603 VPWR VPWR a_11958_5467# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X604 a_2343_5051# Y VPWR w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X605 VGND VGND a_13369_2135# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X606 VGND VPWR a_13802_4955# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X607 a_7173_15235# a_6635_15235# VPWR w_6570_15449# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X608 a_24234_14385# a_24774_14701# a_24962_14701# sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1274 pd=1.16667 as=0.09209 ps=0.99 w=0.42 l=0.15
**devattr s=3683,198 d=10752,424
X609 a_6726_5409# VPWR a_5975_5299# VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X610 VPWR VPWR a_6029_5043# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X611 a_2313_1791# a_2259_2047# a_1920_1765# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X612 a_12881_13987# a_12135_15219# a_12809_13987# w_12566_13951# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X613 a_4576_5413# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X614 a_4755_12857# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X615 VGND a_4515_11543# a_4849_11293# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X616 VPWR a_7506_5013# a_7454_5039# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X617 a_9515_1777# VPWR a_9419_1777# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X618 VGND a_12976_1743# a_12924_1769# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X619 a_13201_2135# VPWR a_13105_2135# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X620 a_15185_2021# a_14255_1769# a_15602_2131# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X621 VGND VGND a_12292_5833# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X622 a_10088_5471# VGND VPWR w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X623 a_4585_16339# VPWR a_4503_16339# w_4430_16303# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X624 VGND a_9477_11527# a_9811_11277# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X625 VPWR a_14946_4905# a_16006_4585# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X626 VPWR a_4839_12857# a_5809_14763# w_5712_14949# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X627 a_7635_5039# VGND VPWR w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X628 VGND VGND a_9465_16323# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X629 a_4595_14775# VPWR a_4513_14775# w_4440_14739# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X630 VGND VGND a_12250_2139# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X631 VPWR a_9360_4571# a_9308_4597# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X632 a_15309_4951# a_15255_4841# a_14916_4559# VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X633 a_9585_4963# VPWR a_9489_4963# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X634 VPWR VGND a_7899_5039# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X635 a_15978_5825# VPWR a_15227_5715# VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X636 a_3790_1761# a_3199_1791# a_4015_2153# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X637 a_11958_5833# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X638 a_4015_1787# VPWR a_3919_1787# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X639 sky130_fd_sc_hd__mux2_1_0.A1 a_15255_4841# VPWR w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X640 VGND VPWR a_8232_2145# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X641 a_2049_1791# VGND VPWR w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X642 a_2145_2157# VPWR a_2049_2157# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X643 a_14916_4559# a_14325_4589# a_15141_4585# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X644 sky130_fd_sc_hd__inv_1_2.A a_12631_13987# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4075,198 d=7020,368
X645 a_11351_13753# a_10813_13753# VPWR w_10748_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X646 a_11916_2139# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X647 a_13271_4589# VPWR a_13175_4589# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X648 a_6389_13769# a_5851_13769# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X649 a_4839_12857# a_4505_13107# a_4755_13107# w_4432_13071# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X650 VGND VGND a_6726_5409# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X651 VGND VPWR a_4183_2153# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X652 VGND VPWR a_11553_2139# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X653 VGND a_4839_12857# a_6127_13769# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X654 VGND a_11351_13753# a_11824_13629# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4010,197
X655 a_3010_1791# VPWR a_2259_2047# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X656 a_13369_1769# a_13243_1743# VPWR w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X657 a_23511_14335# ui_in[1] ui_in[0] VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.09322 ps=1.07 w=0.42 l=0.15
**devattr s=3409,185 d=4368,272
X658 a_9725_14759# VGND VPWR w_9402_14723# sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X659 a_4765_11293# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X660 VPWR VGND a_6029_5043# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X661 a_5999_1783# a_5945_2039# a_5606_1757# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X662 VPWR VGND a_15281_5459# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X663 VPWR VPWR a_9597_13793# w_9500_13979# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X664 a_4903_15345# a_4625_15373# VPWR w_4528_15559# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X665 a_9629_2033# a_8755_1779# a_10046_2143# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X666 VGND a_9799_16073# a_11873_15219# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X667 a_9465_16323# VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X668 a_14066_2135# VPWR a_13315_2025# VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X669 a_9799_16073# VPWR a_9715_16073# VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X670 VGND VPWR a_8262_5405# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X671 a_11595_5467# a_11541_5723# a_11202_5441# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X672 VGND a_13018_5437# a_12966_5463# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X673 VGND VPWR a_15602_2131# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X674 a_2343_5051# a_2289_5307# a_1950_5025# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X675 a_7669_14003# a_4915_10549# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=4368,272 d=2772,150
X676 a_15071_1765# VPWR a_14975_1765# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X677 a_9683_2143# a_8755_1779# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X678 a_16006_4951# VPWR a_15255_4841# VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X679 VPWR a_6389_13769# a_6944_13645# w_6756_13609# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5830,267
X680 VPWR sky130_fd_sc_hd__mux2_1_0.S a_16871_4938# sky130_fd_sc_hd__mux2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2772,150
X681 a_13411_5463# a_13285_5437# VPWR w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X682 a_13357_5719# a_13285_5437# a_13774_5829# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X683 VPWR VGND a_9549_13091# w_9394_13055# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X684 VGND VPWR a_9675_12125# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X685 VGND VGND a_9477_11527# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X686 a_24407_14651# a_23731_14309# a_24234_14385# sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09013 pd=0.995 as=0.1274 ps=1.16667 w=0.42 l=0.15
**devattr s=2268,138 d=3605,199
X687 VGND a_4839_12857# a_6129_12927# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5266,228
X688 a_2676_2157# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X689 a_11679_15219# a_8113_13753# a_11597_15219# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
X690 VGND VPWR a_9685_10561# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X691 a_4213_5413# a_4159_5303# a_3820_5021# VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X692 a_9699_4853# VPWR a_10116_4597# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X693 a_15141_4951# VPWR a_15045_4951# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X694 a_9587_15357# VGND VPWR w_9490_15543# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X695 a_11019_12911# a_9811_11277# a_10937_12911# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X696 a_11243_11891# a_10965_11919# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X697 VGND VPWR a_11916_2139# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X698 a_14136_4589# VPWR a_13385_4845# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X699 a_4159_5303# a_3229_5051# a_4576_5047# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X700 VPWR VPWR a_15672_4585# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X701 VGND sky130_fd_sc_hd__mux2_1_0.S a_17346_5265# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=4514,209
X702 VGND VGND a_4183_2153# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X703 a_8596_5039# VPWR a_7845_5295# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X704 VGND a_9290_1751# a_9238_1777# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X705 a_9875_13765# a_9597_13793# VPWR w_9500_13979# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X706 a_7869_2145# a_6885_1783# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X707 a_8113_13753# a_7669_14003# VPWR w_7604_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5930,268 d=10800,508
X708 a_6329_12927# a_5975_12927# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=5266,228 d=6760,364
X709 sky130_fd_sc_hd__inv_1_0.A a_15185_2021# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X710 VPWR VGND a_15936_1765# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X711 VGND VGND a_14066_2135# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X712 a_9725_5837# a_9671_5727# a_9332_5445# VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X713 a_5945_2039# a_5873_1757# a_6362_1783# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X714 a_11455_4959# VPWR a_11359_4959# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X715 a_10965_11919# a_9811_11277# VPWR w_10868_12105# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X716 a_24318_14385# sky130_fd_sc_hd__inv_1_0.A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10858 pd=1.36 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X717 a_11623_4593# a_11569_4849# a_11230_4567# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X718 a_9801_12841# VPWR a_9717_12841# VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X719 VPWR VPWR a_4627_12141# w_4530_12327# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X720 a_6281_11907# a_6003_11935# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X721 a_10380_1777# VPWR a_9629_2033# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X722 VGND VPWR a_10046_2143# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X723 a_4915_10549# a_4637_10577# VPWR w_4540_10763# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X724 a_2343_5417# Y VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X725 a_9290_1751# a_8755_1779# a_9515_1777# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X726 a_12976_1743# a_13243_1743# a_13201_2135# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X727 a_5831_1783# VPWR a_5735_1783# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X728 a_24318_14385# a_23731_14309# a_24234_14385# VNB sky130_fd_pr__nfet_01v8 ad=0.10858 pd=1.36 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=4318,272
X729 a_9549_13091# VPWR a_9467_13091# w_9394_13055# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X730 a_9477_11527# VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X731 a_3229_5051# a_2289_5307# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X732 a_6087_14735# a_5809_14763# VPWR w_5712_14949# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X733 VPWR VPWR a_4637_10577# w_4540_10763# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X734 VGND VPWR a_6029_5409# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X735 a_12481_5467# a_11541_5723# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X736 a_11499_2029# a_10569_1777# a_11916_1773# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X737 a_13369_1769# a_13315_2025# a_12976_1743# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X738 a_11427_5467# VPWR a_11331_5467# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X739 VGND VPWR a_13369_2135# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X740 a_4753_16339# VGND VPWR w_4430_16303# sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X741 a_2175_5051# VPWR a_2079_5051# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X742 a_10450_4963# VPWR a_9699_4853# VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X743 VPWR VPWR a_9683_1777# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X744 a_4763_14775# VGND VPWR w_4440_14739# sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X745 a_9360_4571# VPWR a_9585_4963# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X746 sky130_fd_sc_hd__inv_1_5.Y sky130_fd_sc_hd__inv_1_5.A VPWR sky130_fd_sc_hd__inv_1_5.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X747 a_4910_5413# VPWR a_4159_5303# VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X748 a_13439_4955# a_13385_4845# a_13046_4563# VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X749 VPWR VGND a_8596_5039# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X750 a_10088_5837# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X751 a_15017_5825# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X752 a_7899_5405# a_7845_5295# a_7506_5013# VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X753 a_10422_5471# VPWR a_9671_5727# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X754 VGND VPWR a_6362_2149# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X755 VPWR VPWR a_10116_4597# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X756 a_13046_4563# a_13313_4563# a_13271_4589# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X757 a_9332_5445# VGND a_9557_5471# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X758 a_9599_10561# VGND VPWR w_9502_10747# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X759 a_11359_4593# VGND VPWR w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X760 sky130_fd_sc_hd__mux2_1_0.S a_7845_5295# VPWR w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X761 VGND a_3820_5021# a_3768_5047# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X762 a_11595_5833# a_10611_5471# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X763 VPWR VPWR a_7869_1779# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X764 VPWR VPWR a_13439_4589# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X765 a_7506_5013# a_6915_5043# a_7731_5039# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X766 VGND VPWR a_15281_5825# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X767 VGND VGND a_7869_2145# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X768 a_9717_12841# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X769 a_8262_5039# VGND VPWR w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X770 VPWR VGND a_9557_14759# w_9402_14723# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X771 a_9867_12097# a_9589_12125# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X772 VPWR VPWR a_9725_5471# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X773 VPWR VGND a_10380_1777# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X774 a_4839_12857# VPWR a_4755_12857# VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X775 a_3199_1791# a_2259_2047# VPWR w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X776 a_12439_1773# a_11499_2029# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X777 a_9799_16073# a_9465_16323# a_9715_16323# w_9392_16287# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X778 a_12809_13987# a_11243_11891# a_12713_13987# w_12566_13951# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X779 a_2313_2157# a_2259_2047# a_1920_1765# VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X780 VPWR ui_in[1] a_23731_14309# sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.1083 ps=1.36 w=0.42 l=0.15
**devattr s=4332,272 d=4316,272
X781 a_1920_1765# sky130_fd_sc_hd__inv_1_0.Y a_2145_1791# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X782 VPWR VGND a_4585_16339# w_4430_16303# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X783 a_17053_4938# a_16871_4938# VPWR sky130_fd_sc_hd__mux2_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X784 a_12075_13379# a_11824_13629# VPWR w_11718_13593# sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5830,267 d=13600,536
X785 VPWR VGND a_4595_14775# w_4440_14739# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X786 a_7701_2145# VPWR a_7605_2145# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X787 VGND VGND a_10450_4963# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X788 a_15281_5825# a_15227_5715# a_14888_5433# VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X789 a_10046_1777# VGND VPWR w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X790 a_9419_1777# VGND VPWR w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X791 VPWR VPWR a_2313_1791# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X792 a_13105_2135# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X793 VGND VGND a_4910_5413# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X794 a_2706_5051# VGND VPWR w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X795 a_15227_5715# a_14297_5463# a_15644_5459# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X796 sky130_fd_sc_hd__inv_1_5.A sky130_fd_sc_hd__inv_1_4.A VPWR sky130_fd_sc_hd__inv_1_4.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X797 VGND VGND a_6029_5409# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X798 a_14846_1739# a_14255_1769# a_15071_1765# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X799 a_6635_15235# a_6087_14735# VPWR w_6570_15449# sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X800 a_5975_5299# a_5903_5017# a_6392_5043# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X801 a_11553_1773# a_10569_1777# VPWR w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X802 ui_in[0] a_23731_14309# a_23511_14701# sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X803 VPWR VGND a_10422_5471# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X804 VPWR VGND a_9683_1777# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X805 VPWR VPWR a_15239_1765# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X806 a_10116_4963# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X807 a_9489_4963# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X808 a_13385_4845# a_13313_4563# a_13802_4955# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X809 a_24962_14701# ui_in[0] ui_in[0] sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09209 pd=0.99 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=3683,198
X810 a_3919_1787# VGND VPWR w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X811 VPWR a_13046_4563# a_12994_4589# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X812 VGND a_7113_13395# a_7669_14003# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2268,138 d=4075,198
X813 VGND a_9467_13091# a_9801_12841# VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X814 a_10611_5471# a_9671_5727# VPWR w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20523 ps=1.98249 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X815 a_2049_2157# VGND VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X816 a_9557_14759# VPWR a_9475_14759# w_9402_14723# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X817 a_2343_5417# a_2289_5307# a_1950_5025# VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X818 a_7845_5295# a_6915_5043# a_8262_5405# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X819 VPWR a_9332_5445# a_9280_5471# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X820 VGND sky130_fd_sc_hd__inv_1_0.A sky130_fd_sc_hd__inv_1_0.Y VNB sky130_fd_pr__nfet_01v8 ad=0.12778 pd=1.31426 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X821 a_14946_4905# VPWR a_15309_4951# VNB sky130_fd_pr__nfet_01v8 ad=0.07384 pd=0.80236 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X822 VGND VGND a_9753_4963# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X823 VPWR VPWR a_9725_14759# w_9402_14723# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X824 a_13175_4589# VGND VPWR w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X825 a_4849_11293# VPWR a_4765_11293# VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X826 a_13411_5829# a_13285_5437# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08256 ps=0.84921 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X827 a_7731_5405# VPWR a_7635_5405# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X828 a_14297_5463# a_13357_5719# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X829 VPWR VGND a_13439_4589# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X830 a_9461_5471# VGND VPWR w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X831 a_15239_2131# a_15185_2021# a_14846_1739# VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X832 a_3010_2157# VPWR a_2259_2047# VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X833 a_7173_15235# a_6635_15235# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X834 a_13243_5463# VPWR a_13147_5463# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X835 a_5851_13769# a_4837_16089# VPWR w_5786_13983# sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X836 a_4849_11293# a_4515_11543# a_4765_11543# w_4442_11507# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X837 VPWR VGND a_9725_5471# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X838 a_14255_1769# a_13315_2025# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12778 ps=1.31426 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X839 VGND a_4905_12113# a_6089_11935# VNB sky130_fd_pr__nfet_01v8 ad=0.08256 pd=0.84921 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X840 a_4213_5047# a_3229_5051# VPWR w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0862 ps=0.83264 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X841 a_5999_2149# a_5945_2039# a_5606_1757# VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X842 a_4129_2043# a_3199_1791# a_4546_2153# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X843 a_9811_11277# a_9477_11527# a_9727_11527# w_9404_11491# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X844 a_6911_15235# a_6087_14735# a_6805_15235# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X845 VPWR a_4839_12857# a_5851_13769# w_5786_13983# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X846 VPWR a_1950_5025# a_1898_5051# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.20523 pd=1.98249 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X847 a_8566_2145# VPWR a_7815_2035# VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X848 VPWR VPWR a_2676_1791# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X849 VPWR VPWR a_7899_5039# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.0862 pd=0.83264 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
C0 a_7701_1779# sky130_fd_sc_hd__inv_1_0.A 0
C1 a_11291_12911# w_10868_12105# 0
C2 a_2289_5307# a_2706_5417# 0.06611f
C3 sky130_fd_sc_hd__mux2_1_0.A0 w_14736_5374# 0.02073f
C4 a_12994_4589# w_11078_4508# 0.00227f
C5 a_11230_4567# a_11541_5723# 0
C6 a_11916_2139# sky130_fd_sc_hd__inv_1_0.A 0
C7 a_4129_2043# w_3638_1702# 0.10454f
C8 a_2676_2157# VPWR 0.02063f
C9 w_11718_13593# a_9877_10533# 0.00404f
C10 a_4905_12113# a_5975_12927# 0
C11 a_12292_5467# A 0
C12 a_11202_5441# a_11150_5467# 0.1439f
C13 VGND a_5584_5043# 0.08665f
C14 w_9394_13055# a_9467_13091# 0.06993f
C15 a_7731_5405# VPWR 0
C16 a_14066_1769# VGND 0
C17 a_4635_13809# w_4530_12327# 0
C18 ui_in[5] ui_in[6] 0.03102f
C19 a_24318_14385# a_24234_14385# 0.0296f
C20 a_5765_5409# VPWR 0
C21 a_12509_4593# a_13313_4563# 0.02844f
C22 VGND a_5895_14763# 0.00618f
C23 a_13046_4563# a_13018_5437# 0
C24 w_12566_13951# a_11243_11891# 0.03664f
C25 a_9875_13765# a_11351_13753# 0
C26 a_5999_1783# a_5945_2039# 0.00386f
C27 a_6029_5043# a_5903_5017# 0.08094f
C28 a_7845_5295# a_8596_5405# 0.00696f
C29 a_13802_4589# a_13385_4845# 0.03016f
C30 a_13369_2135# VPWR 0.00905f
C31 a_8566_1779# VGND 0
C32 a_4576_5413# w_3668_4962# 0.00139f
C33 w_11050_5382# VGND 0.31674f
C34 a_15255_4841# VPWR 0.35508f
C35 a_5606_1757# w_5454_1698# 0.05213f
C36 a_4753_16339# sky130_fd_sc_hd__inv_1_2.Y 0
C37 VPWR a_9725_5471# 0.16959f
C38 a_9867_12097# a_11243_11891# 0.03573f
C39 a_14946_4905# a_14297_5463# 0.01842f
C40 a_5903_5017# w_3668_4962# 0.00743f
C41 a_14916_4559# w_14764_4500# 0.05213f
C42 a_4763_14775# a_4503_16339# 0
C43 a_11553_2139# sky130_fd_sc_hd__inv_1_0.A 0
C44 a_14946_4905# a_16871_4938# 0.00632f
C45 a_1920_1765# a_2145_1791# 0.00487f
C46 a_11597_15219# a_12135_15219# 0.08446f
C47 sky130_fd_sc_hd__inv_1_0.Y a_1920_1765# 0.08244f
C48 a_9865_15329# w_9392_16287# 0
C49 a_15141_4585# a_14916_4559# 0.00487f
C50 a_10813_13753# a_9811_11277# 0.17627f
C51 VGND VPWR 61.5446f
C52 VPWR a_9799_16073# 1.07863f
C53 a_11178_4593# a_9699_4853# 0
C54 a_14888_5433# a_14297_5463# 0.11887f
C55 a_4913_13781# a_4505_13107# 0
C56 VGND sky130_fd_sc_hd__mux4_1_0.VPB 0.01738f
C57 a_6944_13645# VGND 0
C58 a_8232_1779# a_7815_2035# 0.03016f
C59 a_4513_14775# a_4635_13809# 0.00144f
C60 a_5831_1783# VGND 0
C61 a_11597_15219# a_11767_15219# 0.00167f
C62 a_9727_11277# a_4915_10549# 0
C63 a_14836_5459# w_14736_5374# 0.01793f
C64 a_4129_2043# sky130_fd_sc_hd__inv_1_0.Y 0.00305f
C65 a_6635_15235# VPWR 0.33595f
C66 a_6281_11907# VGND 0.5959f
C67 a_12135_15219# a_10771_14747# 0
C68 a_4915_10549# a_7847_14003# 0
C69 a_13802_4589# a_13285_5437# 0
C70 a_6862_13645# a_4837_16089# 0
C71 a_5831_2149# VGND 0.00231f
C72 sky130_fd_sc_hd__inv_1_2.A VGND 0.70676f
C73 sky130_fd_sc_hd__inv_1_2.A a_9799_16073# 0
C74 a_4915_10549# a_6089_11935# 0
C75 a_11623_4593# a_11986_4593# 0.00985f
C76 a_7476_1753# a_7815_2035# 0.04737f
C77 a_17125_4938# A 0.1015f
C78 a_15644_5825# VGND 0.18635f
C79 a_4837_16089# w_4528_15559# 0.00251f
C80 a_9515_2143# sky130_fd_sc_hd__inv_1_0.A 0
C81 a_14136_4589# sky130_fd_sc_hd__inv_1_0.A 0
C82 ua[4] a_15071_1765# 0
C83 a_4765_11543# a_4849_11293# 0.08177f
C84 a_4503_16339# sky130_fd_sc_hd__inv_1_2.Y 0
C85 a_9809_14509# a_11597_15219# 0.17824f
C86 VPWR a_15239_1765# 0.17252f
C87 a_14066_2135# sky130_fd_sc_hd__inv_1_0.A 0
C88 a_11230_4567# w_11078_4508# 0.05213f
C89 a_10088_5837# A 0.00192f
C90 a_3199_1791# a_4129_2043# 0.21188f
C91 w_9394_13055# VPWR 0.16326f
C92 a_7845_5295# a_7731_5405# 0
C93 a_9360_4571# w_9208_4512# 0.05213f
C94 a_13046_4563# a_13175_4955# 0.00792f
C95 a_4913_13781# w_5906_12121# 0
C96 a_23677_14335# VGND 0.00194f
C97 a_14255_1769# VPWR 1.04578f
C98 a_12924_1769# w_12824_1684# 0.01793f
C99 w_6756_13609# a_7173_15235# 0
C100 a_1920_1765# a_2313_1791# 0.02283f
C101 a_2289_5307# w_1798_4966# 0.10454f
C102 w_12866_5378# a_13018_5437# 0.05213f
C103 a_10639_4597# a_11569_4849# 0.21188f
C104 a_4765_11293# VGND 0.00834f
C105 VGND a_12809_13987# 0
C106 a_5809_14763# w_5910_13141# 0
C107 a_6911_15235# a_6087_14735# 0.00651f
C108 a_11230_4567# a_11455_4593# 0.00487f
C109 a_11385_1773# VPWR 0
C110 a_15309_4585# a_14297_5463# 0
C111 a_4627_12141# a_4765_11543# 0
C112 a_11916_1773# a_13243_1743# 0
C113 a_15281_5459# a_14297_5463# 0.08312f
C114 a_7476_1753# a_5945_2039# 0.00446f
C115 a_3790_1761# w_3638_1702# 0.05213f
C116 a_17125_5265# VPWR 0
C117 VGND ui_in[1] 0.11268f
C118 a_17125_4938# sky130_fd_sc_hd__mux2_1_0.A0 0.06947f
C119 a_11873_15219# VGND 0.00384f
C120 a_11873_15219# a_9799_16073# 0.00241f
C121 a_9809_14509# a_10771_14747# 0.00524f
C122 a_9238_1777# a_9290_1751# 0.1439f
C123 VGND a_4585_16339# 0.00117f
C124 a_11427_5833# A 0
C125 a_2049_1791# VPWR 0.00125f
C126 a_14297_5463# sky130_fd_sc_hd__mux2_1_0.S 0.04835f
C127 a_10639_4597# a_11595_5833# 0
C128 a_7845_5295# a_9725_5471# 0
C129 a_7605_1779# a_7869_1779# 0
C130 a_10813_13753# w_10748_13967# 0.08205f
C131 a_16871_4938# sky130_fd_sc_hd__mux2_1_0.S 0.25154f
C132 VPWR a_17346_5265# 0
C133 a_13175_4589# a_13313_4563# 0
C134 a_13046_4563# a_12509_4593# 0
C135 w_14694_1680# a_15602_2131# 0.00139f
C136 a_2676_1791# w_1768_1706# 0.01154f
C137 a_4635_13809# a_4839_12857# 0.00246f
C138 a_4849_11293# a_5975_12927# 0.18651f
C139 a_15239_2131# VPWR 0.00775f
C140 w_5786_13983# a_5975_12927# 0
C141 a_6003_11935# a_4905_12113# 0.18618f
C142 a_24962_14701# ua[0] 0.13397f
C143 a_11019_12911# VGND 0.00238f
C144 a_15045_4951# a_15309_4951# 0
C145 a_7845_5295# VGND 1.20783f
C146 a_5809_14763# w_5712_14949# 0.05631f
C147 a_11986_4959# w_11078_4508# 0.00139f
C148 a_9801_12841# a_11824_13629# 0.00327f
C149 a_4849_11293# w_6756_13609# 0
C150 a_3820_5021# VPWR 0.29445f
C151 a_9867_12097# a_9811_11277# 0.25265f
C152 a_17339_4938# VGND 0
C153 a_8566_2145# a_7815_2035# 0.00696f
C154 a_6862_13645# a_5851_13769# 0
C155 a_11553_1773# sky130_fd_sc_hd__inv_1_0.A 0
C156 a_9308_4597# A 0
C157 w_9500_13979# VGND 0.11975f
C158 a_9875_13765# a_10771_14747# 0
C159 a_10088_5837# a_9671_5727# 0.06611f
C160 a_11623_4593# a_10611_5471# 0
C161 w_14694_1680# a_13315_2025# 0
C162 a_2706_5051# a_2343_5051# 0.00985f
C163 a_9559_11527# VGND 0.00172f
C164 a_5999_1783# VGND 0.01528f
C165 a_8113_13753# a_11351_13753# 0
C166 a_5554_1783# w_5454_1698# 0.01793f
C167 a_4763_14775# a_4847_14525# 0.07979f
C168 VGND a_9549_13091# 0.00171f
C169 a_15672_4585# w_14764_4500# 0.01154f
C170 w_11050_5382# a_11541_5723# 0.10454f
C171 sky130_fd_sc_hd__inv_1_5.A VGND 0.27564f
C172 sky130_fd_sc_hd__inv_1_0.Y a_4880_1787# 0
C173 a_7506_5013# a_6915_5043# 0.11887f
C174 w_11050_5382# a_12966_5463# 0.00227f
C175 a_3790_1761# sky130_fd_sc_hd__inv_1_0.Y 0.00242f
C176 a_24774_14701# ua[0] 0.00406f
C177 a_4903_15345# a_4625_15373# 0.12165f
C178 w_3638_1702# VPWR 0.51511f
C179 a_10857_14747# a_9811_11277# 0.00121f
C180 a_4755_12857# VGND 0.00847f
C181 VGND a_9715_16323# 0.01705f
C182 a_13385_4845# a_13285_5437# 0
C183 a_9489_4963# A 0
C184 a_4915_10549# a_7751_14003# 0
C185 a_9715_16323# a_9799_16073# 0.07445f
C186 a_13732_1769# a_13243_1743# 0.08907f
C187 w_6570_15449# a_7173_15235# 0.01567f
C188 a_11499_2029# w_12824_1684# 0
C189 w_10872_13125# a_10937_12911# 0.04996f
C190 a_14846_1739# a_13315_2025# 0.00446f
C191 VGND a_4763_14525# 0.00834f
C192 a_13802_4589# sky130_fd_sc_hd__inv_1_0.A 0
C193 a_15045_4951# a_14946_4905# 0.0029f
C194 VPWR a_11541_5723# 0.33241f
C195 a_11049_14719# a_9475_14759# 0
C196 a_3199_1791# a_3790_1761# 0.11887f
C197 a_4513_14775# a_5809_14763# 0
C198 VPWR a_12966_5463# 0.06844f
C199 a_8596_5405# A 0
C200 VPWR sky130_fd_sc_hd__inv_1_4.VPB 0.07223f
C201 w_5484_4958# a_5903_5017# 0.24672f
C202 a_12135_15219# w_11718_13593# 0
C203 a_11150_5467# w_9180_5386# 0.00188f
C204 a_13439_4589# a_13271_4589# 0
C205 a_4847_14525# a_4505_13107# 0
C206 sky130_fd_sc_hd__inv_1_2.Y a_4847_14525# 0.29596f
C207 VGND a_10895_13753# 0.00382f
C208 a_9589_12125# a_9867_12097# 0.1206f
C209 a_10895_13753# a_9799_16073# 0
C210 a_6389_13769# a_6127_13769# 0
C211 VGND a_11243_11891# 0.5959f
C212 a_2175_5417# a_2289_5307# 0
C213 a_15978_5825# VGND 0.00228f
C214 a_11958_5467# a_10611_5471# 0.08907f
C215 a_13439_4589# a_13313_4563# 0.08094f
C216 VGND a_9515_1777# 0
C217 a_9699_4853# a_9585_4963# 0
C218 a_9629_2033# w_9138_1692# 0.10454f
C219 a_3768_5047# VGND 0.08661f
C220 w_4430_16303# a_4903_15345# 0
C221 a_13175_4589# a_13046_4563# 0.00758f
C222 w_10674_14933# VGND 0.0161f
C223 a_10116_4597# VGND 0.01145f
C224 w_10674_14933# a_9799_16073# 0.00872f
C225 a_9467_13091# w_9492_12311# 0.0035f
C226 a_8232_1779# VGND 0.01329f
C227 a_4045_5047# a_3229_5051# 0
C228 a_9477_11527# a_9867_12097# 0
C229 a_6885_1783# a_7701_1779# 0
C230 a_7605_1779# VPWR 0.00115f
C231 a_7506_5013# a_9360_4571# 0
C232 VGND a_4910_5413# 0.00246f
C233 a_6392_5043# a_5903_5017# 0.08907f
C234 VGND a_10983_13753# 0.00475f
C235 a_10983_13753# a_9799_16073# 0.00246f
C236 a_4903_15345# w_4538_13995# 0.00397f
C237 a_5861_5409# VPWR 0
C238 a_11916_2139# w_11008_1688# 0.00139f
C239 a_7476_1753# VGND 0.40126f
C240 a_2145_1791# VPWR 0.00107f
C241 a_9875_13765# a_11291_12911# 0.0204f
C242 a_13201_1769# VPWR 0
C243 sky130_fd_sc_hd__inv_1_0.Y VPWR 1.34565f
C244 a_6057_12927# VPWR 0
C245 a_9332_5445# a_9557_5471# 0.00487f
C246 a_9809_14509# w_11718_13593# 0
C247 VGND a_2343_5417# 0.20137f
C248 a_9717_12841# VGND 0.00847f
C249 a_9801_12841# a_11089_13753# 0.00253f
C250 a_6389_13769# a_7751_14003# 0
C251 a_4913_13781# w_5910_13141# 0.09336f
C252 w_9392_16287# a_9587_15357# 0
C253 sky130_fd_sc_hd__inv_1_0.Y a_5831_1783# 0
C254 a_9801_12841# a_9467_13091# 0.16952f
C255 a_6003_11935# a_4849_11293# 0.10332f
C256 a_9683_2143# VGND 0.20145f
C257 a_5809_14763# a_4839_12857# 0.21988f
C258 a_2706_5417# VPWR 0.01961f
C259 a_9865_15329# a_11824_13629# 0
C260 VGND a_23731_14309# 0.12017f
C261 a_8113_13753# a_11597_15219# 0.1684f
C262 a_9629_2033# sky130_fd_sc_hd__inv_1_0.A 0.00296f
C263 a_4765_11543# a_4637_10577# 0
C264 a_15071_1765# VPWR 0
C265 w_12866_5378# a_13774_5829# 0.00139f
C266 a_5831_2149# sky130_fd_sc_hd__inv_1_0.Y 0
C267 a_13411_5829# VPWR 0.00606f
C268 a_9332_5445# a_9280_5471# 0.1439f
C269 a_15045_4585# a_14916_4559# 0.00758f
C270 a_7731_5405# A 0
C271 a_3199_1791# VPWR 1.05387f
C272 a_9725_14509# VGND 0.00834f
C273 a_11427_5833# a_11595_5833# 0
C274 Y a_2706_5051# 0.08994f
C275 sky130_fd_sc_hd__mux2_1_0.S a_13018_5437# 0
C276 VGND a_13147_5829# 0.00333f
C277 a_9465_16323# a_9715_16073# 0.00723f
C278 a_11230_4567# a_9699_4853# 0.00446f
C279 a_4903_15345# a_5895_14763# 0
C280 a_5735_1783# a_5873_1757# 0
C281 a_6003_11935# a_4627_12141# 0
C282 a_9419_2143# VPWR 0
C283 w_9490_15543# a_9475_14759# 0
C284 a_11553_2139# w_11008_1688# 0
C285 a_6127_13769# a_4839_12857# 0.00253f
C286 w_11078_4508# VPWR 0.52749f
C287 a_15017_5459# VPWR 0.00132f
C288 a_8113_13753# a_10771_14747# 0
C289 a_4913_13781# w_5712_14949# 0
C290 sky130_fd_sc_hd__mux2_1_0.S a_11202_5441# 0
C291 a_15255_4841# A 0
C292 w_4432_13071# a_4635_13809# 0.00101f
C293 VGND a_23511_14701# 0.00202f
C294 a_9725_5471# A 0
C295 a_9867_12097# a_9675_12125# 0
C296 a_9475_14759# w_9402_14723# 0.06993f
C297 a_2313_1791# VPWR 0.17194f
C298 a_11455_4593# VPWR 0.00101f
C299 a_13369_2135# a_13315_2025# 0.03622f
C300 a_15602_2131# VGND 0.18859f
C301 a_12320_4593# VGND 0
C302 a_13385_4845# sky130_fd_sc_hd__inv_1_0.A 0
C303 a_4213_5413# w_3668_4962# 0
C304 a_14946_4905# a_15644_5459# 0.00474f
C305 VPWR w_9492_12311# 0.17848f
C306 a_3768_5047# a_3820_5021# 0.1439f
C307 a_11051_11919# VPWR 0
C308 a_8566_2145# VGND 0.00244f
C309 a_4903_15345# VPWR 0.24554f
C310 VGND A 2.34296f
C311 sky130_fd_sc_hd__inv_1_5.A sky130_fd_sc_hd__inv_1_4.VPB 0.02727f
C312 VPWR a_23677_14701# 0.18463f
C313 a_5873_1757# a_5069_1787# 0.02844f
C314 a_23677_14701# sky130_fd_sc_hd__mux4_1_0.VPB 0.01733f
C315 a_11385_2139# VPWR 0
C316 a_9585_4963# a_9753_4963# 0
C317 a_6087_14735# VGND 0.35053f
C318 a_6329_12927# a_4505_13107# 0
C319 a_13439_4589# a_13046_4563# 0.02283f
C320 a_15255_4841# sky130_fd_sc_hd__mux2_1_0.A0 0
C321 a_10813_13753# a_11351_13753# 0.07901f
C322 VGND a_9811_11277# 1.26863f
C323 a_9597_13793# a_9475_14759# 0.00144f
C324 a_14946_4905# a_14136_4955# 0
C325 a_9811_11277# a_9799_16073# 0.03118f
C326 w_7604_13967# a_7669_14003# 0.05168f
C327 a_13315_2025# VGND 1.19935f
C328 a_17053_4938# sky130_fd_sc_hd__mux2_1_0.A1 0.00136f
C329 a_10965_11919# a_9867_12097# 0.18618f
C330 sky130_fd_sc_hd__inv_1_2.A a_23677_14701# 0
C331 a_13357_5719# VGND 1.20852f
C332 a_6087_14735# a_6635_15235# 0.08954f
C333 ui_in[0] sky130_fd_sc_hd__inv_1_0.A 0.24408f
C334 a_6389_13769# a_4913_13781# 0
C335 a_9801_12841# VPWR 0.75043f
C336 a_4837_16089# a_6021_13769# 0.00246f
C337 a_15602_2131# a_14255_1769# 0.03325f
C338 a_4183_2153# a_4546_2153# 0.00847f
C339 a_11230_4567# a_10611_5471# 0
C340 a_14325_4589# a_15227_5715# 0
C341 a_5999_2149# VPWR 0.00848f
C342 a_5903_5017# a_5584_5043# 0.04799f
C343 a_4513_14775# a_4913_13781# 0
C344 a_5999_1783# sky130_fd_sc_hd__inv_1_0.Y 0
C345 sky130_fd_sc_hd__mux2_1_0.A0 VGND 0.40622f
C346 a_13105_1769# a_13243_1743# 0
C347 a_9489_4597# a_9753_4597# 0
C348 a_7113_13395# VGND 0.35166f
C349 a_14846_1739# w_12824_1684# 0
C350 VGND a_4587_13107# 0.00171f
C351 a_9671_5727# a_9725_5471# 0.00386f
C352 a_6329_12927# w_5906_12121# 0
C353 a_9699_4853# a_9753_4597# 0.00386f
C354 w_9394_13055# a_9811_11277# 0.00299f
C355 a_15281_5825# a_15227_5715# 0.03622f
C356 a_5831_2149# a_5999_2149# 0
C357 a_12135_15219# a_11049_14719# 0.00425f
C358 a_4755_13107# VPWR 0.31944f
C359 a_6635_15235# a_7113_13395# 0
C360 VPWR w_1798_4966# 0.51758f
C361 a_7424_1779# sky130_fd_sc_hd__inv_1_0.A 0.00118f
C362 a_9865_15329# a_11089_13753# 0
C363 a_17125_5265# A 0
C364 a_9557_14759# VPWR 0.02511f
C365 a_14255_1769# a_13315_2025# 0.13962f
C366 a_13439_4955# a_13385_4845# 0.03622f
C367 ui_in[1] a_23677_14701# 0.02095f
C368 a_4513_14775# a_4503_16339# 0.00102f
C369 a_15602_2131# a_15239_2131# 0.00847f
C370 a_24318_14385# VGND 0.09477f
C371 a_7869_1779# a_7701_1779# 0
C372 ua[0] VPWR 0.07056f
C373 a_9671_5727# VGND 1.46609f
C374 A a_17346_5265# 0.00101f
C375 ua[0] sky130_fd_sc_hd__mux4_1_0.VPB 0.02132f
C376 a_15281_5459# a_15644_5459# 0.00985f
C377 a_14325_4589# a_13802_4589# 0
C378 a_9683_1777# a_9290_1751# 0.02283f
C379 a_14794_1765# VPWR 0.07423f
C380 a_11824_13629# a_12075_13379# 0.10945f
C381 a_6129_12927# a_5975_12927# 0.00401f
C382 a_11049_14719# a_11767_15219# 0.00366f
C383 a_9461_5837# a_9725_5837# 0
C384 a_4576_5413# VPWR 0.01963f
C385 VGND w_10748_13967# 0.01862f
C386 w_10748_13967# a_9799_16073# 0.06973f
C387 a_11553_1773# w_11008_1688# 0.01092f
C388 a_9589_12125# VGND 0.24254f
C389 sky130_fd_sc_hd__mux2_1_0.VPB VPWR 0.1138f
C390 a_11986_4959# a_10611_5471# 0
C391 a_5903_5017# VPWR 0.97115f
C392 a_5765_5043# VGND 0
C393 a_4849_11293# a_4905_12113# 0.25265f
C394 uio_out[6] uio_out[5] 0.03102f
C395 uo_out[1] uo_out[2] 0.03102f
C396 a_7506_5013# a_7731_5039# 0.00487f
C397 sky130_fd_sc_hd__mux2_1_0.S a_6915_5043# 0
C398 w_12566_13951# a_11351_13753# 0
C399 a_17125_5265# sky130_fd_sc_hd__mux2_1_0.A0 0.00576f
C400 a_7454_5039# VGND 0.08651f
C401 a_9809_14509# a_11049_14719# 0.3196f
C402 a_12250_2139# sky130_fd_sc_hd__inv_1_0.A 0
C403 a_4913_13781# a_4839_12857# 0.44871f
C404 a_12631_13987# a_11824_13629# 0
C405 a_9477_11527# VGND 0.29765f
C406 sky130_fd_sc_hd__mux2_1_0.A0 a_17346_5265# 0
C407 a_7899_5039# a_6915_5043# 0.08312f
C408 a_13802_4955# a_13385_4845# 0.06611f
C409 a_5851_13769# a_6021_13769# 0.00167f
C410 a_13147_5829# a_12966_5463# 0
C411 a_13439_4955# a_13285_5437# 0
C412 a_15185_2021# sky130_fd_sc_hd__inv_1_0.A 0.1531f
C413 a_7476_1753# a_7605_1779# 0.00758f
C414 w_7604_13967# VPWR 0.07722f
C415 a_4576_5047# a_4213_5047# 0.00985f
C416 a_9801_12841# a_11019_12911# 0.00149f
C417 VGND a_14836_5459# 0.08665f
C418 a_4627_12141# a_4905_12113# 0.1206f
C419 a_9589_12125# w_9394_13055# 0
C420 a_2079_5417# VGND 0.00311f
C421 sky130_fd_sc_hd__inv_1_0.A w_9138_1692# 0.00331f
C422 a_13243_5463# VGND 0
C423 ua[0] ui_in[1] 0.36102f
C424 a_9801_12841# w_9500_13979# 0.00445f
C425 w_7604_13967# a_6281_11907# 0.03664f
C426 a_7635_5405# VPWR 0
C427 a_4847_14525# w_5712_14949# 0.00381f
C428 a_9332_5445# a_9557_5837# 0.00559f
C429 a_9875_13765# a_11049_14719# 0
C430 a_1868_1791# w_1768_1706# 0.01793f
C431 w_9394_13055# a_9477_11527# 0
C432 a_5873_1757# sky130_fd_sc_hd__inv_1_0.A 0
C433 a_9801_12841# a_9549_13091# 0
C434 a_4903_15345# a_4763_14525# 0
C435 a_11541_5723# A 0.00769f
C436 a_14864_4585# VGND 0
C437 a_13774_5463# VGND 0.01425f
C438 a_10380_2143# a_9629_2033# 0.00696f
C439 a_11569_4849# VGND 1.20507f
C440 a_2343_5417# a_2706_5417# 0.00847f
C441 a_10813_13753# a_10771_14747# 0
C442 VGND a_9683_13793# 0.00661f
C443 a_13802_4955# a_13285_5437# 0
C444 a_6362_1783# a_5873_1757# 0.08907f
C445 a_9865_15329# VPWR 0.24549f
C446 a_12966_5463# A 0.00303f
C447 a_11986_4593# VPWR 0.20848f
C448 a_3040_5051# a_2289_5307# 0.00682f
C449 a_9489_4597# VPWR 0.0015f
C450 uio_out[2] uio_out[1] 0.03102f
C451 a_4837_16089# sky130_fd_sc_hd__inv_1_2.Y 0.27498f
C452 a_13369_2135# w_12824_1684# 0
C453 a_9360_4571# sky130_fd_sc_hd__mux2_1_0.S 0
C454 VGND a_11595_5833# 0.20021f
C455 a_4915_10549# a_7919_14003# 0
C456 a_13732_2135# sky130_fd_sc_hd__inv_1_0.A 0
C457 VGND a_9725_14759# 0.02642f
C458 a_9699_4853# VPWR 0.60063f
C459 a_7424_1779# w_7324_1694# 0.01793f
C460 a_11051_11919# a_11243_11891# 0
C461 a_7506_5013# a_7635_5039# 0.00758f
C462 a_9290_1751# a_7815_2035# 0.00511f
C463 a_7899_5039# a_9360_4571# 0
C464 VGND a_6805_15235# 0.00334f
C465 a_9675_12125# VGND 0.00662f
C466 a_4849_11293# a_7173_15235# 0
C467 a_15255_4841# w_14764_4500# 0.10454f
C468 a_6362_1783# sky130_fd_sc_hd__inv_1_0.A 0
C469 a_13147_5829# a_13411_5829# 0
C470 a_9419_2143# a_9683_2143# 0
C471 a_2175_5417# VPWR 0
C472 VGND a_12713_13987# 0
C473 a_11160_1747# a_11499_2029# 0.04737f
C474 w_5786_13983# a_7173_15235# 0
C475 a_5975_5299# a_5636_5017# 0.04737f
C476 a_6389_13769# a_4847_14525# 0
C477 a_6635_15235# a_6805_15235# 0.00167f
C478 sky130_fd_sc_hd__mux2_1_0.S w_9180_5386# 0.00671f
C479 a_9727_11527# a_9467_13091# 0
C480 a_7701_1779# VPWR 0
C481 a_15255_4841# a_15141_4585# 0
C482 VGND w_12824_1684# 0.29354f
C483 a_11427_5467# a_11202_5441# 0.00487f
C484 a_9801_12841# a_10895_13753# 0
C485 a_4513_14775# a_4847_14525# 0.1679f
C486 a_14325_4589# a_13385_4845# 0.13962f
C487 a_13439_4589# a_14946_4905# 0
C488 a_4837_16089# w_5906_12121# 0
C489 a_11916_2139# VPWR 0.01968f
C490 a_4635_13809# VGND 0.24546f
C491 a_9801_12841# a_11243_11891# 0.02336f
C492 a_13147_5463# VPWR 0.00103f
C493 a_10639_4597# w_9208_4512# 0.02026f
C494 a_16006_4951# a_14946_4905# 0.0022f
C495 a_9809_14509# w_9402_14723# 0.02435f
C496 a_11553_1773# a_11289_1773# 0
C497 VGND w_14764_4500# 0.00461f
C498 a_9629_2033# w_11008_1688# 0
C499 a_9801_12841# w_10674_14933# 0.08813f
C500 a_10965_11919# VGND 0.13487f
C501 Y a_3040_5417# 0
C502 w_11050_5382# a_10611_5471# 0.25055f
C503 a_10965_11919# a_9799_16073# 0
C504 a_2676_1791# VPWR 0.20903f
C505 a_6329_12927# w_5910_13141# 0.02303f
C506 a_8262_5039# w_7354_4954# 0.01154f
C507 a_13313_4563# a_10639_4597# 0
C508 a_13201_1769# a_13315_2025# 0
C509 a_9801_12841# a_10983_13753# 0
C510 a_23731_14309# a_23677_14701# 0.09132f
C511 a_13411_5829# A 0.00117f
C512 a_9465_16323# a_9475_14759# 0.00102f
C513 uio_in[6] uio_in[5] 0.03102f
C514 a_7669_14003# w_6756_13609# 0
C515 Y a_3949_5047# 0
C516 a_24241_14651# a_24407_14651# 0.00988f
C517 a_4849_11293# w_5786_13983# 0.10705f
C518 a_3768_5047# w_1798_4966# 0.00188f
C519 a_12439_1773# a_13243_1743# 0.02844f
C520 a_11958_5467# a_13285_5437# 0
C521 a_14255_1769# w_12824_1684# 0.02026f
C522 a_11108_1773# a_9629_2033# 0
C523 a_9801_12841# a_9717_12841# 0.00208f
C524 a_9809_14509# a_9597_13793# 0
C525 a_15644_5459# a_14297_5463# 0.08907f
C526 a_8113_13753# a_7919_14003# 0
C527 a_10611_5471# VPWR 1.069f
C528 a_13201_2135# a_13369_2135# 0
C529 a_11553_2139# VPWR 0.00968f
C530 VGND a_4045_5047# 0
C531 a_9875_13765# w_9402_14723# 0
C532 a_11595_5467# a_11427_5467# 0
C533 a_15017_5459# A 0
C534 w_11078_4508# A 0
C535 a_13802_4589# w_12894_4504# 0.01154f
C536 a_13357_5719# a_13411_5829# 0.03622f
C537 a_10813_13753# a_11291_12911# 0
C538 a_4627_12141# a_4849_11293# 0.0022f
C539 a_9801_12841# a_9725_14509# 0
C540 a_6362_2149# a_5945_2039# 0.06611f
C541 a_9865_15329# w_9500_13979# 0.00397f
C542 a_10937_12911# w_10868_12105# 0
C543 a_5933_13769# a_6389_13769# 0
C544 a_23511_14701# a_23677_14701# 0.05551f
C545 a_12976_1743# sky130_fd_sc_hd__inv_1_0.A 0.00202f
C546 a_7845_5295# a_9699_4853# 0
C547 a_4847_14525# a_4839_12857# 0.20053f
C548 a_15672_4951# a_15309_4951# 0.00847f
C549 a_4765_11543# VPWR 0.31817f
C550 a_2343_5417# w_1798_4966# 0
C551 a_11178_4593# sky130_fd_sc_hd__inv_1_0.A 0
C552 a_2145_2157# a_2313_2157# 0
C553 w_12866_5378# a_12481_5467# 0.0025f
C554 a_10569_1777# a_11160_1747# 0.11887f
C555 VPWR a_4753_16089# 0.00472f
C556 a_13201_2135# VGND 0.00231f
C557 a_9875_13765# a_9597_13793# 0.1205f
C558 a_15309_4951# sky130_fd_sc_hd__mux2_1_0.A1 0
C559 a_9753_4963# VPWR 0.05505f
C560 a_9727_11277# VGND 0.00834f
C561 a_5851_13769# w_5906_12121# 0
C562 w_4432_13071# a_4913_13781# 0.00226f
C563 a_9727_11527# VPWR 0.31817f
C564 a_7847_14003# VGND 0
C565 sky130_fd_sc_hd__inv_1_0.A w_7324_1694# 0.00331f
C566 a_23677_14701# A 0
C567 a_4576_5047# w_3668_4962# 0.01154f
C568 VGND a_6089_11935# 0.00568f
C569 a_10857_14747# a_10771_14747# 0.00658f
C570 a_8113_13753# a_11049_14719# 0.09735f
C571 VPWR a_12075_13379# 0.24586f
C572 a_9811_11277# w_9492_12311# 0.00145f
C573 a_6087_14735# a_4903_15345# 0
C574 a_23731_14309# ua[0] 0
C575 a_9515_2143# VPWR 0
C576 a_14136_4589# VPWR 0
C577 a_11051_11919# a_9811_11277# 0
C578 a_11623_4593# sky130_fd_sc_hd__inv_1_0.A 0
C579 a_11569_4849# a_11541_5723# 0.00177f
C580 a_10813_13753# w_11718_13593# 0.00132f
C581 a_14066_2135# VPWR 0
C582 a_13369_1769# VGND 0.01514f
C583 a_5975_5299# a_6915_5043# 0.13962f
C584 VGND a_11351_13753# 0.25955f
C585 sky130_fd_sc_hd__inv_1_2.A a_12075_13379# 0.03027f
C586 a_11351_13753# a_9799_16073# 0.00515f
C587 a_24962_14701# ui_in[0] 0.12838f
C588 a_4213_5047# w_3668_4962# 0.01092f
C589 a_5975_12927# VPWR 0.1592f
C590 a_10380_1777# VGND 0
C591 a_6389_13769# a_6329_12927# 0.20048f
C592 a_11595_5833# a_11541_5723# 0.03622f
C593 a_12631_13987# VPWR 0.07848f
C594 a_4903_15345# a_7113_13395# 0
C595 a_24241_14651# sky130_fd_sc_hd__inv_1_5.Y 0
C596 a_6885_1783# a_7424_1779# 0.0725f
C597 a_9547_16323# VPWR 0.0251f
C598 a_9801_12841# a_9811_11277# 0.82158f
C599 a_4129_2043# a_4183_1787# 0.00386f
C600 a_15672_4951# a_14946_4905# 0.18442f
C601 a_11906_13629# a_11824_13629# 0.00477f
C602 a_9865_15329# a_10895_13753# 0.0035f
C603 a_17053_4938# a_17125_4938# 0
C604 a_6281_11907# a_5975_12927# 0
C605 w_6756_13609# VPWR 0.08767f
C606 a_5933_13769# a_4839_12857# 0
C607 VGND a_14108_5829# 0.00248f
C608 sky130_fd_sc_hd__inv_1_2.A a_12631_13987# 0.10369f
C609 a_14946_4905# sky130_fd_sc_hd__mux2_1_0.A1 0.08128f
C610 a_3010_1791# VPWR 0
C611 a_4849_11293# w_4440_14739# 0.00324f
C612 a_15309_4951# a_14916_4559# 0.02301f
C613 w_10674_14933# a_9865_15329# 0.00546f
C614 a_13105_2135# sky130_fd_sc_hd__inv_1_0.A 0
C615 a_12809_13987# a_12075_13379# 0.00121f
C616 a_7899_5405# a_6915_5043# 0.04534f
C617 a_3820_5021# a_4045_5047# 0.00487f
C618 w_6756_13609# a_6281_11907# 0.00315f
C619 VGND a_5809_14763# 0.13243f
C620 a_1868_1791# a_1920_1765# 0.1439f
C621 a_24774_14701# ui_in[0] 0.63058f
C622 a_9290_1751# VGND 0.40141f
C623 a_4915_10549# a_9597_13793# 0.00124f
C624 a_9865_15329# a_10983_13753# 0.00818f
C625 a_7731_5039# a_7899_5039# 0
C626 a_13439_4955# a_13802_4955# 0.00847f
C627 a_10116_4597# a_9699_4853# 0.03016f
C628 a_10450_4963# a_10639_4597# 0
C629 a_9589_12125# w_9492_12311# 0.05631f
C630 a_2313_2157# w_1768_1706# 0
C631 a_11553_1773# VPWR 0.17705f
C632 Y a_5975_5299# 0
C633 sky130_fd_sc_hd__mux2_1_0.VPB A 0.03021f
C634 a_4837_16089# w_5910_13141# 0
C635 a_12631_13987# a_12809_13987# 0.00412f
C636 a_7845_5295# a_9753_4963# 0
C637 a_5903_5017# A 0
C638 a_6129_12927# a_4905_12113# 0
C639 a_13315_2025# a_14794_1765# 0
C640 a_6127_13769# VGND 0.00413f
C641 a_15227_5715# VPWR 0.32967f
C642 a_4015_2153# VGND 0.00231f
C643 a_10380_2143# sky130_fd_sc_hd__inv_1_0.A 0
C644 a_13385_4845# w_12894_4504# 0.10454f
C645 a_11595_5467# a_11202_5441# 0.02283f
C646 a_14325_4589# sky130_fd_sc_hd__inv_1_0.A 0
C647 a_6696_2149# a_5945_2039# 0.00696f
C648 sky130_fd_sc_hd__inv_1_2.Y w_4528_15559# 0
C649 VGND sky130_fd_sc_hd__inv_1_0.VPB 0.02955f
C650 VPWR a_9587_15357# 0.38646f
C651 a_4129_2043# a_5069_1787# 0.12975f
C652 a_8113_13753# w_9490_15543# 0.00459f
C653 VPWR a_4213_5413# 0.00874f
C654 a_9477_11527# w_9492_12311# 0
C655 a_13018_5437# a_13243_5829# 0.00559f
C656 a_9585_4597# VGND 0
C657 a_9865_15329# a_9725_14509# 0
C658 a_9801_12841# w_10748_13967# 0.08124f
C659 a_6329_12927# a_4839_12857# 0.08252f
C660 a_11455_4959# VGND 0.00209f
C661 a_13385_4845# a_13271_4955# 0
C662 a_9801_12841# a_9589_12125# 0
C663 a_11160_1747# a_11289_2139# 0.00792f
C664 a_7476_1753# a_7701_1779# 0.00487f
C665 a_2175_5417# a_2343_5417# 0
C666 a_4837_16089# a_4915_10549# 0.01618f
C667 a_15644_5825# a_15227_5715# 0.06611f
C668 a_15141_4951# sky130_fd_sc_hd__mux2_1_0.A1 0
C669 a_14916_4559# a_14946_4905# 0.38909f
C670 a_8113_13753# w_9402_14723# 0.00353f
C671 a_11569_4849# w_11078_4508# 0.10454f
C672 a_12994_4589# sky130_fd_sc_hd__inv_1_0.A 0
C673 a_9332_5445# VPWR 0.29533f
C674 uio_oe[1] uio_oe[2] 0.03102f
C675 a_9308_4597# w_9208_4512# 0.01793f
C676 w_11532_15433# a_11824_13629# 0
C677 a_6362_2149# VGND 0.18643f
C678 sky130_fd_sc_hd__mux2_1_0.A0 sky130_fd_sc_hd__mux2_1_0.VPB 0.1118f
C679 a_7899_5405# a_8262_5405# 0.00847f
C680 a_4837_16089# w_5712_14949# 0.00872f
C681 a_7751_14003# VGND 0
C682 a_15672_4951# sky130_fd_sc_hd__mux2_1_0.S 0
C683 a_6885_1783# a_5873_1757# 0
C684 a_14946_4905# a_15978_5459# 0
C685 a_7635_5405# A 0
C686 a_13802_4589# VPWR 0.2102f
C687 a_7701_2145# sky130_fd_sc_hd__inv_1_0.A 0
C688 a_9801_12841# a_9477_11527# 0
C689 a_11569_4849# a_11455_4593# 0
C690 a_16006_4585# a_14946_4905# 0
C691 a_11597_15219# VGND 0.13063f
C692 a_11108_1773# w_9138_1692# 0.00188f
C693 a_9461_5471# VPWR 0.00116f
C694 a_11597_15219# a_9799_16073# 0.232f
C695 a_14916_4559# a_14888_5433# 0
C696 a_4849_11293# a_4637_10577# 0
C697 sky130_fd_sc_hd__mux2_1_0.A1 sky130_fd_sc_hd__mux2_1_0.S 0.42059f
C698 w_12894_4504# a_13285_5437# 0
C699 a_12320_4959# VGND 0.00281f
C700 w_6570_15449# VPWR 0.08494f
C701 a_8113_13753# a_9597_13793# 0.00382f
C702 a_12976_1743# a_13105_2135# 0.00792f
C703 sky130_fd_sc_hd__inv_1_4.A VPWR 0.25987f
C704 VGND a_11958_5833# 0.1907f
C705 a_7635_5039# a_7899_5039# 0
C706 a_6885_1783# sky130_fd_sc_hd__inv_1_0.A 0.00266f
C707 w_7604_13967# a_7113_13395# 0.04664f
C708 w_11008_1688# sky130_fd_sc_hd__inv_1_0.A 0.00321f
C709 a_9875_13765# w_10872_13125# 0.09336f
C710 a_3790_1761# a_4183_1787# 0.02283f
C711 a_10088_5471# w_9180_5386# 0.01154f
C712 a_6362_1783# a_6885_1783# 0
C713 a_2706_5051# a_3229_5051# 0
C714 w_4432_13071# a_4847_14525# 0
C715 a_10771_14747# VGND 0.13243f
C716 a_3040_5051# VPWR 0
C717 sky130_fd_sc_hd__inv_1_2.A sky130_fd_sc_hd__inv_1_4.A 0
C718 a_10771_14747# a_9799_16073# 0.03093f
C719 a_9865_15329# a_9811_11277# 0.30844f
C720 a_4627_12141# a_4637_10577# 0
C721 a_5851_13769# w_5910_13141# 0.00142f
C722 a_9699_4853# A 0
C723 a_6003_11935# VPWR 0.1599f
C724 a_9465_16323# a_9809_14509# 0
C725 VGND a_6726_5409# 0.00245f
C726 sky130_fd_sc_hd__inv_1_2.VPB VPWR 0.0708f
C727 a_24962_14701# sky130_fd_sc_hd__inv_1_0.A 0.00234f
C728 a_15141_4951# a_14916_4559# 0.00559f
C729 a_9801_12841# a_9683_13793# 0
C730 a_11331_5467# a_11202_5441# 0.00758f
C731 a_11108_1773# sky130_fd_sc_hd__inv_1_0.A 0.00117f
C732 a_5765_5043# a_5903_5017# 0
C733 a_6389_13769# a_4837_16089# 0.00515f
C734 a_11243_11891# a_12075_13379# 0.19825f
C735 VPWR a_11679_15219# 0
C736 a_24241_14651# a_24234_14385# 0.13413f
C737 a_3919_2153# a_3790_1761# 0.00792f
C738 a_6003_11935# a_6281_11907# 0.11706f
C739 a_4515_11543# w_4540_10763# 0.0035f
C740 VPWR a_4045_5413# 0
C741 a_11049_14719# a_10813_13753# 0
C742 a_9599_10561# VPWR 0.36832f
C743 a_4513_14775# a_4837_16089# 0
C744 a_4915_10549# w_4540_10763# 0.0204f
C745 sky130_fd_sc_hd__inv_1_2.A sky130_fd_sc_hd__inv_1_2.VPB 0.05602f
C746 a_15309_4585# a_14916_4559# 0.02283f
C747 a_4915_10549# a_5851_13769# 0.00193f
C748 a_9801_12841# a_9725_14759# 0.00187f
C749 a_4753_16339# VGND 0.01705f
C750 w_9500_13979# a_9587_15357# 0
C751 a_4635_13809# a_4903_15345# 0.00159f
C752 a_13147_5463# A 0
C753 a_8262_5039# VPWR 0.2064f
C754 a_14916_4559# sky130_fd_sc_hd__mux2_1_0.S 0
C755 a_24152_14385# ui_in[0] 0.02237f
C756 a_9629_2033# VPWR 0.34514f
C757 a_12631_13987# a_11243_11891# 0.19153f
C758 a_9332_5445# a_7845_5295# 0
C759 a_10965_11919# w_9492_12311# 0
C760 a_10965_11919# a_11051_11919# 0.00658f
C761 a_4129_2043# a_5873_1757# 0.00412f
C762 uio_in[2] uio_in[3] 0.03102f
C763 a_24774_14701# sky130_fd_sc_hd__inv_1_0.A 0.00262f
C764 a_11230_4567# sky130_fd_sc_hd__inv_1_0.A 0
C765 a_13201_1769# a_13369_1769# 0
C766 a_4849_11293# a_6129_12927# 0
C767 a_4913_13781# VGND 0.70497f
C768 a_11359_4959# VGND 0.00292f
C769 a_9683_2143# a_9515_2143# 0
C770 a_7635_5405# a_7454_5039# 0
C771 a_4513_14775# a_4595_14775# 0.00641f
C772 a_11160_1747# VGND 0.40116f
C773 Y a_5636_5017# 0.0021f
C774 a_4183_1787# VPWR 0.17525f
C775 a_11595_5467# a_11331_5467# 0
C776 a_9865_15329# w_10748_13967# 0.07513f
C777 a_9715_16323# a_9587_15357# 0
C778 a_14946_4905# w_14736_5374# 0.02228f
C779 a_2145_2157# a_1920_1765# 0.00559f
C780 a_9699_4853# a_9671_5727# 0.00177f
C781 a_6696_2149# VGND 0.00244f
C782 ui_in[0] rst_n 0.03102f
C783 a_9877_10533# w_10868_12105# 0
C784 a_10611_5471# A 0.0073f
C785 a_9801_12841# a_10965_11919# 0
C786 a_12976_1743# w_11008_1688# 0
C787 a_9467_13091# a_9717_13091# 0.02504f
C788 a_5606_1757# a_5945_2039# 0.04737f
C789 a_6392_5409# a_5975_5299# 0.06611f
C790 a_5735_1783# VPWR 0.00115f
C791 a_4635_13809# a_4755_13107# 0
C792 a_15672_4585# a_14946_4905# 0.01208f
C793 a_4503_16339# VGND 0.28566f
C794 a_9875_13765# a_10937_12911# 0.08477f
C795 a_13385_4845# VPWR 0.37942f
C796 a_4837_16089# a_4839_12857# 0.4639f
C797 a_11202_5441# w_9180_5386# 0
C798 a_11906_13629# VPWR 0.0014f
C799 a_3010_2157# VPWR 0
C800 a_14888_5433# w_14736_5374# 0.05213f
C801 a_3919_2153# VPWR 0
C802 a_15978_5825# a_15227_5715# 0.00696f
C803 a_6885_1783# w_7324_1694# 0.25055f
C804 a_6389_13769# a_5851_13769# 0.07901f
C805 VGND a_11291_12911# 0.19423f
C806 a_14794_1765# w_12824_1684# 0.00188f
C807 sky130_fd_sc_hd__inv_1_4.A sky130_fd_sc_hd__inv_1_5.A 0.1036f
C808 w_12894_4504# sky130_fd_sc_hd__inv_1_0.A 0.00104f
C809 w_11050_5382# a_13285_5437# 0.00743f
C810 a_11289_1773# sky130_fd_sc_hd__inv_1_0.A 0
C811 a_9753_4963# A 0
C812 a_2676_2157# a_2259_2047# 0.06611f
C813 a_1868_1791# VPWR 0.08418f
C814 a_11160_1747# a_11385_1773# 0.00487f
C815 a_15672_4951# a_14297_5463# 0
C816 ui_in[0] VPWR 0.10592f
C817 Y a_2343_5051# 0.0842f
C818 VGND a_13411_5463# 0.01681f
C819 a_5069_1787# VPWR 0.06754f
C820 a_2313_2157# a_1920_1765# 0.02301f
C821 ui_in[0] sky130_fd_sc_hd__mux4_1_0.VPB 0.27045f
C822 a_7845_5295# a_8262_5039# 0.03016f
C823 a_2343_5051# a_1950_5025# 0.02283f
C824 a_9727_11527# a_9811_11277# 0.08177f
C825 a_4595_14775# a_4839_12857# 0
C826 a_4015_2153# sky130_fd_sc_hd__inv_1_0.Y 0
C827 a_11958_5833# a_11541_5723# 0.06611f
C828 a_2289_5307# w_3668_4962# 0
C829 w_9208_4512# VGND 0.28745f
C830 a_9811_11277# a_12075_13379# 0.00118f
C831 sky130_fd_sc_hd__inv_1_0.Y sky130_fd_sc_hd__inv_1_0.VPB 0.02708f
C832 VPWR a_13285_5437# 0.94532f
C833 a_17053_4938# VGND 0
C834 a_16871_4938# sky130_fd_sc_hd__mux2_1_0.A1 0.15182f
C835 a_11986_4593# a_11569_4849# 0.03016f
C836 sky130_fd_sc_hd__inv_1_2.A ui_in[0] 0.00113f
C837 a_13271_4589# VGND 0
C838 VGND w_11718_13593# 0.01919f
C839 a_7869_1779# sky130_fd_sc_hd__inv_1_0.A 0
C840 a_9671_5727# a_10611_5471# 0.13962f
C841 a_6029_5409# w_5484_4958# 0
C842 w_11718_13593# a_9799_16073# 0
C843 a_9753_4597# sky130_fd_sc_hd__inv_1_0.A 0
C844 a_7669_14003# a_7173_15235# 0.16709f
C845 a_15281_5459# w_14736_5374# 0.01092f
C846 a_11230_4567# a_11178_4593# 0.1439f
C847 a_9419_2143# a_9290_1751# 0.00792f
C848 a_14325_4589# a_15281_5825# 0
C849 a_14066_2135# a_13315_2025# 0.00696f
C850 a_6862_13645# a_4915_10549# 0
C851 a_13313_4563# VGND 0.6054f
C852 a_7424_1779# VPWR 0.07407f
C853 VGND a_6717_15235# 0.00151f
C854 a_10857_14747# a_11049_14719# 0
C855 sky130_fd_sc_hd__mux2_1_0.S w_14736_5374# 0.00355f
C856 a_9865_15329# a_9725_14759# 0.00327f
C857 a_4905_12113# VPWR 0.28921f
C858 a_10639_4597# sky130_fd_sc_hd__mux2_1_0.S 0.03363f
C859 a_9597_13793# a_10813_13753# 0
C860 a_15672_4585# a_15309_4585# 0.00985f
C861 a_23677_14335# ui_in[0] 0
C862 a_9801_12841# a_11351_13753# 0.04676f
C863 VPWR a_9717_13091# 0.31944f
C864 a_1920_1765# w_1768_1706# 0.05213f
C865 w_11532_15433# VPWR 0.08492f
C866 a_6635_15235# a_6717_15235# 0.00578f
C867 a_6087_14735# w_6756_13609# 0
C868 a_2259_2047# VGND 1.20011f
C869 a_5851_13769# a_4839_12857# 0.13074f
C870 a_4905_12113# a_6281_11907# 0.03573f
C871 a_13439_4955# w_12894_4504# 0
C872 a_4903_15345# a_5809_14763# 0.0039f
C873 a_11623_4593# a_11230_4567# 0.02283f
C874 a_11091_12911# VPWR 0
C875 Y a_3949_5413# 0
C876 ui_in[0] ui_in[1] 5.4829f
C877 a_8262_5405# a_6915_5043# 0.03325f
C878 a_7113_13395# a_5975_12927# 0
C879 sky130_fd_sc_hd__inv_1_2.A w_11532_15433# 0
C880 a_5999_1783# a_5735_1783# 0
C881 a_13439_4955# a_13271_4955# 0
C882 a_3919_1787# VGND 0
C883 a_6696_1783# sky130_fd_sc_hd__inv_1_0.A 0
C884 a_7869_2145# a_8232_2145# 0.00847f
C885 a_6029_5043# w_5484_4958# 0.01092f
C886 a_14916_4559# a_14297_5463# 0
C887 a_9465_16323# a_8113_13753# 0.0062f
C888 a_12250_2139# VPWR 0
C889 a_17125_4938# a_14946_4905# 0.00161f
C890 a_9589_12125# a_9727_11527# 0
C891 w_6756_13609# a_7113_13395# 0.03222f
C892 a_7669_14003# w_5786_13983# 0
C893 w_10748_13967# a_12075_13379# 0
C894 a_4903_15345# a_6127_13769# 0
C895 a_15227_5715# A 0.00796f
C896 a_5895_14763# a_7173_15235# 0
C897 a_4159_5303# a_5636_5017# 0.00492f
C898 a_15185_2021# VPWR 0.33214f
C899 a_11331_5833# VPWR 0
C900 a_4849_11293# w_4538_13995# 0.00123f
C901 a_14066_1769# sky130_fd_sc_hd__inv_1_0.A 0
C902 a_11499_2029# a_11916_1773# 0.03016f
C903 a_4847_14525# VGND 0.43095f
C904 a_9477_11527# a_9727_11527# 0.02504f
C905 a_9629_2033# a_9515_1777# 0
C906 a_13802_4955# w_12894_4504# 0.00139f
C907 VPWR w_9138_1692# 0.51534f
C908 a_5606_1757# VGND 0.40141f
C909 a_6862_13645# a_6389_13769# 0.24537f
C910 a_11569_4849# a_10611_5471# 0
C911 a_4576_5047# VPWR 0.20634f
C912 w_10748_13967# a_12631_13987# 0
C913 a_6635_15235# a_4847_14525# 0.17824f
C914 VGND a_11150_5467# 0.08811f
C915 a_9332_5445# A 0.00451f
C916 a_8566_1779# sky130_fd_sc_hd__inv_1_0.A 0
C917 a_6029_5043# a_6392_5043# 0.00985f
C918 a_4513_14775# w_4528_15559# 0
C919 a_4627_12141# w_4538_13995# 0
C920 a_7506_5013# a_7731_5405# 0.00559f
C921 a_5873_1757# VPWR 0.96923f
C922 sky130_fd_sc_hd__mux2_1_0.A0 a_15227_5715# 0.13856f
C923 a_10611_5471# a_11595_5833# 0.04534f
C924 VPWR a_7173_15235# 0.55471f
C925 a_9461_5837# VGND 0.00346f
C926 Y a_1950_5025# 0.08244f
C927 a_4213_5047# VPWR 0.17485f
C928 a_9461_5471# A 0
C929 a_4849_11293# a_5895_14763# 0.00121f
C930 a_5831_1783# a_5873_1757# 0
C931 a_7869_1779# w_7324_1694# 0.01092f
C932 a_12924_1769# a_13243_1743# 0.04799f
C933 a_6911_15235# a_4837_16089# 0.00241f
C934 w_4440_14739# a_4625_15373# 0.00155f
C935 a_3040_5417# a_3229_5051# 0
C936 a_9629_2033# a_9683_2143# 0.03622f
C937 a_6281_11907# a_7173_15235# 0.09936f
C938 a_12135_15219# a_9877_10533# 0.07807f
C939 a_11906_13629# a_11243_11891# 0
C940 a_4711_15373# a_4625_15373# 0.00658f
C941 a_13732_2135# VPWR 0.01969f
C942 a_7919_14003# VGND 0
C943 sky130_fd_sc_hd__inv_1_0.A VPWR 0.2927f
C944 a_5999_2149# a_6362_2149# 0.00847f
C945 a_13046_4563# VGND 0.41147f
C946 a_6087_14735# w_6570_15449# 0.06196f
C947 sky130_fd_sc_hd__inv_1_0.A sky130_fd_sc_hd__mux4_1_0.VPB 0.08268f
C948 a_6362_1783# VPWR 0.20684f
C949 a_3949_5047# a_3229_5051# 0
C950 a_11108_1773# w_11008_1688# 0.01793f
C951 a_9360_4571# w_9180_5386# 0.00104f
C952 a_17125_4938# sky130_fd_sc_hd__mux2_1_0.S 0.31816f
C953 a_2145_2157# VPWR 0
C954 a_5933_13769# VGND 0.00382f
C955 a_10450_4963# VGND 0.00221f
C956 a_7506_5013# VGND 0.40201f
C957 a_4849_11293# VPWR 0.42529f
C958 a_9865_15329# a_11351_13753# 0
C959 a_6862_13645# a_4839_12857# 0.00327f
C960 a_4849_11293# a_6944_13645# 0
C961 w_5786_13983# VPWR 0.0898f
C962 a_9332_5445# a_9671_5727# 0.04737f
C963 a_2259_2047# w_3638_1702# 0
C964 a_10569_1777# a_11916_1773# 0.08907f
C965 a_12713_13987# a_12075_13379# 0.00226f
C966 a_9801_12841# a_10771_14747# 0.21988f
C967 a_4849_11293# a_6281_11907# 0.00683f
C968 a_3790_1761# w_1768_1706# 0
C969 a_14325_4589# w_12894_4504# 0.02026f
C970 a_8596_5039# VPWR 0
C971 w_5786_13983# a_6281_11907# 0
C972 a_11049_14719# VGND 0.35053f
C973 a_8262_5039# A 0
C974 a_14297_5463# w_14736_5374# 0.25055f
C975 a_9599_10561# a_9811_11277# 0
C976 a_11049_14719# a_9799_16073# 0.29394f
C977 a_10813_13753# w_10872_13125# 0.00142f
C978 a_4627_12141# VPWR 0.38028f
C979 sky130_fd_sc_hd__inv_1_0.A ui_in[1] 0.0357f
C980 a_12481_5467# a_13018_5437# 0
C981 a_12631_13987# a_12713_13987# 0.00695f
C982 VGND a_2706_5051# 0.01359f
C983 a_15672_4585# a_14297_5463# 0
C984 a_15017_5825# VGND 0.00305f
C985 a_24962_14701# a_24774_14701# 0.10432f
C986 a_12994_4589# w_12894_4504# 0.01793f
C987 a_4627_12141# a_6281_11907# 0
C988 a_13439_4955# VPWR 0.00924f
C989 VPWR a_9557_5471# 0
C990 a_5861_5043# a_5975_5299# 0
C991 a_4903_15345# a_4913_13781# 0.1161f
C992 a_2313_2157# VPWR 0.00745f
C993 Y a_1898_5051# 0.0073f
C994 a_23731_14309# ui_in[0] 0.35239f
C995 a_4765_11293# a_4849_11293# 0.00206f
C996 a_6329_12927# VGND 0.19423f
C997 uio_oe[0] uio_oe[1] 0.03102f
C998 a_1898_5051# a_1950_5025# 0.1439f
C999 w_9500_13979# a_7173_15235# 0
C1000 a_5999_1783# a_5873_1757# 0.08094f
C1001 a_9809_14509# a_9475_14759# 0.1679f
C1002 a_11160_1747# a_11385_2139# 0.00559f
C1003 a_9280_5471# VPWR 0.07735f
C1004 a_15113_5459# VGND 0
C1005 a_5606_1757# w_3638_1702# 0
C1006 sky130_fd_sc_hd__inv_1_5.Y a_23511_14335# 0.05256f
C1007 a_7476_1753# a_7424_1779# 0.1439f
C1008 a_12976_1743# VPWR 0.29525f
C1009 a_6029_5409# VPWR 0.00962f
C1010 w_12866_5378# VGND 0.31514f
C1011 a_11499_2029# a_13243_1743# 0.00412f
C1012 a_9308_4597# sky130_fd_sc_hd__mux2_1_0.S 0
C1013 a_5554_1783# VGND 0.08664f
C1014 a_11178_4593# VPWR 0.09319f
C1015 a_15045_4951# a_14916_4559# 0.00792f
C1016 w_9392_16287# VPWR 0.16528f
C1017 a_4903_15345# a_4503_16339# 0
C1018 a_8755_1779# a_9419_1777# 0
C1019 a_7731_5039# a_6915_5043# 0
C1020 a_5584_5043# w_3668_4962# 0.00227f
C1021 a_13385_4845# A 0
C1022 a_15255_4841# a_15309_4951# 0.03622f
C1023 a_2259_2047# a_2145_1791# 0
C1024 a_5999_1783# sky130_fd_sc_hd__inv_1_0.A 0
C1025 sky130_fd_sc_hd__inv_1_0.Y a_2259_2047# 0.25757f
C1026 VPWR w_7324_1694# 0.51443f
C1027 ui_in[0] a_23511_14701# 0.05408f
C1028 a_15113_5825# VGND 0.00231f
C1029 a_13313_4563# a_13411_5829# 0
C1030 a_9725_14759# a_9587_15357# 0
C1031 a_9875_13765# w_10868_12105# 0
C1032 a_13802_4955# VPWR 0.02429f
C1033 a_9877_10533# w_9404_11491# 0
C1034 a_11623_4959# a_10639_4597# 0.04534f
C1035 a_6362_1783# a_5999_1783# 0.00985f
C1036 sky130_fd_sc_hd__inv_1_2.A w_9392_16287# 0
C1037 a_9811_11277# a_11906_13629# 0
C1038 Y a_4159_5303# 0.00305f
C1039 w_1768_1706# VPWR 0.51727f
C1040 a_13175_4589# a_13439_4589# 0
C1041 a_9589_12125# a_9599_10561# 0
C1042 a_9585_4597# a_9699_4853# 0
C1043 a_13357_5719# a_13385_4845# 0.00177f
C1044 a_9875_13765# a_9475_14759# 0
C1045 a_11623_4593# VPWR 0.17434f
C1046 a_15309_4951# VGND 0.00129f
C1047 sky130_fd_sc_hd__inv_1_0.Y a_3919_1787# 0
C1048 a_6726_5043# VPWR 0
C1049 uio_out[3] uio_out[4] 0.03102f
C1050 a_3199_1791# a_2259_2047# 0.13962f
C1051 ui_in[0] A 0.07335f
C1052 a_13313_4563# w_11078_4508# 0.00743f
C1053 a_7845_5295# a_8596_5039# 0.00682f
C1054 w_9490_15543# VGND 0.11947f
C1055 w_4440_14739# VPWR 0.16205f
C1056 a_6029_5043# VPWR 0.17685f
C1057 a_9801_12841# a_11291_12911# 0.08252f
C1058 a_6885_1783# a_7869_1779# 0.08312f
C1059 a_9865_15329# a_11597_15219# 0
C1060 w_9490_15543# a_9799_16073# 0.00251f
C1061 a_9477_11527# a_9599_10561# 0.00144f
C1062 a_10046_2143# a_8755_1779# 0.03325f
C1063 a_4721_13809# a_4839_12857# 0
C1064 a_15227_5715# w_14764_4500# 0
C1065 a_4711_15373# VPWR 0.00333f
C1066 a_10813_13753# a_10937_12911# 0
C1067 a_9867_12097# w_10872_13125# 0
C1068 a_8596_5405# sky130_fd_sc_hd__mux2_1_0.S 0
C1069 A a_13285_5437# 0.00473f
C1070 a_3199_1791# a_3919_1787# 0
C1071 VPWR w_3668_4962# 0.51523f
C1072 VGND w_9402_14723# 0.07437f
C1073 w_9402_14723# a_9799_16073# 0
C1074 a_4015_1787# VGND 0
C1075 a_4915_10549# a_9877_10533# 0.00316f
C1076 a_15255_4841# a_14946_4905# 1.1874f
C1077 a_6392_5043# w_5484_4958# 0.01154f
C1078 a_11351_13753# a_12075_13379# 0.06159f
C1079 a_5606_1757# sky130_fd_sc_hd__inv_1_0.Y 0.0021f
C1080 a_2259_2047# a_2313_1791# 0.00386f
C1081 a_4755_12857# a_4849_11293# 0
C1082 a_9865_15329# a_10771_14747# 0.0039f
C1083 w_11050_5382# a_11958_5467# 0.01154f
C1084 a_13105_2135# VPWR 0
C1085 a_13357_5719# a_13285_5437# 0.21146f
C1086 Y VPB 0.02708f
C1087 a_9683_2143# w_9138_1692# 0
C1088 a_10422_5471# VGND 0
C1089 a_7635_5039# a_6915_5043# 0
C1090 a_10569_1777# a_13243_1743# 0
C1091 a_9515_1777# sky130_fd_sc_hd__inv_1_0.A 0
C1092 a_7845_5295# a_9280_5471# 0
C1093 a_4183_2153# VGND 0.20098f
C1094 a_2175_5051# a_2289_5307# 0
C1095 a_9801_12841# w_11718_13593# 0.00515f
C1096 a_10116_4597# sky130_fd_sc_hd__inv_1_0.A 0
C1097 a_8232_1779# sky130_fd_sc_hd__inv_1_0.A 0
C1098 a_9597_13793# VGND 0.24546f
C1099 a_14946_4905# VGND 0.17745f
C1100 a_12881_13987# a_9877_10533# 0
C1101 a_11351_13753# a_12631_13987# 0.00196f
C1102 a_9811_11277# a_9717_13091# 0
C1103 a_11958_5467# VPWR 0.20396f
C1104 a_4915_10549# a_9475_14759# 0
C1105 a_7476_1753# sky130_fd_sc_hd__inv_1_0.A 0.00206f
C1106 a_24318_14385# ui_in[0] 0.04767f
C1107 a_10380_2143# VPWR 0
C1108 a_14325_4589# VPWR 1.12038f
C1109 a_9811_11277# a_11091_12911# 0
C1110 a_15602_2131# a_15185_2021# 0.06611f
C1111 sky130_fd_sc_hd__inv_1_5.Y sky130_fd_sc_hd__inv_1_5.VPB 0.04452f
C1112 a_9290_1751# a_9515_2143# 0.00559f
C1113 a_14888_5433# VGND 0.40147f
C1114 a_9683_2143# sky130_fd_sc_hd__inv_1_0.A 0
C1115 uo_out[3] uo_out[2] 0.03102f
C1116 a_9725_5837# w_9180_5386# 0
C1117 a_23731_14309# sky130_fd_sc_hd__inv_1_0.A 0
C1118 a_11331_5833# A 0
C1119 a_15281_5825# VPWR 0.00604f
C1120 a_5861_5043# a_5636_5017# 0.00487f
C1121 a_15255_4841# a_15141_4951# 0
C1122 a_5975_12927# a_5809_14763# 0
C1123 a_4637_10577# VPWR 0.36832f
C1124 w_9394_13055# a_9597_13793# 0.00101f
C1125 a_5099_5047# a_5636_5017# 0
C1126 a_4837_16089# VGND 0.68517f
C1127 a_12994_4589# VPWR 0.07511f
C1128 a_5554_1783# w_3638_1702# 0.00227f
C1129 a_10422_5837# VGND 0.00262f
C1130 a_9809_14509# a_9673_15357# 0
C1131 a_4903_15345# a_4847_14525# 0.15229f
C1132 w_9502_10747# a_9877_10533# 0.0204f
C1133 a_15255_4841# a_15309_4585# 0.00386f
C1134 w_12866_5378# a_11541_5723# 0
C1135 a_15255_4841# a_15281_5459# 0
C1136 a_10611_5471# a_11958_5833# 0.03325f
C1137 w_9392_16287# a_9715_16323# 0.01327f
C1138 a_4837_16089# a_6635_15235# 0.232f
C1139 a_12135_15219# a_11767_15219# 0
C1140 a_10639_4597# a_11202_5441# 0
C1141 a_7701_2145# VPWR 0
C1142 a_24774_14701# a_24152_14385# 0
C1143 a_15644_5825# a_15281_5825# 0.00847f
C1144 a_6389_13769# a_6021_13769# 0
C1145 w_12866_5378# a_12966_5463# 0.01793f
C1146 a_9867_12097# a_10937_12911# 0
C1147 a_14946_4905# a_17125_5265# 0
C1148 ua[5] w_11008_1688# 0
C1149 a_15255_4841# sky130_fd_sc_hd__mux2_1_0.S 0.00102f
C1150 a_14864_4585# a_13385_4845# 0
C1151 a_13046_4563# w_11078_4508# 0
C1152 a_2289_5307# VPWR 0.34431f
C1153 a_14946_4905# a_17346_5265# 0
C1154 a_5735_2149# VGND 0.00305f
C1155 a_6885_1783# VPWR 1.0518f
C1156 a_9809_14509# a_12135_15219# 0
C1157 w_11008_1688# VPWR 0.51509f
C1158 a_15309_4585# VGND 0
C1159 a_9589_12125# a_9717_13091# 0
C1160 a_15602_2131# sky130_fd_sc_hd__inv_1_0.A 0.00187f
C1161 a_4129_2043# a_4880_1787# 0.00682f
C1162 a_15281_5459# VGND 0.01492f
C1163 a_4595_14775# VGND 0.00172f
C1164 a_5606_1757# a_5999_2149# 0.02301f
C1165 a_12320_4593# sky130_fd_sc_hd__inv_1_0.A 0
C1166 a_6087_14735# a_7173_15235# 0.00425f
C1167 a_9585_4963# VPWR 0
C1168 a_11597_15219# a_12075_13379# 0
C1169 a_8113_13753# a_9475_14759# 0.0055f
C1170 sky130_fd_sc_hd__mux2_1_0.S VGND 1.9195f
C1171 a_3790_1761# a_4129_2043# 0.04737f
C1172 a_11108_1773# ua[5] 0
C1173 a_9557_5837# VPWR 0
C1174 a_13243_5463# a_13285_5437# 0
C1175 w_5484_4958# a_5584_5043# 0.01793f
C1176 a_4546_1787# VGND 0.01333f
C1177 a_8566_2145# sky130_fd_sc_hd__inv_1_0.A 0
C1178 a_11916_1773# VGND 0.01327f
C1179 w_7354_4954# VPWR 0.51208f
C1180 sky130_fd_sc_hd__inv_1_0.A A 0.91673f
C1181 a_9238_1777# a_8755_1779# 0.07352f
C1182 a_4505_13107# w_5910_13141# 0
C1183 a_24962_14701# VPWR 0.21151f
C1184 a_7899_5039# VGND 0.0165f
C1185 uo_out[3] uo_out[4] 0.03102f
C1186 a_24962_14701# sky130_fd_sc_hd__mux4_1_0.VPB 0.07712f
C1187 a_9809_14509# a_11767_15219# 0.00624f
C1188 a_11108_1773# VPWR 0.07418f
C1189 a_11595_5467# a_10639_4597# 0
C1190 a_13315_2025# sky130_fd_sc_hd__inv_1_0.A 0.00291f
C1191 a_13315_2025# a_13732_2135# 0.06611f
C1192 a_13774_5463# a_13285_5437# 0.08907f
C1193 w_4430_16303# a_4625_15373# 0
C1194 a_8232_1779# w_7324_1694# 0.01154f
C1195 a_7113_13395# a_7173_15235# 0.36868f
C1196 sky130_fd_sc_hd__inv_1_0.Y a_5554_1783# 0.0012f
C1197 a_5933_13769# a_4903_15345# 0.0035f
C1198 a_4515_11543# a_4505_13107# 0.00102f
C1199 w_11050_5382# a_11230_4567# 0.00104f
C1200 a_4505_13107# w_4442_11507# 0
C1201 a_6003_11935# a_6089_11935# 0.00658f
C1202 VGND w_4540_10763# 0.12086f
C1203 a_6129_12927# VPWR 0
C1204 a_13385_4845# w_14764_4500# 0
C1205 a_12439_1773# a_12924_1769# 0.02709f
C1206 a_5851_13769# VGND 0.15513f
C1207 a_4183_2153# w_3638_1702# 0
C1208 a_7476_1753# w_7324_1694# 0.05213f
C1209 w_4538_13995# a_4625_15373# 0
C1210 w_12866_5378# a_13411_5829# 0
C1211 a_6087_14735# a_4849_11293# 0.00179f
C1212 a_9699_4853# w_9208_4512# 0.10454f
C1213 a_6021_13769# a_4839_12857# 0
C1214 a_6087_14735# w_5786_13983# 0
C1215 sky130_fd_sc_hd__inv_1_2.Y w_5712_14949# 0
C1216 a_11160_1747# a_11553_2139# 0.02301f
C1217 w_4530_12327# a_4505_13107# 0.0035f
C1218 a_11986_4593# a_13313_4563# 0
C1219 a_1920_1765# VPWR 0.30549f
C1220 a_24774_14701# VPWR 0.0823f
C1221 a_8596_5039# A 0
C1222 a_11824_13629# VPWR 0.09661f
C1223 a_24774_14701# sky130_fd_sc_hd__mux4_1_0.VPB 0.14223f
C1224 VGND a_3040_5417# 0.00244f
C1225 a_11230_4567# VPWR 0.31788f
C1226 a_4910_5047# VPWR 0
C1227 w_5484_4958# VPWR 0.5153f
C1228 a_4513_14775# a_4763_14775# 0.02504f
C1229 a_3768_5047# w_3668_4962# 0.01793f
C1230 a_13147_5463# a_13411_5463# 0
C1231 a_10046_1777# a_8755_1779# 0.08907f
C1232 a_24962_14701# ui_in[1] 0.02448f
C1233 a_15644_5459# w_14736_5374# 0.01154f
C1234 a_4915_10549# w_5906_12121# 0
C1235 w_10872_13125# VGND 0.02002f
C1236 a_24318_14385# sky130_fd_sc_hd__inv_1_0.A 0.05111f
C1237 w_10872_13125# a_9799_16073# 0
C1238 ua[4] VPWR 0.00186f
C1239 a_3949_5047# VGND 0
C1240 a_4849_11293# a_7113_13395# 0.00118f
C1241 a_13439_4955# A 0
C1242 a_9557_5471# A 0
C1243 a_4129_2043# VPWR 0.34563f
C1244 a_12292_5833# A 0
C1245 a_9809_14509# a_9875_13765# 0.0012f
C1246 a_4849_11293# a_4587_13107# 0
C1247 w_5786_13983# a_7113_13395# 0
C1248 a_9801_12841# a_11049_14719# 0.02474f
C1249 a_13732_1769# VGND 0.01325f
C1250 sky130_fd_sc_hd__inv_1_0.Y a_4015_1787# 0
C1251 a_10380_1777# a_9629_2033# 0.00682f
C1252 a_7845_5295# w_7354_4954# 0.10454f
C1253 a_9280_5471# A 0.00331f
C1254 a_6029_5409# A 0
C1255 a_14108_5463# VPWR 0
C1256 a_16006_4951# sky130_fd_sc_hd__mux2_1_0.A1 0
C1257 a_4503_16339# a_4753_16089# 0.00723f
C1258 a_6392_5043# VPWR 0.20634f
C1259 a_11178_4593# A 0
C1260 a_6389_13769# sky130_fd_sc_hd__inv_1_2.Y 0
C1261 a_4913_13781# a_5975_12927# 0.08477f
C1262 a_8113_13753# sky130_fd_sc_hd__inv_1_2.Y 0.03523f
C1263 w_12894_4504# VPWR 0.52921f
C1264 a_4513_14775# a_4505_13107# 0
C1265 a_24774_14701# ui_in[1] 0.02507f
C1266 a_11289_1773# VPWR 0.00117f
C1267 a_4183_2153# sky130_fd_sc_hd__inv_1_0.Y 0
C1268 a_13315_2025# a_12976_1743# 0.04737f
C1269 a_11986_4959# VPWR 0.02086f
C1270 a_11331_5833# a_11595_5833# 0
C1271 a_3199_1791# a_4015_1787# 0
C1272 a_13369_2135# a_13243_1743# 0.04534f
C1273 VPWR a_4625_15373# 0.38724f
C1274 a_13802_4955# A 0
C1275 a_13271_4955# VPWR 0
C1276 Y a_5861_5043# 0
C1277 a_4763_14775# a_4839_12857# 0.00187f
C1278 a_2706_5051# w_1798_4966# 0.01154f
C1279 a_2259_2047# a_2676_1791# 0.03016f
C1280 a_11291_12911# a_12075_13379# 0
C1281 a_9465_16323# VGND 0.28565f
C1282 a_9465_16323# a_9799_16073# 0.16891f
C1283 a_11427_5833# a_11202_5441# 0.00559f
C1284 a_5099_5047# Y 0
C1285 a_13732_1769# a_14255_1769# 0
C1286 a_9629_2033# a_9290_1751# 0.04737f
C1287 a_15255_4841# a_14297_5463# 0
C1288 a_12439_1773# a_11499_2029# 0.12975f
C1289 a_6726_5043# A 0
C1290 a_3199_1791# a_4183_2153# 0.04534f
C1291 a_15255_4841# a_16871_4938# 0
C1292 a_12135_15219# a_12881_13987# 0
C1293 a_4546_1787# w_3638_1702# 0.01154f
C1294 a_11906_13629# a_11351_13753# 0.00183f
C1295 a_10813_13753# a_9877_10533# 0.00193f
C1296 a_9671_5727# a_9557_5471# 0
C1297 a_6029_5043# A 0
C1298 a_7869_1779# VPWR 0.17565f
C1299 a_13243_1743# VGND 0.60976f
C1300 a_9753_4597# VPWR 0.26479f
C1301 sky130_fd_sc_hd__mux2_1_0.S a_11541_5723# 0
C1302 a_9809_14509# a_4915_10549# 0
C1303 a_9753_4963# w_9208_4512# 0
C1304 a_11569_4849# sky130_fd_sc_hd__inv_1_0.A 0
C1305 a_14864_4585# sky130_fd_sc_hd__inv_1_0.A 0
C1306 ua[6] w_7324_1694# 0
C1307 a_14297_5463# VGND 0.67503f
C1308 a_6862_13645# VGND 0.13594f
C1309 a_3768_5047# a_2289_5307# 0
C1310 a_7506_5013# a_7635_5405# 0.00792f
C1311 a_16871_4938# VGND 0.1106f
C1312 a_6805_15235# a_7173_15235# 0
C1313 a_14946_4905# a_15017_5459# 0
C1314 a_11160_1747# a_11553_1773# 0.02283f
C1315 VGND a_10937_12911# 0.14511f
C1316 VGND w_4528_15559# 0.11947f
C1317 a_7476_1753# a_7701_2145# 0.00559f
C1318 a_10937_12911# a_9799_16073# 0
C1319 a_3949_5047# a_3820_5021# 0.00758f
C1320 a_7669_14003# VPWR 0.082f
C1321 a_10813_13753# w_10868_12105# 0
C1322 w_11718_13593# a_12075_13379# 0.03222f
C1323 a_11089_13753# VPWR 0.0014f
C1324 w_4430_16303# VPWR 0.16502f
C1325 a_11597_15219# a_11679_15219# 0.00578f
C1326 a_6862_13645# a_6635_15235# 0
C1327 a_8232_1779# a_6885_1783# 0.08907f
C1328 a_4839_12857# a_4505_13107# 0.16952f
C1329 a_8113_13753# a_12135_15219# 0.002f
C1330 a_9467_13091# VPWR 0.38927f
C1331 a_24152_14385# VPWR 0.00352f
C1332 a_7669_14003# a_6281_11907# 0.19153f
C1333 a_4880_1787# VPWR 0
C1334 a_14888_5433# a_15017_5459# 0.00758f
C1335 a_4905_12113# a_6089_11935# 0
C1336 a_9801_12841# w_9402_14723# 0.00408f
C1337 a_24152_14385# sky130_fd_sc_hd__mux4_1_0.VPB 0.00146f
C1338 a_9597_13793# w_9492_12311# 0
C1339 a_7476_1753# a_6885_1783# 0.11887f
C1340 w_4538_13995# VPWR 0.17926f
C1341 a_14255_1769# a_13243_1743# 0
C1342 a_5735_2149# sky130_fd_sc_hd__inv_1_0.Y 0
C1343 a_2289_5307# a_2343_5417# 0.03622f
C1344 a_9875_13765# a_4915_10549# 0.00401f
C1345 sky130_fd_sc_hd__inv_1_5.Y a_24407_14651# 0
C1346 a_3790_1761# VPWR 0.29465f
C1347 a_7899_5405# a_7731_5405# 0
C1348 Y a_3229_5051# 0.00475f
C1349 a_6696_1783# VPWR 0
C1350 a_2175_5051# VPWR 0.00105f
C1351 a_7815_2035# a_8232_2145# 0.06611f
C1352 a_13732_2135# w_12824_1684# 0.00139f
C1353 w_12824_1684# sky130_fd_sc_hd__inv_1_0.A 0.00315f
C1354 sky130_fd_sc_hd__inv_1_5.Y sky130_fd_sc_hd__inv_1_3.VPB 0.07239f
C1355 w_11718_13593# a_12631_13987# 0
C1356 a_9699_4853# a_10450_4963# 0.00696f
C1357 a_11958_5467# A 0
C1358 a_9715_16073# VGND 0.00773f
C1359 VGND a_5975_5299# 1.20008f
C1360 a_9715_16073# a_9799_16073# 0.00234f
C1361 w_9394_13055# a_10937_12911# 0
C1362 a_9865_15329# a_11049_14719# 0
C1363 sky130_fd_sc_hd__inv_1_0.Y a_4546_1787# 0
C1364 a_14325_4589# A 0
C1365 w_14764_4500# sky130_fd_sc_hd__inv_1_0.A 0.00111f
C1366 w_5906_12121# a_4839_12857# 0.00131f
C1367 a_5584_5043# VPWR 0.07434f
C1368 a_15672_4951# sky130_fd_sc_hd__mux2_1_0.A1 0
C1369 a_10611_5471# a_11150_5467# 0.0725f
C1370 a_14066_1769# VPWR 0
C1371 a_11427_5467# VGND 0
C1372 w_12566_13951# a_9877_10533# 0.0566f
C1373 a_9801_12841# a_9597_13793# 0.00246f
C1374 a_11623_4959# VGND 0.19557f
C1375 a_15141_4585# sky130_fd_sc_hd__inv_1_0.A 0
C1376 a_4915_10549# w_9404_11491# 0.00173f
C1377 a_9809_14509# a_8113_13753# 0.30331f
C1378 a_5895_14763# VPWR 0
C1379 a_11243_11891# a_11824_13629# 0.00248f
C1380 a_15281_5825# A 0.00135f
C1381 a_9725_5471# a_10088_5471# 0.00985f
C1382 a_10116_4963# VGND 0.1833f
C1383 a_4903_15345# a_4837_16089# 0.50561f
C1384 a_24962_14701# a_23731_14309# 0
C1385 a_12994_4589# A 0
C1386 a_3199_1791# a_4546_1787# 0.08907f
C1387 a_4635_13809# a_4849_11293# 0.00317f
C1388 a_9867_12097# a_9877_10533# 0.0298f
C1389 a_6029_5043# a_5765_5043# 0
C1390 a_8566_1779# VPWR 0
C1391 a_4213_5047# a_4045_5047# 0
C1392 a_15281_5459# a_15017_5459# 0
C1393 a_4635_13809# w_5786_13983# 0
C1394 w_11050_5382# VPWR 0.51381f
C1395 a_5945_2039# w_5454_1698# 0.10454f
C1396 a_2079_5051# a_2343_5051# 0
C1397 a_24152_14385# ui_in[1] 0.03464f
C1398 a_7899_5405# VGND 0.20211f
C1399 a_2259_2047# a_3010_1791# 0.00682f
C1400 a_6003_11935# a_4913_13781# 0
C1401 w_11078_4508# sky130_fd_sc_hd__mux2_1_0.S 0.00114f
C1402 VGND a_10088_5471# 0.10448f
C1403 ua[5] VPWR 0.00178f
C1404 a_12250_1773# a_11499_2029# 0.00682f
C1405 a_4627_12141# a_4635_13809# 0
C1406 a_4515_11543# w_4442_11507# 0.06993f
C1407 a_13105_1769# VGND 0
C1408 a_4915_10549# a_4515_11543# 0
C1409 a_4915_10549# w_4442_11507# 0
C1410 a_2049_2157# VGND 0.00311f
C1411 a_9867_12097# w_10868_12105# 0.08119f
C1412 a_5099_5047# a_4159_5303# 0.12975f
C1413 a_4721_13809# VGND 0.00661f
C1414 VPWR sky130_fd_sc_hd__mux4_1_0.VPB 0.22983f
C1415 a_7669_14003# w_9500_13979# 0
C1416 a_6944_13645# VPWR 0.0014f
C1417 a_4903_15345# a_4595_14775# 0
C1418 a_9332_5445# w_9208_4512# 0
C1419 a_24774_14701# a_23731_14309# 0.00253f
C1420 a_9585_4963# A 0
C1421 a_11623_4593# a_11569_4849# 0.00386f
C1422 a_5831_1783# VPWR 0
C1423 w_9500_13979# a_9467_13091# 0
C1424 a_14946_4905# sky130_fd_sc_hd__mux2_1_0.VPB 0.00424f
C1425 a_13201_2135# sky130_fd_sc_hd__inv_1_0.A 0
C1426 a_9557_5837# A 0
C1427 w_4530_12327# a_4515_11543# 0
C1428 w_7354_4954# A 0.00328f
C1429 a_6281_11907# VPWR 0.2162f
C1430 w_6756_13609# a_4847_14525# 0
C1431 a_6281_11907# a_6944_13645# 0
C1432 a_7869_2145# a_7605_2145# 0
C1433 a_5831_2149# VPWR 0
C1434 sky130_fd_sc_hd__inv_1_2.A VPWR 0.93097f
C1435 a_12976_1743# w_12824_1684# 0.05213f
C1436 sky130_fd_sc_hd__inv_1_2.A sky130_fd_sc_hd__mux4_1_0.VPB 0.08143f
C1437 a_14916_4559# sky130_fd_sc_hd__mux2_1_0.A1 0
C1438 a_15644_5825# VPWR 0.01852f
C1439 a_11160_1747# a_9629_2033# 0.00446f
C1440 a_3738_1787# VGND 0.08661f
C1441 a_5735_2149# a_5999_2149# 0
C1442 a_9683_1777# a_8755_1779# 0.08124f
C1443 a_9467_13091# a_9549_13091# 0.00641f
C1444 a_9865_15329# w_9490_15543# 0.01828f
C1445 ui_in[3] ui_in[2] 0.03102f
C1446 a_13802_4589# a_13313_4563# 0.08907f
C1447 a_13369_1769# sky130_fd_sc_hd__inv_1_0.A 0
C1448 w_7604_13967# a_9597_13793# 0
C1449 a_5765_5409# a_5636_5017# 0.00792f
C1450 a_23677_14335# VPWR 0
C1451 a_9290_1751# w_9138_1692# 0.05213f
C1452 a_4903_15345# a_5851_13769# 0.16764f
C1453 a_4765_11293# VPWR 0.00377f
C1454 a_9865_15329# w_9402_14723# 0.00599f
C1455 a_12809_13987# VPWR 0
C1456 a_10380_1777# sky130_fd_sc_hd__inv_1_0.A 0
C1457 a_10088_5837# w_9180_5386# 0.00139f
C1458 a_4849_11293# a_6089_11935# 0
C1459 a_13018_5437# VGND 0.42749f
C1460 w_11532_15433# a_11597_15219# 0.08205f
C1461 a_9685_10561# a_9877_10533# 0
C1462 a_11873_15219# VPWR 0
C1463 VPWR ui_in[1] 0.40159f
C1464 a_5809_14763# a_7173_15235# 0
C1465 a_9683_1777# a_9419_1777# 0
C1466 ui_in[1] sky130_fd_sc_hd__mux4_1_0.VPB 0.35053f
C1467 a_8232_1779# a_7869_1779# 0.00985f
C1468 VPWR a_4585_16339# 0.0251f
C1469 a_24774_14701# A 0
C1470 a_10116_4597# a_9753_4597# 0.00985f
C1471 a_10569_1777# a_8755_1779# 0
C1472 a_4159_5303# a_3229_5051# 0.21188f
C1473 a_11230_4567# A 0
C1474 a_6389_13769# a_4915_10549# 0.00254f
C1475 w_5484_4958# A 0.00188f
C1476 a_24407_14651# a_24234_14385# 0.00222f
C1477 a_8113_13753# a_4915_10549# 0.13594f
C1478 a_4915_10549# w_9502_10747# 0.00202f
C1479 a_4635_13809# w_4440_14739# 0
C1480 w_7604_13967# a_4837_16089# 0
C1481 sky130_fd_sc_hd__inv_1_2.A ui_in[1] 0.00242f
C1482 a_11202_5441# VGND 0.40461f
C1483 a_7476_1753# a_7869_1779# 0.02283f
C1484 a_9811_11277# a_11824_13629# 0
C1485 a_9557_5837# a_9671_5727# 0
C1486 a_9865_15329# a_9597_13793# 0.00159f
C1487 a_13201_1769# a_13243_1743# 0
C1488 VGND a_5636_5017# 0.40145f
C1489 VGND a_23511_14335# 0.23646f
C1490 w_4432_13071# a_4505_13107# 0.06993f
C1491 a_5873_1757# sky130_fd_sc_hd__inv_1_0.VPB 0
C1492 a_11019_12911# VPWR 0
C1493 a_14864_4585# a_14325_4589# 0.0725f
C1494 a_9290_1751# sky130_fd_sc_hd__inv_1_0.A 0.00208f
C1495 a_12135_15219# a_10813_13753# 0
C1496 a_4513_14775# w_5712_14949# 0
C1497 a_7845_5295# VPWR 0.34676f
C1498 a_9360_4571# a_9308_4597# 0.1439f
C1499 sky130_fd_sc_hd__mux2_1_0.VPB sky130_fd_sc_hd__mux2_1_0.S 0.17704f
C1500 a_4597_11543# a_4515_11543# 0.00641f
C1501 a_11427_5467# a_11541_5723# 0
C1502 a_17339_4938# VPWR 0.00182f
C1503 a_2079_5051# a_1950_5025# 0.00758f
C1504 clk rst_n 0.03102f
C1505 a_13201_2135# a_12976_1743# 0.00559f
C1506 w_9500_13979# VPWR 0.17935f
C1507 w_14694_1680# a_15602_1765# 0.01154f
C1508 uio_oe[5] uio_oe[4] 0.03102f
C1509 a_8232_2145# VGND 0.18643f
C1510 a_5999_1783# VPWR 0.17398f
C1511 a_14108_5463# A 0
C1512 a_9559_11527# VPWR 0.02511f
C1513 a_4849_11293# a_5809_14763# 0.10553f
C1514 a_9801_12841# w_10872_13125# 0.05199f
C1515 a_6392_5043# A 0
C1516 sky130_fd_sc_hd__inv_1_0.A sky130_fd_sc_hd__inv_1_0.VPB 0.05211f
C1517 a_11569_4849# a_12994_4589# 0
C1518 a_7454_5039# w_7354_4954# 0.01793f
C1519 a_6362_2149# a_5873_1757# 0.03325f
C1520 w_6570_15449# a_4847_14525# 0.07233f
C1521 w_5786_13983# a_5809_14763# 0
C1522 a_4839_12857# w_5910_13141# 0.05199f
C1523 w_5454_1698# VGND 0.29362f
C1524 a_9332_5445# a_9461_5837# 0.00792f
C1525 a_5999_1783# a_5831_1783# 0
C1526 VPWR a_9549_13091# 0.02512f
C1527 w_12894_4504# A 0
C1528 a_9717_12841# a_9467_13091# 0.00723f
C1529 a_9585_4597# sky130_fd_sc_hd__inv_1_0.A 0
C1530 sky130_fd_sc_hd__inv_1_5.A VPWR 0.262f
C1531 a_11986_4959# A 0
C1532 a_6329_12927# a_5975_12927# 0.09582f
C1533 a_13369_1769# a_12976_1743# 0.02283f
C1534 a_13385_4845# a_13411_5463# 0
C1535 a_8755_1779# a_7815_2035# 0.13781f
C1536 a_4713_12141# VGND 0.00662f
C1537 a_24774_14701# a_24318_14385# 0.01242f
C1538 a_13357_5719# a_14108_5463# 0.00682f
C1539 a_9360_4571# a_9489_4963# 0.00792f
C1540 a_11595_5467# VGND 0.01545f
C1541 a_13271_4955# A 0
C1542 a_4913_13781# a_4905_12113# 0.00627f
C1543 a_4849_11293# a_6127_13769# 0
C1544 a_5861_5409# a_5975_5299# 0
C1545 a_9809_14509# a_10813_13753# 0
C1546 a_4755_12857# VPWR 0.00415f
C1547 a_6362_2149# sky130_fd_sc_hd__inv_1_0.A 0
C1548 a_24152_14385# a_23731_14309# 0.01881f
C1549 a_4515_11543# a_4839_12857# 0
C1550 a_13175_4955# VGND 0.00329f
C1551 a_14297_5463# a_15017_5459# 0
C1552 a_9715_16323# VPWR 0.32305f
C1553 a_4839_12857# w_4442_11507# 0
C1554 VGND a_2343_5051# 0.01592f
C1555 sky130_fd_sc_hd__inv_1_2.A sky130_fd_sc_hd__inv_1_5.A 0
C1556 a_4915_10549# a_4839_12857# 0.00243f
C1557 a_13357_5719# w_12894_4504# 0
C1558 w_6756_13609# a_6329_12927# 0.04962f
C1559 VPWR a_4763_14525# 0.00474f
C1560 a_13271_4589# a_13385_4845# 0
C1561 a_14325_4589# w_14764_4500# 0.25055f
C1562 uio_in[1] uio_in[2] 0.03102f
C1563 a_4839_12857# w_5712_14949# 0.08813f
C1564 sky130_fd_sc_hd__inv_1_5.Y a_24234_14385# 0
C1565 a_15672_4585# sky130_fd_sc_hd__mux2_1_0.A1 0
C1566 a_3738_1787# w_3638_1702# 0.01793f
C1567 a_13313_4563# a_13385_4845# 0.21146f
C1568 w_7604_13967# a_5851_13769# 0
C1569 a_15141_4585# a_14325_4589# 0
C1570 VGND a_13243_5829# 0.00268f
C1571 a_9332_5445# a_7506_5013# 0
C1572 VGND a_9877_10533# 0.9946f
C1573 a_9877_10533# a_9799_16073# 0.01618f
C1574 a_10895_13753# VPWR 0
C1575 a_7454_5039# w_5484_4958# 0.00188f
C1576 a_12509_4593# VGND 0.06513f
C1577 a_6862_13645# a_4903_15345# 0
C1578 a_12135_15219# w_12566_13951# 0.11864f
C1579 a_11243_11891# VPWR 0.21318f
C1580 a_4183_1787# a_3919_1787# 0
C1581 a_13411_5463# a_13285_5437# 0.08094f
C1582 a_9875_13765# a_10813_13753# 0.0094f
C1583 a_4915_10549# a_4723_10577# 0
C1584 a_3768_5047# VPWR 0.07396f
C1585 a_9515_1777# VPWR 0
C1586 a_4903_15345# w_4528_15559# 0.01828f
C1587 a_3010_2157# a_2259_2047# 0.00696f
C1588 a_6021_13769# VGND 0.00475f
C1589 a_9699_4853# sky130_fd_sc_hd__mux2_1_0.S 0
C1590 w_10674_14933# VPWR 0.07858f
C1591 a_10116_4597# VPWR 0.30078f
C1592 a_15644_5459# VGND 0.01334f
C1593 a_8232_1779# VPWR 0.20639f
C1594 a_7869_2145# a_7815_2035# 0.03622f
C1595 a_15045_4585# sky130_fd_sc_hd__inv_1_0.A 0
C1596 sky130_fd_sc_hd__inv_1_2.A a_11243_11891# 0.00295f
C1597 a_12439_1773# VGND 0.06377f
C1598 VGND w_10868_12105# 0.02048f
C1599 a_24152_14385# A 0.01336f
C1600 w_10868_12105# a_9799_16073# 0
C1601 a_9811_11277# a_11089_13753# 0
C1602 a_4910_5413# VPWR 0
C1603 a_15113_5459# a_15227_5715# 0
C1604 a_10983_13753# VPWR 0
C1605 VGND a_6915_5043# 0.68138f
C1606 VGND a_3949_5413# 0.00305f
C1607 a_7476_1753# VPWR 0.29442f
C1608 a_11623_4959# w_11078_4508# 0
C1609 a_9290_1751# w_7324_1694# 0
C1610 a_9811_11277# a_9467_13091# 0.00376f
C1611 a_2049_2157# sky130_fd_sc_hd__inv_1_0.Y 0
C1612 a_14916_4559# w_14736_5374# 0.00104f
C1613 sky130_fd_sc_hd__inv_1_5.VPB VGND 0.01751f
C1614 a_13018_5437# a_11541_5723# 0.00492f
C1615 a_11160_1747# w_9138_1692# 0
C1616 VGND a_9475_14759# 0.29736f
C1617 a_9801_12841# a_10937_12911# 0.30276f
C1618 a_14136_4955# VGND 0.00215f
C1619 a_9475_14759# a_9799_16073# 0
C1620 a_13313_4563# a_13285_5437# 0.00249f
C1621 a_2343_5417# VPWR 0.00857f
C1622 a_10422_5837# a_10611_5471# 0
C1623 a_9717_12841# VPWR 0.00415f
C1624 a_6389_13769# a_4839_12857# 0.04676f
C1625 a_13018_5437# a_12966_5463# 0.1439f
C1626 a_11230_4567# a_11569_4849# 0.04737f
C1627 a_9683_2143# VPWR 0.00879f
C1628 a_11331_5467# VGND 0
C1629 a_4513_14775# a_4839_12857# 0.00442f
C1630 w_4440_14739# a_5809_14763# 0
C1631 Y a_5765_5409# 0
C1632 a_7669_14003# a_7113_13395# 0.28206f
C1633 a_5606_1757# a_5735_1783# 0.00758f
C1634 a_23731_14309# VPWR 0.15203f
C1635 a_15113_5825# a_15227_5715# 0
C1636 a_11243_11891# a_12809_13987# 0.00264f
C1637 a_23731_14309# sky130_fd_sc_hd__mux4_1_0.VPB 0.22258f
C1638 a_11202_5441# a_11541_5723# 0.04737f
C1639 a_10857_14747# a_12135_15219# 0
C1640 a_9725_14509# VPWR 0.00474f
C1641 a_4546_2153# VGND 0.18648f
C1642 a_10088_5837# a_9725_5837# 0.00847f
C1643 a_3738_1787# sky130_fd_sc_hd__inv_1_0.Y 0.00167f
C1644 a_13774_5829# VGND 0.1873f
C1645 a_13147_5829# VPWR 0
C1646 a_4880_2153# VGND 0.00245f
C1647 a_4837_16089# a_4753_16089# 0.00234f
C1648 a_9865_15329# w_10872_13125# 0.00114f
C1649 w_9394_13055# a_9475_14759# 0
C1650 a_14066_1769# a_13315_2025# 0.00682f
C1651 a_6087_14735# a_5895_14763# 0
C1652 a_11049_14719# a_11679_15219# 0.00232f
C1653 a_11160_1747# sky130_fd_sc_hd__inv_1_0.A 0.00203f
C1654 w_11050_5382# A 0.00615f
C1655 w_9490_15543# a_9587_15357# 0.05631f
C1656 a_10611_5471# sky130_fd_sc_hd__mux2_1_0.S 0.04731f
C1657 a_6696_2149# sky130_fd_sc_hd__inv_1_0.A 0
C1658 a_3199_1791# a_3738_1787# 0.0725f
C1659 a_23511_14701# VPWR 0.07721f
C1660 a_16871_4938# sky130_fd_sc_hd__mux2_1_0.VPB 0.07806f
C1661 a_23511_14701# sky130_fd_sc_hd__mux4_1_0.VPB 0.02285f
C1662 a_4763_14775# VGND 0.02642f
C1663 a_24152_14385# a_24318_14385# 0.05583f
C1664 Y VGND 1.11075f
C1665 a_5606_1757# a_5069_1787# 0
C1666 a_8262_5405# VGND 0.18713f
C1667 a_15602_2131# VPWR 0.01894f
C1668 a_14864_4585# w_12894_4504# 0.00188f
C1669 VGND a_1950_5025# 0.40871f
C1670 a_11569_4849# w_12894_4504# 0
C1671 a_12320_4593# VPWR 0
C1672 a_17125_4938# sky130_fd_sc_hd__mux2_1_0.A1 0.19521f
C1673 a_4849_11293# a_4913_13781# 0.26616f
C1674 w_9402_14723# a_9587_15357# 0.00155f
C1675 a_9360_4571# VGND 0.41248f
C1676 a_9725_5471# w_9180_5386# 0.01092f
C1677 a_11986_4959# a_11569_4849# 0.06611f
C1678 a_13046_4563# a_13385_4845# 0.04737f
C1679 a_9589_12125# a_9467_13091# 0.00144f
C1680 a_9875_13765# a_9867_12097# 0.00627f
C1681 a_4837_16089# a_5975_12927# 0
C1682 w_5786_13983# a_4913_13781# 0.00175f
C1683 sky130_fd_sc_hd__inv_1_2.A a_23511_14701# 0.04613f
C1684 a_8566_2145# VPWR 0
C1685 VPWR A 0.3547f
C1686 a_11595_5467# a_11541_5723# 0.00386f
C1687 a_23731_14309# ui_in[1] 0.48785f
C1688 a_13175_4589# VGND 0
C1689 A sky130_fd_sc_hd__mux4_1_0.VPB 0.08221f
C1690 a_13018_5437# a_13411_5829# 0.02301f
C1691 a_5861_5409# a_5636_5017# 0.00559f
C1692 a_15936_2131# VGND 0.00236f
C1693 a_6087_14735# VPWR 0.36336f
C1694 w_6756_13609# a_4837_16089# 0
C1695 a_9811_11277# VPWR 0.42529f
C1696 a_9465_16323# a_9865_15329# 0
C1697 a_9477_11527# a_9467_13091# 0.00102f
C1698 VGND w_9180_5386# 0.56712f
C1699 a_3949_5413# a_3820_5021# 0.00792f
C1700 VGND a_15602_1765# 0.01439f
C1701 a_14946_4905# a_15227_5715# 0.04605f
C1702 a_13315_2025# VPWR 0.34548f
C1703 sky130_fd_sc_hd__inv_1_2.A A 0.00503f
C1704 a_9597_13793# a_9587_15357# 0
C1705 a_15644_5825# A 0.00186f
C1706 a_13357_5719# VPWR 0.35551f
C1707 a_10046_1777# a_9683_1777# 0.00985f
C1708 a_5903_5017# a_5975_5299# 0.21146f
C1709 a_9867_12097# w_9404_11491# 0.00119f
C1710 a_8755_1779# VGND 0.67634f
C1711 VGND a_4505_13107# 0.29689f
C1712 sky130_fd_sc_hd__inv_1_2.Y VGND 0.40404f
C1713 a_23511_14701# ui_in[1] 0.00322f
C1714 sky130_fd_sc_hd__mux2_1_0.A0 VPWR 0.13683f
C1715 a_12250_1773# VGND 0
C1716 w_4432_13071# a_4515_11543# 0
C1717 w_9208_4512# sky130_fd_sc_hd__inv_1_0.A 0.00107f
C1718 a_6717_15235# a_7173_15235# 0
C1719 a_7113_13395# VPWR 0.24839f
C1720 ua[6] VPWR 0
C1721 a_14888_5433# a_15227_5715# 0.04737f
C1722 w_11050_5382# a_9671_5727# 0
C1723 a_13046_4563# a_13285_5437# 0
C1724 a_4587_13107# VPWR 0.02512f
C1725 a_23677_14335# A 0
C1726 a_6944_13645# a_7113_13395# 0
C1727 sky130_fd_sc_hd__inv_1_0.Y w_5454_1698# 0.00152f
C1728 a_13271_4589# sky130_fd_sc_hd__inv_1_0.A 0
C1729 w_11078_4508# a_11202_5441# 0
C1730 a_6635_15235# sky130_fd_sc_hd__inv_1_2.Y 0.1684f
C1731 a_15239_1765# a_15602_1765# 0.00985f
C1732 a_4635_13809# a_4625_15373# 0
C1733 a_11499_2029# a_12924_1769# 0
C1734 a_6281_11907# a_7113_13395# 0.19825f
C1735 a_14946_4905# a_13802_4589# 0
C1736 a_9865_15329# a_10937_12911# 0
C1737 a_13313_4563# sky130_fd_sc_hd__inv_1_0.A 0
C1738 a_14255_1769# a_15602_1765# 0.08907f
C1739 a_11178_4593# a_11359_4959# 0
C1740 ui_in[1] A 0.08699f
C1741 a_10046_1777# a_10569_1777# 0
C1742 VGND a_9419_1777# 0
C1743 a_9238_1777# a_7815_2035# 0
C1744 a_24318_14385# VPWR 0
C1745 a_9671_5727# VPWR 0.35696f
C1746 a_9867_12097# a_4915_10549# 0.00417f
C1747 a_24318_14385# sky130_fd_sc_hd__mux4_1_0.VPB 0.00426f
C1748 VGND w_5906_12121# 0.02048f
C1749 a_9673_15357# VGND 0.00661f
C1750 a_5851_13769# a_5975_12927# 0
C1751 a_11331_5833# a_11150_5467# 0
C1752 Y a_3820_5021# 0.00242f
C1753 a_1898_5051# VGND 0.09486f
C1754 w_10748_13967# VPWR 0.0898f
C1755 a_4546_2153# w_3638_1702# 0.00139f
C1756 w_12866_5378# a_13385_4845# 0.00166f
C1757 a_9589_12125# VPWR 0.38028f
C1758 a_16006_4951# a_15255_4841# 0.00696f
C1759 a_7869_2145# VGND 0.20146f
C1760 a_7845_5295# A 0.00297f
C1761 a_11351_13753# a_11824_13629# 0.24537f
C1762 a_5765_5043# VPWR 0.00115f
C1763 uo_out[0] uo_out[1] 0.03102f
C1764 w_6756_13609# a_5851_13769# 0.00132f
C1765 a_15281_5459# a_15227_5715# 0.00386f
C1766 a_2145_2157# a_2259_2047# 0
C1767 a_11916_1773# a_11553_1773# 0.00985f
C1768 a_17339_4938# A 0.0023f
C1769 a_7454_5039# VPWR 0.07407f
C1770 a_4913_13781# w_4440_14739# 0
C1771 a_5606_1757# a_5873_1757# 0.11512f
C1772 a_11019_12911# a_9811_11277# 0.00146f
C1773 a_4847_14525# a_7173_15235# 0
C1774 a_15227_5715# sky130_fd_sc_hd__mux2_1_0.S 0
C1775 a_12135_15219# VGND 0.32171f
C1776 a_9477_11527# VPWR 0.3853f
C1777 a_10046_2143# VGND 0.1864f
C1778 a_12135_15219# a_9799_16073# 0.04819f
C1779 a_7635_5405# a_7899_5405# 0
C1780 a_13439_4589# VGND 0.01261f
C1781 a_13411_5829# a_13243_5829# 0
C1782 w_6570_15449# a_4837_16089# 0.09702f
C1783 w_9500_13979# a_9811_11277# 0.00123f
C1784 a_15045_4585# a_14325_4589# 0
C1785 a_16006_4951# VGND 0
C1786 VPWR a_14836_5459# 0.07614f
C1787 a_4513_14775# w_4432_13071# 0
C1788 a_4635_13809# w_4538_13995# 0.05631f
C1789 w_11050_5382# a_11569_4849# 0.00166f
C1790 a_9559_11527# a_9811_11277# 0
C1791 w_11532_15433# a_11049_14719# 0.06196f
C1792 a_2079_5417# VPWR 0
C1793 a_5554_1783# a_5069_1787# 0.02709f
C1794 VGND a_4159_5303# 1.20044f
C1795 a_10450_4597# VGND 0
C1796 a_11767_15219# VGND 0.00334f
C1797 a_13243_5463# VPWR 0
C1798 a_24318_14385# ui_in[1] 0.00255f
C1799 a_13439_4955# a_13313_4563# 0.04534f
C1800 a_11767_15219# a_9799_16073# 0
C1801 w_4440_14739# a_4503_16339# 0
C1802 w_12866_5378# a_13285_5437# 0.24672f
C1803 a_4183_1787# a_4015_1787# 0
C1804 a_9332_5445# sky130_fd_sc_hd__mux2_1_0.S 0
C1805 a_9811_11277# a_9549_13091# 0
C1806 a_9699_4853# a_10116_4963# 0.06611f
C1807 a_11178_4593# w_9208_4512# 0.00188f
C1808 a_6003_11935# a_4837_16089# 0
C1809 a_12509_4593# w_11078_4508# 0.01094f
C1810 w_11050_5382# a_11595_5833# 0
C1811 a_7113_13395# w_9500_13979# 0
C1812 a_2313_2157# a_2259_2047# 0.03622f
C1813 a_13774_5463# VPWR 0.20622f
C1814 a_6392_5409# VGND 0.18646f
C1815 a_11569_4849# VPWR 0.35469f
C1816 a_14864_4585# VPWR 0.09402f
C1817 a_5999_2149# w_5454_1698# 0
C1818 a_9809_14509# VGND 0.43095f
C1819 a_7919_14003# a_7173_15235# 0
C1820 a_4849_11293# a_4847_14525# 0.00506f
C1821 a_9683_13793# VPWR 0.003f
C1822 a_9809_14509# a_9799_16073# 0.46421f
C1823 sky130_fd_sc_hd__inv_1_0.Y a_4546_2153# 0
C1824 a_7845_5295# a_9671_5727# 0
C1825 sky130_fd_sc_hd__inv_1_0.Y a_4880_2153# 0
C1826 a_11051_11919# a_9877_10533# 0
C1827 a_11595_5833# VPWR 0.00668f
C1828 VPWR a_9725_14759# 0.32009f
C1829 a_7731_5039# VGND 0
C1830 a_13046_4563# sky130_fd_sc_hd__inv_1_0.A 0
C1831 a_13313_4563# a_13802_4955# 0.03325f
C1832 a_15978_5825# A 0
C1833 a_24241_14651# ui_in[0] 0.00168f
C1834 a_9675_12125# VPWR 0.00297f
C1835 a_5903_5017# a_5636_5017# 0.11512f
C1836 a_6805_15235# VPWR 0.00151f
C1837 a_11230_4567# a_11455_4959# 0.00559f
C1838 uio_in[3] uio_in[4] 0.03102f
C1839 VGND VPB 0.0297f
C1840 a_3199_1791# a_4546_2153# 0.03325f
C1841 a_4015_2153# a_4129_2043# 0
C1842 a_14946_4905# a_13385_4845# 0.00318f
C1843 a_3919_2153# a_4183_2153# 0
C1844 a_9811_11277# a_10895_13753# 0
C1845 a_13774_5829# a_13411_5829# 0.00847f
C1846 a_9465_16323# a_9547_16323# 0.00641f
C1847 a_4903_15345# a_6021_13769# 0.00818f
C1848 Y a_5861_5409# 0
C1849 a_7669_14003# a_7847_14003# 0.00412f
C1850 a_9589_12125# w_9500_13979# 0
C1851 w_4432_13071# a_4839_12857# 0.02723f
C1852 a_9811_11277# a_11243_11891# 0.00683f
C1853 a_14846_1739# a_14975_2131# 0.00792f
C1854 a_11359_4593# a_10639_4597# 0
C1855 a_9809_14509# w_9394_13055# 0
C1856 a_10937_12911# a_12075_13379# 0
C1857 a_9875_13765# VGND 0.70497f
C1858 a_9801_12841# a_9877_10533# 0.00243f
C1859 VGND sky130_fd_sc_hd__inv_1_3.VPB 0.01283f
C1860 a_9875_13765# a_9799_16073# 0.01745f
C1861 a_2259_2047# w_1768_1706# 0.10454f
C1862 w_12824_1684# VPWR 0.51515f
C1863 a_11427_5467# a_10611_5471# 0
C1864 VGND a_9725_5837# 0.25449f
C1865 a_11623_4959# a_10611_5471# 0
C1866 a_2343_5051# w_1798_4966# 0.01092f
C1867 w_10674_14933# a_9811_11277# 0.08584f
C1868 a_23731_14309# a_23511_14701# 0.00549f
C1869 a_4635_13809# VPWR 0.37531f
C1870 a_11597_15219# a_11824_13629# 0
C1871 a_6862_13645# a_5975_12927# 0
C1872 Y a_2706_5417# 0.0357f
C1873 w_14764_4500# VPWR 0.52659f
C1874 a_15672_4951# a_15255_4841# 0.06611f
C1875 a_11089_13753# a_11351_13753# 0
C1876 a_15978_5825# sky130_fd_sc_hd__mux2_1_0.A0 0
C1877 a_9811_11277# a_10983_13753# 0
C1878 a_9477_11527# a_9559_11527# 0.00641f
C1879 a_8262_5039# sky130_fd_sc_hd__mux2_1_0.S 0
C1880 a_10965_11919# VPWR 0.1599f
C1881 a_15141_4585# VPWR 0
C1882 a_6862_13645# w_6756_13609# 0.06114f
C1883 a_15255_4841# sky130_fd_sc_hd__mux2_1_0.A1 0.14436f
C1884 a_3820_5021# a_4159_5303# 0.04737f
C1885 a_9801_12841# w_10868_12105# 0.00131f
C1886 a_4849_11293# a_5933_13769# 0
C1887 VGND w_9404_11491# 0.07411f
C1888 a_23731_14309# A 0.1036f
C1889 a_7899_5039# a_8262_5039# 0.00985f
C1890 a_9717_12841# a_9811_11277# 0
C1891 a_10611_5471# a_10088_5471# 0
C1892 w_9394_13055# a_9875_13765# 0.00226f
C1893 a_9801_12841# a_9475_14759# 0.00442f
C1894 a_11160_1747# w_11008_1688# 0.05213f
C1895 ui_in[7] ui_in[6] 0.03102f
C1896 a_15672_4951# VGND 0
C1897 a_13147_5829# A 0
C1898 a_9465_16323# a_9587_15357# 0.00144f
C1899 a_6885_1783# a_6696_2149# 0
C1900 a_9461_5837# a_9280_5471# 0
C1901 a_9753_4963# a_10116_4963# 0.00847f
C1902 a_5554_1783# a_5873_1757# 0.04799f
C1903 VGND w_5910_13141# 0.02002f
C1904 a_13439_4955# a_13046_4563# 0.02301f
C1905 a_10569_1777# a_11499_2029# 0.21188f
C1906 a_9238_1777# VGND 0.08667f
C1907 a_7635_5039# VGND 0
C1908 sky130_fd_sc_hd__mux2_1_0.A1 VGND 0.08121f
C1909 a_4045_5047# VPWR 0
C1910 a_4183_1787# a_4546_1787# 0.00985f
C1911 w_10748_13967# a_11243_11891# 0
C1912 a_23511_14701# A 0.00138f
C1913 a_9589_12125# a_11243_11891# 0
C1914 a_13147_5463# a_13018_5437# 0.00758f
C1915 a_9597_13793# a_9717_13091# 0
C1916 w_4440_14739# a_4847_14525# 0.02435f
C1917 a_11160_1747# a_11108_1773# 0.1439f
C1918 a_4763_14775# a_4903_15345# 0.00327f
C1919 a_14325_4589# a_13313_4563# 0
C1920 a_15227_5715# a_14297_5463# 0.21188f
C1921 a_4515_11543# VGND 0.29765f
C1922 VGND w_4442_11507# 0.07411f
C1923 a_9585_4597# a_9753_4597# 0
C1924 a_13385_4845# sky130_fd_sc_hd__mux2_1_0.S 0
C1925 a_4915_10549# VGND 1.01177f
C1926 a_9557_14759# a_9475_14759# 0.00641f
C1927 a_4913_13781# a_6129_12927# 0
C1928 a_4847_14525# a_4711_15373# 0
C1929 sky130_fd_sc_hd__inv_1_5.Y VGND 0.39119f
C1930 a_13201_2135# VPWR 0
C1931 a_12481_5467# VGND 0.08017f
C1932 a_4849_11293# a_6329_12927# 0.00976f
C1933 a_9727_11277# VPWR 0.00377f
C1934 VGND w_5712_14949# 0.0161f
C1935 a_15255_4841# a_14916_4559# 0.04737f
C1936 a_7847_14003# VPWR 0
C1937 w_4530_12327# VGND 0.11704f
C1938 a_13313_4563# a_12994_4589# 0.04799f
C1939 a_6089_11935# VPWR 0
C1940 a_4837_16089# a_4905_12113# 0
C1941 a_5903_5017# a_6915_5043# 0
C1942 a_24318_14385# a_23731_14309# 0.02707f
C1943 a_6635_15235# w_5712_14949# 0
C1944 a_11230_4567# a_11359_4959# 0.00792f
C1945 VGND a_12881_13987# 0
C1946 a_4015_2153# a_3790_1761# 0.00559f
C1947 a_7847_14003# a_6281_11907# 0.00264f
C1948 a_13369_1769# VPWR 0.17557f
C1949 a_16006_4585# a_15255_4841# 0.00682f
C1950 a_6281_11907# a_6089_11935# 0
C1951 a_5809_14763# a_5895_14763# 0.00658f
C1952 a_13357_5719# A 0.00759f
C1953 w_9394_13055# a_4915_10549# 0.00179f
C1954 a_10046_1777# VGND 0.01329f
C1955 sky130_fd_sc_hd__mux2_1_0.A1 a_17125_5265# 0.00499f
C1956 a_11351_13753# VPWR 0.38708f
C1957 a_14916_4559# VGND 0
C1958 a_10813_13753# w_12566_13951# 0
C1959 a_7669_14003# a_7751_14003# 0.00695f
C1960 a_4903_15345# sky130_fd_sc_hd__inv_1_2.Y 0
C1961 a_10380_1777# VPWR 0
C1962 sky130_fd_sc_hd__mux2_1_0.S a_13285_5437# 0.04118f
C1963 a_6862_13645# w_6570_15449# 0
C1964 sky130_fd_sc_hd__mux2_1_0.A0 A 0.00975f
C1965 a_24241_14651# sky130_fd_sc_hd__inv_1_0.A 0.03575f
C1966 Y w_1798_4966# 0.25023f
C1967 a_10611_5471# a_11202_5441# 0.11887f
C1968 a_15978_5459# VGND 0
C1969 a_1950_5025# w_1798_4966# 0.05213f
C1970 uio_oe[7] uio_oe[6] 0.03102f
C1971 a_16006_4585# VGND 0
C1972 a_4753_16339# a_4625_15373# 0
C1973 a_11291_12911# a_11824_13629# 0.10646f
C1974 VPWR a_14108_5829# 0
C1975 a_2079_5417# a_2343_5417# 0
C1976 a_6389_13769# VGND 0.25955f
C1977 a_8113_13753# VGND 0.15767f
C1978 VGND a_14975_2131# 0.00305f
C1979 w_9502_10747# VGND 0.12086f
C1980 a_8113_13753# a_9799_16073# 0.36356f
C1981 Y a_4576_5413# 0
C1982 a_4513_14775# VGND 0.29736f
C1983 a_5809_14763# VPWR 0.1486f
C1984 a_24318_14385# A 0.04268f
C1985 a_9671_5727# A 0.00739f
C1986 a_9290_1751# VPWR 0.29556f
C1987 Y a_5903_5017# 0.0011f
C1988 a_11243_11891# a_12713_13987# 0.00373f
C1989 a_11160_1747# a_11289_1773# 0.00758f
C1990 a_14946_4905# sky130_fd_sc_hd__inv_1_0.A 0
C1991 a_9865_15329# a_9475_14759# 0.00566f
C1992 a_14846_1739# a_14975_1765# 0.00758f
C1993 a_4505_13107# a_4755_13107# 0.02504f
C1994 a_14846_1739# a_15071_2131# 0.00559f
C1995 a_4597_11543# VGND 0.00172f
C1996 a_11230_4567# w_9208_4512# 0
C1997 a_6127_13769# VPWR 0.0014f
C1998 a_4015_2153# VPWR 0
C1999 a_9811_11277# w_10748_13967# 0.10705f
C2000 VPWR sky130_fd_sc_hd__inv_1_0.VPB 0.06793f
C2001 a_11595_5467# a_10611_5471# 0.08312f
C2002 w_11718_13593# a_11824_13629# 0.06114f
C2003 a_4837_16089# a_7173_15235# 0.04819f
C2004 a_9589_12125# a_9811_11277# 0.0022f
C2005 a_9332_5445# a_7899_5405# 0
C2006 a_7454_5039# A 0.00118f
C2007 a_4753_16339# w_4430_16303# 0.01327f
C2008 a_12924_1769# VGND 0.08648f
C2009 a_4503_16339# a_4625_15373# 0.00144f
C2010 a_9585_4597# VPWR 0.00132f
C2011 a_10965_11919# a_11243_11891# 0.11706f
C2012 a_11455_4959# VPWR 0
C2013 a_14836_5459# A 0.003f
C2014 a_9477_11527# a_9811_11277# 0.16782f
C2015 a_13046_4563# a_12994_4589# 0.1439f
C2016 a_1920_1765# a_2259_2047# 0.04737f
C2017 a_6362_2149# VPWR 0.01976f
C2018 a_15255_4841# w_14736_5374# 0.00166f
C2019 w_11050_5382# a_11958_5833# 0.00139f
C2020 a_5861_5043# VGND 0
C2021 a_13243_5463# A 0
C2022 a_7751_14003# VPWR 0
C2023 VGND a_4839_12857# 1.32139f
C2024 a_5099_5047# VGND 0.06389f
C2025 a_9801_12841# a_12135_15219# 0.00685f
C2026 a_1898_5051# w_1798_4966# 0.01793f
C2027 a_12320_4593# a_11569_4849# 0.00682f
C2028 a_11597_15219# VPWR 0.3359f
C2029 a_15672_4585# a_15255_4841# 0.03016f
C2030 VGND a_24234_14385# 0.05676f
C2031 a_13357_5719# a_14836_5459# 0
C2032 a_15239_2131# a_14975_2131# 0
C2033 a_4546_1787# a_5873_1757# 0
C2034 a_6281_11907# a_7751_14003# 0.00373f
C2035 a_12320_4959# VPWR 0
C2036 a_4913_13781# w_4538_13995# 0.01958f
C2037 a_12481_5467# a_11541_5723# 0.12975f
C2038 a_13385_4845# a_14297_5463# 0
C2039 a_4849_11293# a_4837_16089# 0.03118f
C2040 a_13439_4955# a_14946_4905# 0
C2041 a_11569_4849# A 0
C2042 VGND w_14736_5374# 0.29321f
C2043 a_13774_5463# A 0
C2044 a_14864_4585# A 0
C2045 sky130_fd_sc_hd__inv_1_5.Y sky130_fd_sc_hd__inv_1_4.VPB 0.00994f
C2046 a_9360_4571# a_9489_4597# 0.00758f
C2047 a_11958_5833# VPWR 0.01821f
C2048 a_13243_5463# a_13357_5719# 0
C2049 a_4837_16089# w_5786_13983# 0.06973f
C2050 a_12481_5467# a_12966_5463# 0.02709f
C2051 a_10639_4597# VGND 0.65621f
C2052 a_15309_4585# sky130_fd_sc_hd__inv_1_0.A 0
C2053 w_4430_16303# a_4503_16339# 0.06993f
C2054 sky130_fd_sc_hd__inv_1_2.A a_11597_15219# 0
C2055 a_9360_4571# a_9699_4853# 0.04737f
C2056 a_13313_4563# w_12894_4504# 0.24672f
C2057 VGND a_4723_10577# 0.00697f
C2058 a_15672_4585# VGND 0
C2059 a_10771_14747# VPWR 0.1486f
C2060 a_2175_5417# Y 0
C2061 a_11595_5833# A 0.00169f
C2062 a_11916_1773# sky130_fd_sc_hd__inv_1_0.A 0
C2063 a_2175_5417# a_1950_5025# 0.00559f
C2064 a_13357_5719# a_13774_5463# 0.03016f
C2065 a_9877_10533# a_12075_13379# 0.16207f
C2066 a_15045_4585# VPWR 0.00135f
C2067 a_6726_5409# VPWR 0
C2068 a_11291_12911# a_9467_13091# 0
C2069 a_9801_12841# a_9809_14509# 0.20053f
C2070 a_5851_13769# a_7173_15235# 0
C2071 a_15017_5825# a_15281_5825# 0
C2072 a_11331_5467# a_10611_5471# 0
C2073 a_9753_4597# w_9208_4512# 0.01092f
C2074 a_7605_2145# VGND 0.00305f
C2075 a_9811_11277# a_9725_14759# 0
C2076 a_6087_14735# a_6805_15235# 0.00366f
C2077 a_9699_4853# w_9180_5386# 0.00166f
C2078 w_14694_1680# a_14846_1739# 0.05213f
C2079 a_9675_12125# a_9811_11277# 0
C2080 a_9589_12125# a_9477_11527# 0
C2081 a_7506_5013# w_7354_4954# 0.05213f
C2082 a_14946_4905# a_13802_4955# 0
C2083 a_14297_5463# a_13285_5437# 0
C2084 a_10895_13753# a_11351_13753# 0
C2085 VGND a_3229_5051# 0.67714f
C2086 a_12292_5467# VGND 0
C2087 a_4129_2043# a_5606_1757# 0.00492f
C2088 a_4753_16339# VPWR 0.32314f
C2089 a_11597_15219# a_11873_15219# 0.00119f
C2090 a_12631_13987# a_9877_10533# 0.0762f
C2091 a_11351_13753# a_11243_11891# 0.00255f
C2092 a_4576_5413# a_4159_5303# 0.06611f
C2093 a_11499_2029# VGND 1.19976f
C2094 a_9238_1777# a_9419_2143# 0
C2095 w_14764_4500# A 0
C2096 a_13315_2025# w_12824_1684# 0.10454f
C2097 a_9557_14759# a_9809_14509# 0
C2098 a_2289_5307# a_2706_5051# 0.03016f
C2099 a_4159_5303# a_5903_5017# 0.00412f
C2100 a_9308_4597# a_9489_4963# 0
C2101 a_11160_1747# ua[5] 0
C2102 a_9801_12841# a_9875_13765# 0.44871f
C2103 a_3949_5047# a_4213_5047# 0
C2104 a_11351_13753# a_10983_13753# 0
C2105 a_4913_13781# VPWR 0.60287f
C2106 a_15309_4951# a_14325_4589# 0.04534f
C2107 a_15113_5825# a_15281_5825# 0
C2108 a_9865_15329# a_9673_15357# 0.00101f
C2109 a_11359_4959# VPWR 0
C2110 a_10965_11919# a_9811_11277# 0.10332f
C2111 a_4849_11293# a_5851_13769# 0.17627f
C2112 a_11160_1747# VPWR 0.29475f
C2113 w_5786_13983# a_5851_13769# 0.08205f
C2114 a_6392_5409# a_5903_5017# 0.03325f
C2115 a_14975_1765# VGND 0
C2116 a_15071_2131# VGND 0.00231f
C2117 a_4847_14525# a_4625_15373# 0.00215f
C2118 a_10813_13753# VGND 0.15513f
C2119 a_6696_2149# VPWR 0
C2120 a_4903_15345# w_5910_13141# 0.00114f
C2121 a_10813_13753# a_9799_16073# 0.08387f
C2122 a_10937_12911# a_11091_12911# 0.00401f
C2123 a_7506_5013# w_5484_4958# 0
C2124 a_15255_4841# a_17125_4938# 0
C2125 a_9801_12841# w_9404_11491# 0
C2126 a_4627_12141# w_4540_10763# 0
C2127 a_9290_1751# a_9515_1777# 0.00487f
C2128 a_4503_16339# VPWR 0.39579f
C2129 a_9683_1777# VGND 0.01556f
C2130 a_9280_5471# sky130_fd_sc_hd__mux2_1_0.S 0
C2131 a_13732_1769# sky130_fd_sc_hd__inv_1_0.A 0
C2132 uo_out[7] uio_out[0] 0.03102f
C2133 a_4837_16089# w_4440_14739# 0
C2134 a_10611_5471# w_9180_5386# 0.02026f
C2135 a_11499_2029# a_11385_1773# 0
C2136 a_9589_12125# a_9675_12125# 0.00658f
C2137 a_9865_15329# a_12135_15219# 0
C2138 a_4915_10549# w_9492_12311# 0.00193f
C2139 a_3790_1761# a_2259_2047# 0.00446f
C2140 a_11291_12911# VPWR 0.23898f
C2141 a_5903_5017# VPB 0
C2142 a_11049_14719# a_11824_13629# 0
C2143 a_9360_4571# a_9753_4963# 0.02301f
C2144 a_14975_1765# a_15239_1765# 0
C2145 sky130_fd_sc_hd__inv_1_5.Y a_23677_14701# 0.01449f
C2146 a_13046_4563# w_12894_4504# 0.05213f
C2147 a_17125_4938# VGND 0.16937f
C2148 a_15644_5459# a_15227_5715# 0.03016f
C2149 a_14255_1769# a_14975_1765# 0
C2150 a_4903_15345# w_5712_14949# 0.00546f
C2151 a_1868_1791# a_2049_2157# 0
C2152 a_3790_1761# a_3919_1787# 0.00758f
C2153 a_14325_4589# a_14946_4905# 0.58451f
C2154 w_4430_16303# a_4847_14525# 0
C2155 a_10088_5837# VGND 0.22304f
C2156 a_3919_2153# a_3738_1787# 0
C2157 a_13046_4563# a_13271_4955# 0.00559f
C2158 a_10569_1777# VGND 0.6772f
C2159 a_13411_5463# VPWR 0.16932f
C2160 a_3820_5021# a_3229_5051# 0.11887f
C2161 a_9290_1751# a_9683_2143# 0.02301f
C2162 a_9727_11277# a_9811_11277# 0.00206f
C2163 a_13201_2135# a_13315_2025# 0
C2164 a_9801_12841# a_4915_10549# 0
C2165 a_4765_11543# a_4505_13107# 0
C2166 a_10450_4597# a_9699_4853# 0.00682f
C2167 a_6911_15235# VGND 0.00384f
C2168 a_9589_12125# a_10965_11919# 0
C2169 a_14946_4905# a_15281_5825# 0.00186f
C2170 a_3949_5413# a_4213_5413# 0
C2171 a_10639_4597# a_11541_5723# 0
C2172 a_9475_14759# a_9587_15357# 0
C2173 w_9208_4512# VPWR 0.78497f
C2174 a_17053_4938# VPWR 0
C2175 a_9809_14509# a_9865_15329# 0.15229f
C2176 a_14325_4589# a_14888_5433# 0
C2177 a_13271_4589# VPWR 0
C2178 w_4432_13071# VGND 0.07276f
C2179 a_13243_1743# sky130_fd_sc_hd__inv_1_0.A 0.00204f
C2180 a_13732_2135# a_13243_1743# 0.03325f
C2181 w_11718_13593# VPWR 0.08767f
C2182 VGND a_15936_1765# 0
C2183 a_6911_15235# a_6635_15235# 0.00119f
C2184 a_11569_4849# a_11595_5833# 0
C2185 a_4503_16339# a_4585_16339# 0.00641f
C2186 a_13369_1769# a_13315_2025# 0.00386f
C2187 a_11427_5833# VGND 0.00241f
C2188 a_15239_2131# a_15071_2131# 0
C2189 a_9811_11277# a_11351_13753# 0.00488f
C2190 a_13313_4563# VPWR 0.97733f
C2191 w_10674_14933# a_11597_15219# 0
C2192 w_12566_13951# VGND 0.00711f
C2193 a_7847_14003# a_7113_13395# 0.00121f
C2194 a_6717_15235# VPWR 0
C2195 w_12566_13951# a_9799_16073# 0
C2196 a_15281_5825# a_14888_5433# 0.02301f
C2197 sky130_fd_sc_hd__mux2_1_0.A1 sky130_fd_sc_hd__mux2_1_0.VPB 0.09504f
C2198 a_14108_5829# A 0
C2199 a_7669_14003# a_7919_14003# 0.00876f
C2200 a_4129_2043# a_5554_1783# 0
C2201 a_4903_15345# a_6389_13769# 0
C2202 a_6057_12927# a_4839_12857# 0.00149f
C2203 a_2259_2047# VPWR 0.3445f
C2204 a_9867_12097# VGND 0.43935f
C2205 a_9867_12097# a_9799_16073# 0
C2206 ua[7] w_1768_1706# 0
C2207 w_14694_1680# VGND 0.29099f
C2208 a_4513_14775# a_4903_15345# 0.00566f
C2209 a_12292_5467# a_11541_5723# 0.00682f
C2210 a_5975_12927# a_4505_13107# 0
C2211 a_17125_4938# a_17346_5265# 0.00783f
C2212 a_10569_1777# a_11385_1773# 0
C2213 a_9875_13765# a_9865_15329# 0.1161f
C2214 w_10674_14933# a_10771_14747# 0.05631f
C2215 a_7815_2035# VGND 1.2f
C2216 a_6087_14735# a_5809_14763# 0.1109f
C2217 a_9308_4597# VGND 0.08793f
C2218 a_9599_10561# a_9877_10533# 0.1296f
C2219 a_6862_13645# a_4849_11293# 0
C2220 sky130_fd_sc_hd__inv_1_4.A sky130_fd_sc_hd__inv_1_5.VPB 0
C2221 a_14864_4585# w_14764_4500# 0.01793f
C2222 a_13357_5719# a_14108_5829# 0.00696f
C2223 a_3919_1787# VPWR 0.00117f
C2224 a_15309_4585# a_14325_4589# 0.08312f
C2225 a_14325_4589# a_15281_5459# 0
C2226 a_13018_5437# a_13285_5437# 0.11512f
C2227 Y a_4213_5413# 0
C2228 a_24241_14651# a_24774_14701# 0.0098f
C2229 a_9699_4853# a_9725_5837# 0
C2230 VGND a_2079_5051# 0
C2231 a_9801_12841# a_8113_13753# 0.00389f
C2232 a_14325_4589# sky130_fd_sc_hd__mux2_1_0.S 0.03312f
C2233 w_11050_5382# a_11150_5467# 0.01793f
C2234 w_9394_13055# a_9867_12097# 0
C2235 ui_in[0] a_23511_14335# 0.08552f
C2236 a_10857_14747# VGND 0.00618f
C2237 w_14694_1680# a_15239_1765# 0.01092f
C2238 a_10857_14747# a_9799_16073# 0
C2239 w_7604_13967# a_4915_10549# 0.05671f
C2240 a_14846_1739# VGND 0.40101f
C2241 a_5975_12927# w_5906_12121# 0
C2242 a_9477_11527# a_9727_11277# 0.00723f
C2243 w_14694_1680# a_14255_1769# 0.25055f
C2244 a_4847_14525# VPWR 0.36398f
C2245 a_9332_5445# a_8262_5405# 0
C2246 w_10748_13967# a_11351_13753# 0.01492f
C2247 a_5945_2039# VGND 1.20001f
C2248 a_11455_4959# A 0
C2249 a_5606_1757# VPWR 0.29521f
C2250 a_9332_5445# a_9360_4571# 0
C2251 a_9465_16323# w_9392_16287# 0.06993f
C2252 a_12135_15219# a_12075_13379# 0.36868f
C2253 a_9489_4963# VGND 0.00325f
C2254 a_4513_14775# a_4755_13107# 0
C2255 a_4129_2043# a_4015_1787# 0
C2256 a_12976_1743# a_13243_1743# 0.11512f
C2257 VPWR a_11150_5467# 0.07689f
C2258 a_5606_1757# a_5831_1783# 0.00487f
C2259 a_10639_4597# w_11078_4508# 0.25055f
C2260 a_8262_5039# a_6915_5043# 0.08907f
C2261 a_5831_2149# a_5606_1757# 0.00559f
C2262 a_8596_5405# VGND 0.00249f
C2263 a_4903_15345# a_4839_12857# 0.1369f
C2264 a_5069_1787# w_5454_1698# 0.0025f
C2265 a_11289_2139# VGND 0.00305f
C2266 a_9461_5837# VPWR 0
C2267 a_14794_1765# a_14975_2131# 0
C2268 a_9332_5445# w_9180_5386# 0.05213f
C2269 a_14846_1739# a_15239_1765# 0.02283f
C2270 a_10639_4597# a_11455_4593# 0
C2271 a_4637_10577# w_4540_10763# 0.05631f
C2272 a_12135_15219# a_12631_13987# 0.16709f
C2273 a_4129_2043# a_4183_2153# 0.03622f
C2274 w_14694_1680# a_15239_2131# 0
C2275 a_14846_1739# a_14255_1769# 0.11887f
C2276 VGND a_9685_10561# 0.00697f
C2277 a_13105_1769# sky130_fd_sc_hd__inv_1_0.A 0
C2278 a_11958_5833# A 0.00158f
C2279 a_3040_5051# Y 0
C2280 a_11916_1773# w_11008_1688# 0.01154f
C2281 a_7919_14003# VPWR 0
C2282 a_13046_4563# VPWR 0.2975f
C2283 a_7424_1779# w_5454_1698# 0.00188f
C2284 a_11291_12911# a_11243_11891# 0.00298f
C2285 w_7354_4954# sky130_fd_sc_hd__mux2_1_0.S 0.0206f
C2286 a_6281_11907# a_7919_14003# 0
C2287 a_7751_14003# a_7113_13395# 0.00226f
C2288 w_7604_13967# a_6389_13769# 0
C2289 a_9673_15357# a_9587_15357# 0.00658f
C2290 Y a_4045_5413# 0
C2291 a_7899_5039# w_7354_4954# 0.01092f
C2292 a_8113_13753# w_7604_13967# 0.01891f
C2293 a_6726_5409# A 0
C2294 a_11331_5833# a_11202_5441# 0.00792f
C2295 a_5933_13769# VPWR 0
C2296 a_10450_4963# VPWR 0
C2297 a_4905_12113# a_4713_12141# 0
C2298 a_10771_14747# a_9811_11277# 0.10553f
C2299 a_7506_5013# VPWR 0.29452f
C2300 w_6570_15449# sky130_fd_sc_hd__inv_1_2.Y 0.097f
C2301 a_6029_5409# a_5975_5299# 0.03622f
C2302 a_14136_4955# a_13385_4845# 0.00696f
C2303 a_14946_4905# w_12894_4504# 0.00104f
C2304 a_4839_12857# a_4755_13107# 0.08134f
C2305 a_14846_1739# a_15239_2131# 0.02301f
C2306 a_11427_5833# a_11541_5723# 0
C2307 uio_out[3] uio_out[2] 0.03102f
C2308 a_8262_5039# a_9360_4571# 0
C2309 a_2676_2157# VGND 0.18903f
C2310 a_2289_5307# a_3040_5417# 0.00696f
C2311 a_14946_4905# a_13271_4955# 0
C2312 a_11049_14719# VPWR 0.36334f
C2313 a_7731_5405# VGND 0.00235f
C2314 w_11718_13593# a_11243_11891# 0.00315f
C2315 ua[0] a_24234_14385# 0
C2316 a_10116_4597# w_9208_4512# 0.01154f
C2317 sky130_fd_sc_hd__inv_1_2.Y sky130_fd_sc_hd__inv_1_2.VPB 0.02743f
C2318 a_11351_13753# a_12713_13987# 0
C2319 VGND a_5765_5409# 0.00306f
C2320 a_13369_1769# w_12824_1684# 0.01092f
C2321 a_11499_2029# a_11385_2139# 0
C2322 ui_in[2] ui_in[1] 0.03102f
C2323 a_5861_5043# a_5903_5017# 0
C2324 a_8113_13753# a_9865_15329# 0.00176f
C2325 a_11230_4567# sky130_fd_sc_hd__mux2_1_0.S 0
C2326 a_5999_1783# a_5606_1757# 0.02283f
C2327 a_5099_5047# a_5903_5017# 0.02844f
C2328 a_6726_5043# a_5975_5299# 0.00682f
C2329 a_2706_5051# VPWR 0.20629f
C2330 a_15017_5825# VPWR 0
C2331 a_13369_2135# VGND 0.20063f
C2332 a_9727_11527# w_9404_11491# 0.01327f
C2333 a_2049_2157# a_2313_2157# 0
C2334 a_4159_5303# a_4213_5413# 0.03622f
C2335 a_15255_4841# VGND 0.00379f
C2336 a_6029_5043# a_5975_5299# 0.00386f
C2337 VGND a_9725_5471# 0.10237f
C2338 a_4837_16089# a_4625_15373# 0
C2339 a_6329_12927# VPWR 0.23898f
C2340 a_6087_14735# a_4913_13781# 0
C2341 a_9629_2033# a_8755_1779# 0.21161f
C2342 a_4129_2043# a_4546_1787# 0.03016f
C2343 a_13439_4589# a_13802_4589# 0.00985f
C2344 a_3790_1761# a_4015_1787# 0.00487f
C2345 a_13105_1769# a_12976_1743# 0.00758f
C2346 a_7669_14003# a_9597_13793# 0
C2347 a_6003_11935# w_5906_12121# 0.05631f
C2348 w_7604_13967# a_4839_12857# 0
C2349 a_15113_5459# VPWR 0
C2350 w_12866_5378# VPWR 0.51463f
C2351 a_4880_2153# a_5069_1787# 0
C2352 a_4765_11543# a_4515_11543# 0.02504f
C2353 a_6281_11907# a_6329_12927# 0.00298f
C2354 a_10771_14747# w_10748_13967# 0
C2355 a_5873_1757# w_5454_1698# 0.24672f
C2356 a_9809_14509# a_9587_15357# 0.00215f
C2357 a_14325_4589# a_14297_5463# 0.00251f
C2358 a_4765_11543# w_4442_11507# 0.01327f
C2359 a_5554_1783# VPWR 0.07437f
C2360 a_3229_5051# w_1798_4966# 0.02026f
C2361 a_4847_14525# a_4763_14525# 0.00206f
C2362 a_9597_13793# a_9467_13091# 0.00115f
C2363 VGND a_9799_16073# 0.68227f
C2364 a_11455_4959# a_11569_4849# 0
C2365 a_13774_5829# a_13285_5437# 0.03325f
C2366 a_3790_1761# a_4183_2153# 0.02301f
C2367 a_9717_13091# a_9475_14759# 0
C2368 a_8232_2145# sky130_fd_sc_hd__inv_1_0.A 0
C2369 a_11873_15219# a_11049_14719# 0.00651f
C2370 a_9801_12841# a_10813_13753# 0.13074f
C2371 a_15281_5825# a_14297_5463# 0.04534f
C2372 a_9727_11527# a_4915_10549# 0
C2373 a_15113_5825# VPWR 0
C2374 a_6635_15235# VGND 0.13063f
C2375 sky130_fd_sc_hd__mux2_1_0.S w_12894_4504# 0.00112f
C2376 a_7506_5013# a_7845_5295# 0.04737f
C2377 w_5454_1698# sky130_fd_sc_hd__inv_1_0.A 0.00165f
C2378 a_5975_12927# w_5910_13141# 0.04996f
C2379 a_4576_5413# a_3229_5051# 0.03325f
C2380 a_9811_11277# a_11291_12911# 0.00976f
C2381 a_12439_1773# a_12250_2139# 0
C2382 a_6362_1783# w_5454_1698# 0.01154f
C2383 w_4430_16303# a_4837_16089# 0.02445f
C2384 a_5903_5017# a_3229_5051# 0
C2385 a_15309_4951# VPWR 0.00889f
C2386 a_12135_15219# a_11679_15219# 0
C2387 VGND a_15239_1765# 0.01387f
C2388 w_9394_13055# VGND 0.07276f
C2389 a_13411_5463# A 0
C2390 a_11569_4849# a_12320_4959# 0.00696f
C2391 w_9490_15543# VPWR 0.18191f
C2392 a_13243_1743# w_11008_1688# 0.00743f
C2393 a_14255_1769# VGND 0.67529f
C2394 a_3738_1787# w_1768_1706# 0.00188f
C2395 a_24241_14651# VPWR 0.25337f
C2396 w_9208_4512# A 0
C2397 a_17053_4938# A 0
C2398 a_24241_14651# sky130_fd_sc_hd__mux4_1_0.VPB 0.0237f
C2399 a_12881_13987# a_12075_13379# 0.00207f
C2400 a_11385_1773# VGND 0
C2401 VPWR w_9402_14723# 0.16205f
C2402 a_11986_4593# a_10639_4597# 0.08907f
C2403 sky130_fd_sc_hd__inv_1_2.A w_9490_15543# 0
C2404 uio_oe[0] uio_out[7] 0.03102f
C2405 a_4849_11293# a_4713_12141# 0
C2406 a_17125_5265# VGND 0.00352f
C2407 a_9629_2033# a_10046_2143# 0.06611f
C2408 a_13357_5719# a_13411_5463# 0.00386f
C2409 a_4159_5303# a_4045_5413# 0
C2410 a_4015_1787# VPWR 0
C2411 w_6756_13609# a_4915_10549# 0.00404f
C2412 sky130_fd_sc_hd__inv_1_0.Y a_5945_2039# 0
C2413 a_9332_5445# a_9725_5837# 0.02301f
C2414 a_11958_5833# a_11595_5833# 0.00847f
C2415 a_2049_1791# VGND 0
C2416 ui_in[3] ui_in[4] 0.03102f
C2417 a_13313_4563# A 0
C2418 VGND a_17346_5265# 0.00328f
C2419 a_12509_4593# sky130_fd_sc_hd__inv_1_0.A 0
C2420 a_9699_4853# a_10639_4597# 0.13962f
C2421 a_9811_11277# w_11718_13593# 0
C2422 a_14846_1739# a_15071_1765# 0.00487f
C2423 a_11178_4593# a_11202_5441# 0
C2424 a_10422_5471# VPWR 0
C2425 a_6029_5409# a_5636_5017# 0.02301f
C2426 a_6087_14735# a_6717_15235# 0.00232f
C2427 a_14255_1769# a_15239_1765# 0.08312f
C2428 a_12881_13987# a_12631_13987# 0.00876f
C2429 a_9867_12097# w_9492_12311# 0.0247f
C2430 a_4183_2153# VPWR 0.00888f
C2431 a_9809_14509# a_11679_15219# 0.00159f
C2432 uio_oe[2] uio_oe[3] 0.03102f
C2433 a_15239_2131# VGND 0.19769f
C2434 a_9867_12097# a_11051_11919# 0
C2435 a_4837_16089# a_5895_14763# 0
C2436 a_4627_12141# a_4713_12141# 0.00658f
C2437 a_9597_13793# VPWR 0.37502f
C2438 sky130_fd_sc_hd__inv_1_4.A sky130_fd_sc_hd__inv_1_3.VPB 0.02625f
C2439 a_14946_4905# VPWR 1.2932f
C2440 a_13357_5719# a_13313_4563# 0
C2441 a_12439_1773# sky130_fd_sc_hd__inv_1_0.A 0
C2442 a_9801_12841# w_12566_13951# 0
C2443 VGND a_3820_5021# 0.40141f
C2444 a_4905_12113# a_4505_13107# 0
C2445 a_24241_14651# ui_in[1] 0.06316f
C2446 w_4432_13071# a_4755_13107# 0.01327f
C2447 a_13439_4589# a_13385_4845# 0.00386f
C2448 a_17125_4938# sky130_fd_sc_hd__mux2_1_0.VPB 0.04809f
C2449 a_13439_4955# a_13175_4955# 0
C2450 a_4849_11293# a_6021_13769# 0
C2451 a_9801_12841# a_9867_12097# 0.04364f
C2452 a_7669_14003# a_5851_13769# 0
C2453 a_14888_5433# VPWR 0.30504f
C2454 a_15644_5825# a_14946_4905# 0.00336f
C2455 w_7354_4954# a_5975_5299# 0
C2456 a_9671_5727# w_9208_4512# 0
C2457 a_8232_2145# w_7324_1694# 0.00139f
C2458 a_4576_5047# Y 0
C2459 a_15239_2131# a_14255_1769# 0.04534f
C2460 a_4837_16089# VPWR 1.09775f
C2461 a_6029_5043# a_5636_5017# 0.02283f
C2462 a_10937_12911# a_11824_13629# 0
C2463 a_15936_2131# a_15185_2021# 0.00696f
C2464 a_5851_13769# w_4538_13995# 0
C2465 w_6756_13609# a_6389_13769# 0.06723f
C2466 a_10422_5837# VPWR 0
C2467 VGND w_3638_1702# 0.2935f
C2468 w_10674_14933# a_11049_14719# 0.02211f
C2469 a_15185_2021# a_15602_1765# 0.03016f
C2470 a_6087_14735# a_4847_14525# 0.3196f
C2471 a_5636_5017# w_3668_4962# 0
C2472 a_10639_4597# a_10611_5471# 0.00251f
C2473 a_9865_15329# a_10813_13753# 0.16764f
C2474 a_4905_12113# w_5906_12121# 0.08119f
C2475 a_14916_4559# a_15227_5715# 0
C2476 a_2676_2157# sky130_fd_sc_hd__inv_1_0.Y 0.03547f
C2477 a_11150_5467# A 0.00306f
C2478 VGND a_11541_5723# 1.23723f
C2479 w_11050_5382# sky130_fd_sc_hd__mux2_1_0.S 0.00342f
C2480 a_15141_4951# VPWR 0
C2481 a_9801_12841# a_10857_14747# 0
C2482 Y a_4213_5047# 0
C2483 a_11499_2029# a_11916_2139# 0.06611f
C2484 a_7899_5405# w_7354_4954# 0
C2485 VGND a_12966_5463# 0.10729f
C2486 w_10872_13125# a_9467_13091# 0
C2487 VGND sky130_fd_sc_hd__inv_1_4.VPB 0.01319f
C2488 a_5735_2149# VPWR 0
C2489 a_13439_4589# a_13285_5437# 0
C2490 a_15978_5459# a_15227_5715# 0.00682f
C2491 a_6003_11935# w_5910_13141# 0
C2492 a_9599_10561# w_9404_11491# 0
C2493 a_9461_5837# A 0
C2494 w_14694_1680# a_14794_1765# 0.01793f
C2495 a_13243_5463# a_13411_5463# 0
C2496 a_8755_1779# w_9138_1692# 0.24998f
C2497 a_15309_4585# VPWR 0.17334f
C2498 a_15281_5459# VPWR 0.16927f
C2499 sky130_fd_sc_hd__inv_1_5.Y sky130_fd_sc_hd__inv_1_4.A 0.14977f
C2500 a_5999_2149# a_5945_2039# 0.03622f
C2501 a_4595_14775# VPWR 0.02511f
C2502 w_5484_4958# a_5975_5299# 0.10454f
C2503 a_9360_4571# sky130_fd_sc_hd__inv_1_0.A 0
C2504 a_4635_13809# a_4913_13781# 0.1205f
C2505 sky130_fd_sc_hd__mux2_1_0.S VPWR 2.23739f
C2506 a_4546_1787# VPWR 0.20643f
C2507 a_11916_1773# VPWR 0.20655f
C2508 a_13046_4563# A 0
C2509 uo_out[6] uo_out[7] 0.03102f
C2510 a_13175_4589# sky130_fd_sc_hd__inv_1_0.A 0
C2511 a_8113_13753# a_9587_15357# 0.00113f
C2512 a_11623_4959# a_11230_4567# 0.02301f
C2513 a_12439_1773# a_12976_1743# 0
C2514 a_12994_4589# a_13018_5437# 0
C2515 a_7899_5039# VPWR 0.1761f
C2516 a_13774_5463# a_13411_5463# 0.00985f
C2517 a_6003_11935# a_4915_10549# 0
C2518 a_15936_2131# sky130_fd_sc_hd__inv_1_0.A 0
C2519 w_11532_15433# a_12135_15219# 0.01567f
C2520 a_5975_12927# a_4839_12857# 0.30276f
C2521 a_4837_16089# a_4585_16339# 0
C2522 a_9597_13793# w_9500_13979# 0.05631f
C2523 a_7605_1779# VGND 0
C2524 a_4763_14775# a_4849_11293# 0
C2525 sky130_fd_sc_hd__inv_1_2.Y a_7173_15235# 0.002f
C2526 w_4528_15559# a_4625_15373# 0.05631f
C2527 a_11499_2029# a_11553_2139# 0.03622f
C2528 sky130_fd_sc_hd__inv_1_0.A a_15602_1765# 0
C2529 a_5861_5409# VGND 0.00233f
C2530 a_14846_1739# a_14794_1765# 0.1439f
C2531 a_6003_11935# w_4530_12327# 0
C2532 a_4915_10549# a_9599_10561# 0
C2533 a_2145_1791# VGND 0
C2534 w_9392_16287# a_9475_14759# 0
C2535 a_13201_1769# VGND 0
C2536 w_6756_13609# a_4839_12857# 0.00515f
C2537 a_13357_5719# a_13046_4563# 0
C2538 a_7506_5013# A 0.00206f
C2539 VPWR w_4540_10763# 0.166f
C2540 sky130_fd_sc_hd__inv_1_0.Y VGND 1.11393f
C2541 a_6057_12927# VGND 0.00238f
C2542 a_8755_1779# sky130_fd_sc_hd__inv_1_0.A 0.00258f
C2543 uio_in[5] uio_in[4] 0.03102f
C2544 a_5851_13769# VPWR 0.3558f
C2545 a_6392_5043# a_5975_5299# 0.03016f
C2546 a_13313_4563# a_11569_4849# 0.00412f
C2547 a_9671_5727# a_11150_5467# 0
C2548 a_12250_1773# sky130_fd_sc_hd__inv_1_0.A 0
C2549 a_7113_13395# a_7919_14003# 0.00207f
C2550 VGND a_2706_5417# 0.18671f
C2551 uo_out[5] uo_out[4] 0.03102f
C2552 a_5851_13769# a_6281_11907# 0
C2553 a_15071_1765# VGND 0
C2554 a_2049_2157# a_1920_1765# 0.00792f
C2555 VGND a_13411_5829# 0.20231f
C2556 a_11595_5467# a_11958_5467# 0.00985f
C2557 a_3040_5417# VPWR 0
C2558 a_3199_1791# VGND 0.67808f
C2559 ua[7] VPWR 0
C2560 a_9809_14509# w_11532_15433# 0.07233f
C2561 a_6862_13645# a_7669_14003# 0
C2562 a_10569_1777# a_11916_2139# 0.03325f
C2563 a_10046_2143# w_9138_1692# 0.00139f
C2564 a_4849_11293# a_4505_13107# 0.00376f
C2565 a_11623_4959# a_11986_4959# 0.00847f
C2566 sky130_fd_sc_hd__inv_1_0.A a_9419_1777# 0
C2567 a_11049_14719# a_9811_11277# 0.00179f
C2568 a_9419_2143# VGND 0.00305f
C2569 w_10872_13125# VPWR 0.0888f
C2570 w_5786_13983# sky130_fd_sc_hd__inv_1_2.Y 0
C2571 a_15017_5825# A 0
C2572 a_3949_5047# VPWR 0.00114f
C2573 a_15017_5459# VGND 0
C2574 w_11078_4508# VGND 0.28981f
C2575 a_10937_12911# a_9467_13091# 0
C2576 a_6029_5409# Y 0
C2577 a_10046_1777# a_9629_2033# 0.03016f
C2578 a_8113_13753# sky130_fd_sc_hd__inv_1_2.VPB 0.00457f
C2579 a_15071_1765# a_15239_1765# 0
C2580 a_15978_5825# a_14946_4905# 0
C2581 a_2313_1791# VGND 0.01474f
C2582 a_4576_5047# a_4159_5303# 0.03016f
C2583 a_7845_5295# sky130_fd_sc_hd__mux2_1_0.S 0.13855f
C2584 a_13732_1769# VPWR 0.20646f
C2585 a_4627_12141# a_4505_13107# 0.00144f
C2586 a_6087_14735# a_6329_12927# 0
C2587 a_12994_4589# a_13175_4955# 0
C2588 a_14255_1769# a_15071_1765# 0
C2589 a_15227_5715# w_14736_5374# 0.10454f
C2590 a_7869_2145# sky130_fd_sc_hd__inv_1_0.A 0
C2591 a_15113_5459# A 0
C2592 a_6885_1783# a_8232_2145# 0.03325f
C2593 a_24241_14651# a_23731_14309# 0.02645f
C2594 w_12866_5378# A 0.00618f
C2595 a_17339_4938# sky130_fd_sc_hd__mux2_1_0.S 0.00688f
C2596 a_7845_5295# a_7899_5039# 0.00386f
C2597 a_10813_13753# a_12075_13379# 0
C2598 VGND w_9492_12311# 0.11704f
C2599 a_9599_10561# w_9502_10747# 0.05631f
C2600 ena clk 0.03102f
C2601 a_10857_14747# a_9865_15329# 0
C2602 a_11051_11919# VGND 0.00568f
C2603 a_4849_11293# w_5906_12121# 0.0984f
C2604 a_4903_15345# VGND 0.98587f
C2605 a_6885_1783# w_5454_1698# 0.02026f
C2606 a_10569_1777# a_11553_2139# 0.04534f
C2607 VGND a_23677_14701# 0.00402f
C2608 a_9875_13765# a_11091_12911# 0
C2609 a_9280_5471# w_9180_5386# 0.01793f
C2610 a_10046_2143# sky130_fd_sc_hd__inv_1_0.A 0
C2611 a_13439_4589# sky130_fd_sc_hd__inv_1_0.A 0
C2612 a_11385_2139# VGND 0.00231f
C2613 a_4213_5047# a_4159_5303# 0.00386f
C2614 a_7701_1779# a_7815_2035# 0
C2615 a_13357_5719# w_12866_5378# 0.10454f
C2616 a_4903_15345# a_6635_15235# 0
C2617 a_15113_5825# A 0
C2618 a_12509_4593# a_12994_4589# 0.02709f
C2619 a_2289_5307# a_2343_5051# 0.00386f
C2620 a_6329_12927# a_7113_13395# 0
C2621 a_4763_14775# w_4440_14739# 0.01327f
C2622 a_9465_16323# VPWR 0.3941f
C2623 a_10813_13753# a_12631_13987# 0
C2624 a_12966_5463# a_11541_5723# 0
C2625 a_7506_5013# a_7454_5039# 0.1439f
C2626 a_10450_4597# sky130_fd_sc_hd__inv_1_0.A 0
C2627 a_6029_5043# Y 0
C2628 a_4627_12141# w_5906_12121# 0
C2629 a_9801_12841# VGND 1.32139f
C2630 a_4847_14525# a_6805_15235# 0.00624f
C2631 sky130_fd_sc_hd__inv_1_5.Y ui_in[0] 0.06787f
C2632 a_14916_4559# a_13385_4845# 0.00446f
C2633 a_9801_12841# a_9799_16073# 0.4639f
C2634 a_11230_4567# a_11202_5441# 0
C2635 a_15309_4951# A 0
C2636 a_11049_14719# w_10748_13967# 0
C2637 a_14325_4589# a_14136_4955# 0
C2638 a_5999_2149# VGND 0.20086f
C2639 a_4905_12113# w_5910_13141# 0
C2640 a_11499_2029# a_11553_1773# 0.00386f
C2641 a_4913_13781# a_5809_14763# 0
C2642 a_11291_12911# a_11351_13753# 0.20048f
C2643 w_5484_4958# a_5636_5017# 0.05213f
C2644 Y w_3668_4962# 0.00346f
C2645 a_9465_16323# sky130_fd_sc_hd__inv_1_2.A 0
C2646 a_13243_1743# VPWR 0.97021f
C2647 a_8755_1779# w_7324_1694# 0.01935f
C2648 a_4213_5413# a_3229_5051# 0.04534f
C2649 a_2049_1791# a_2313_1791# 0
C2650 a_12481_5467# a_13285_5437# 0.02844f
C2651 a_24241_14651# A 0.03341f
C2652 a_6003_11935# a_4839_12857# 0
C2653 a_13046_4563# a_11569_4849# 0.00492f
C2654 VGND a_4755_13107# 0.02544f
C2655 a_4635_13809# a_4847_14525# 0
C2656 a_14297_5463# VPWR 1.06327f
C2657 a_6862_13645# VPWR 0.09661f
C2658 VGND w_1798_4966# 0.29762f
C2659 a_4905_12113# a_4515_11543# 0
C2660 a_16871_4938# VPWR 0.07431f
C2661 a_6862_13645# a_6944_13645# 0.00477f
C2662 a_4905_12113# w_4442_11507# 0.00119f
C2663 sky130_fd_sc_hd__inv_1_0.Y w_3638_1702# 0.00351f
C2664 a_4915_10549# a_4905_12113# 0.0298f
C2665 a_15255_4841# sky130_fd_sc_hd__mux2_1_0.VPB 0.00175f
C2666 a_13018_5437# w_12894_4504# 0
C2667 a_9557_14759# VGND 0.00172f
C2668 a_4913_13781# a_6127_13769# 0
C2669 w_4528_15559# VPWR 0.18191f
C2670 a_10937_12911# VPWR 0.1592f
C2671 a_9801_12841# w_9394_13055# 0.02723f
C2672 a_4915_10549# a_9717_13091# 0
C2673 VGND ua[0] 0.06916f
C2674 a_9811_11277# w_9402_14723# 0.00324f
C2675 a_6862_13645# a_6281_11907# 0.00248f
C2676 a_14794_1765# VGND 0.08635f
C2677 a_10422_5471# A 0
C2678 w_4530_12327# a_4905_12113# 0.0247f
C2679 w_12566_13951# a_12075_13379# 0.04664f
C2680 a_15644_5825# a_14297_5463# 0.03325f
C2681 a_4576_5413# VGND 0.18649f
C2682 a_12439_1773# w_11008_1688# 0.01094f
C2683 a_3199_1791# w_3638_1702# 0.25055f
C2684 w_11718_13593# a_11351_13753# 0.06723f
C2685 a_15017_5825# a_14836_5459# 0
C2686 uo_out[0] uio_in[7] 0.03102f
C2687 sky130_fd_sc_hd__mux2_1_0.VPB VGND 0.01288f
C2688 w_4432_13071# a_5975_12927# 0
C2689 a_4129_2043# w_5454_1698# 0
C2690 a_14946_4905# A 0.01569f
C2691 VGND a_5903_5017# 0.61211f
C2692 a_9715_16073# VPWR 0.00472f
C2693 w_7354_4954# a_6915_5043# 0.25055f
C2694 a_9238_1777# w_9138_1692# 0.01793f
C2695 a_5975_5299# VPWR 0.34516f
C2696 a_7869_2145# w_7324_1694# 0
C2697 a_9597_13793# a_9811_11277# 0.00317f
C2698 w_12566_13951# a_12631_13987# 0.05168f
C2699 w_12866_5378# a_14836_5459# 0.00188f
C2700 uio_in[1] uio_in[0] 0.03102f
C2701 a_13357_5719# a_14946_4905# 0
C2702 a_14888_5433# A 0.00509f
C2703 a_9877_10533# a_11824_13629# 0
C2704 a_11427_5467# VPWR 0.00102f
C2705 w_7604_13967# VGND 0.00757f
C2706 a_3790_1761# a_3738_1787# 0.1439f
C2707 a_24241_14651# a_24318_14385# 0.01352f
C2708 a_14255_1769# a_14794_1765# 0.0725f
C2709 w_11078_4508# a_11541_5723# 0
C2710 a_11623_4959# VPWR 0.00948f
C2711 a_10569_1777# a_11553_1773# 0.08312f
C2712 a_11553_2139# a_11289_2139# 0
C2713 a_10116_4963# VPWR 0.05672f
C2714 a_14946_4905# sky130_fd_sc_hd__mux2_1_0.A0 0.01594f
C2715 a_9597_13793# a_7113_13395# 0
C2716 a_7635_5405# VGND 0.00305f
C2717 a_10422_5837# A 0
C2718 a_6087_14735# a_4837_16089# 0.29394f
C2719 a_13357_5719# a_14888_5433# 0.00446f
C2720 a_6029_5409# a_6392_5409# 0.00847f
C2721 w_10872_13125# a_11243_11891# 0
C2722 w_12866_5378# a_13774_5463# 0.01154f
C2723 a_7899_5405# VPWR 0.00948f
C2724 Y a_2289_5307# 0.25757f
C2725 a_9489_4963# a_9753_4963# 0
C2726 a_8113_13753# w_11532_15433# 0.097f
C2727 a_9238_1777# sky130_fd_sc_hd__inv_1_0.A 0.00119f
C2728 a_9671_5727# a_10422_5471# 0.00682f
C2729 a_2289_5307# a_1950_5025# 0.04737f
C2730 a_4915_10549# a_7173_15235# 0.07716f
C2731 sky130_fd_sc_hd__mux2_1_0.A1 sky130_fd_sc_hd__inv_1_0.A 0
C2732 a_9699_4853# a_9725_5471# 0
C2733 VPWR a_10088_5471# 0.2062f
C2734 a_15141_4951# A 0
C2735 a_9809_14509# w_9392_16287# 0
C2736 a_3820_5021# w_1798_4966# 0
C2737 a_11019_12911# a_10937_12911# 0.00517f
C2738 w_5484_4958# a_6915_5043# 0.02026f
C2739 a_3199_1791# sky130_fd_sc_hd__inv_1_0.Y 0.0046f
C2740 a_9865_15329# VGND 0.98587f
C2741 a_9865_15329# a_9799_16073# 0.50561f
C2742 a_11986_4593# VGND 0.01315f
C2743 a_9489_4597# VGND 0
C2744 a_13105_1769# VPWR 0.00117f
C2745 a_10046_1777# w_9138_1692# 0.01154f
C2746 w_5712_14949# a_7173_15235# 0
C2747 a_2049_2157# VPWR 0
C2748 a_9465_16323# a_9715_16323# 0.02504f
C2749 a_8262_5405# w_7354_4954# 0.00139f
C2750 a_9360_4571# a_9585_4963# 0.00559f
C2751 a_4837_16089# a_7113_13395# 0
C2752 a_4721_13809# VPWR 0.003f
C2753 a_15281_5459# A 0
C2754 a_4849_11293# w_5910_13141# 0.05304f
C2755 a_9360_4571# w_7354_4954# 0
C2756 a_9597_13793# w_10748_13967# 0
C2757 a_9699_4853# VGND 1.17357f
C2758 uio_out[6] uio_out[7] 0.03102f
C2759 sky130_fd_sc_hd__inv_1_5.Y sky130_fd_sc_hd__inv_1_0.A 0
C2760 a_9589_12125# a_9597_13793# 0
C2761 a_12509_4593# w_12894_4504# 0.0025f
C2762 sky130_fd_sc_hd__mux2_1_0.S A 0.02419f
C2763 ui_in[0] a_24234_14385# 0.34724f
C2764 a_4159_5303# w_3668_4962# 0.10454f
C2765 a_2175_5417# VGND 0.0024f
C2766 a_2145_1791# a_2313_1791# 0
C2767 a_7899_5039# A 0
C2768 sky130_fd_sc_hd__inv_1_0.Y a_2313_1791# 0.08436f
C2769 a_3738_1787# VPWR 0.07401f
C2770 a_6885_1783# a_8755_1779# 0
C2771 a_7701_1779# VGND 0
C2772 a_4849_11293# a_4515_11543# 0.16782f
C2773 w_11050_5382# a_13018_5437# 0
C2774 a_4849_11293# w_4442_11507# 0.02399f
C2775 a_6392_5043# a_6915_5043# 0
C2776 a_5584_5043# a_5636_5017# 0.1439f
C2777 a_11597_15219# w_11718_13593# 0
C2778 a_4849_11293# a_4915_10549# 0.00639f
C2779 a_4847_14525# a_5809_14763# 0.00524f
C2780 a_4753_16339# a_4503_16339# 0.02504f
C2781 a_13357_5719# sky130_fd_sc_hd__mux2_1_0.S 0
C2782 a_10422_5837# a_9671_5727# 0.00696f
C2783 a_4129_2043# a_4546_2153# 0.06611f
C2784 w_5786_13983# a_4915_10549# 0
C2785 VGND a_11916_2139# 0.1864f
C2786 a_13147_5463# VGND 0
C2787 a_4905_12113# a_4839_12857# 0.04364f
C2788 a_10046_1777# sky130_fd_sc_hd__inv_1_0.A 0
C2789 a_14946_4905# a_14836_5459# 0.00175f
C2790 a_4129_2043# a_4880_2153# 0.00696f
C2791 a_9683_1777# a_9629_2033# 0.00386f
C2792 a_14916_4559# sky130_fd_sc_hd__inv_1_0.A 0
C2793 a_4849_11293# w_5712_14949# 0.08584f
C2794 a_4849_11293# w_4530_12327# 0.00145f
C2795 sky130_fd_sc_hd__mux2_1_0.A0 sky130_fd_sc_hd__mux2_1_0.S 0.1717f
C2796 w_11050_5382# a_11202_5441# 0.05213f
C2797 a_6389_13769# a_7173_15235# 0.00152f
C2798 a_7845_5295# a_10116_4963# 0
C2799 Y a_4910_5047# 0
C2800 Y w_5484_4958# 0.00152f
C2801 a_4627_12141# a_4515_11543# 0
C2802 a_2676_1791# VGND 0.01464f
C2803 a_6087_14735# a_5851_13769# 0
C2804 a_4627_12141# w_4442_11507# 0.00155f
C2805 a_9332_5445# a_9308_4597# 0
C2806 a_8113_13753# a_7173_15235# 0.00434f
C2807 a_13018_5437# VPWR 0.28383f
C2808 a_15045_4951# VPWR 0
C2809 w_9402_14723# a_9725_14759# 0.01327f
C2810 a_16006_4585# sky130_fd_sc_hd__inv_1_0.A 0
C2811 a_14888_5433# a_14836_5459# 0.1439f
C2812 a_2175_5051# a_2343_5051# 0
C2813 a_7899_5405# a_7845_5295# 0.03622f
C2814 a_7869_2145# a_7701_2145# 0
C2815 a_14864_4585# a_14946_4905# 0.07951f
C2816 a_15309_4951# w_14764_4500# 0
C2817 a_11243_11891# a_10937_12911# 0
C2818 a_7845_5295# a_10088_5471# 0
C2819 a_9597_13793# a_9683_13793# 0.00658f
C2820 a_4627_12141# w_4530_12327# 0.05631f
C2821 sky130_fd_sc_hd__inv_1_0.Y a_5999_2149# 0
C2822 a_11202_5441# VPWR 0.30708f
C2823 sky130_fd_sc_hd__inv_1_0.A a_14975_2131# 0
C2824 a_9671_5727# sky130_fd_sc_hd__mux2_1_0.S 0
C2825 a_10611_5471# VGND 0.69145f
C2826 a_11553_2139# VGND 0.20244f
C2827 a_10569_1777# a_9629_2033# 0.13962f
C2828 a_12481_5467# a_12292_5833# 0
C2829 a_5851_13769# a_7113_13395# 0
C2830 a_5636_5017# VPWR 0.29509f
C2831 a_7605_2145# a_7424_1779# 0
C2832 VPWR a_23511_14335# 0.00214f
C2833 a_7869_2145# a_6885_1783# 0.04534f
C2834 a_23511_14335# sky130_fd_sc_hd__mux4_1_0.VPB 0.00324f
C2835 a_9238_1777# w_7324_1694# 0.00227f
C2836 a_11049_14719# a_11351_13753# 0.00427f
C2837 a_9597_13793# a_9725_14759# 0
C2838 w_10872_13125# a_9811_11277# 0.05304f
C2839 a_14864_4585# a_14888_5433# 0
C2840 a_4765_11543# VGND 0.02702f
C2841 a_4849_11293# a_6389_13769# 0.00488f
C2842 a_6389_13769# w_5786_13983# 0.01492f
C2843 w_11050_5382# a_11595_5467# 0.01092f
C2844 sky130_fd_sc_hd__inv_1_2.A a_23511_14335# 0.04403f
C2845 a_8232_2145# VPWR 0.01966f
C2846 a_4513_14775# a_4849_11293# 0.00146f
C2847 VGND a_4753_16089# 0.00773f
C2848 a_2706_5417# w_1798_4966# 0.00139f
C2849 a_4763_14775# a_4625_15373# 0
C2850 a_9753_4963# VGND 0.19554f
C2851 a_9467_13091# a_9475_14759# 0
C2852 w_5454_1698# VPWR 0.51609f
C2853 a_12924_1769# sky130_fd_sc_hd__inv_1_0.A 0.00116f
C2854 a_9727_11527# VGND 0.02702f
C2855 a_13732_1769# a_13315_2025# 0.03016f
C2856 uio_out[1] uio_out[0] 0.03102f
C2857 a_4839_12857# a_7173_15235# 0.00685f
C2858 VGND a_12075_13379# 0.34868f
C2859 a_12075_13379# a_9799_16073# 0
C2860 a_9515_2143# VGND 0.00231f
C2861 a_14136_4589# VGND 0
C2862 a_23677_14335# a_23511_14335# 0.00648f
C2863 a_4713_12141# VPWR 0.00297f
C2864 a_14946_4905# w_14764_4500# 0.28173f
C2865 a_11595_5467# VPWR 0.17063f
C2866 a_4849_11293# a_4597_11543# 0
C2867 a_14066_2135# VGND 0.00244f
C2868 a_4837_16089# a_6805_15235# 0
C2869 a_13175_4955# VPWR 0
C2870 a_2343_5051# VPWR 0.17446f
C2871 ui_in[1] a_23511_14335# 0.01792f
C2872 a_5975_12927# VGND 0.14511f
C2873 a_9360_4571# a_9753_4597# 0.02283f
C2874 a_12250_2139# a_11499_2029# 0.00696f
C2875 VGND a_12631_13987# 0.24002f
C2876 a_14888_5433# w_14764_4500# 0
C2877 sky130_fd_sc_hd__inv_1_0.A a_24234_14385# 0.04346f
C2878 a_9547_16323# VGND 0.00117f
C2879 w_11718_13593# a_11291_12911# 0.04962f
C2880 a_11569_4849# sky130_fd_sc_hd__mux2_1_0.S 0
C2881 a_9547_16323# a_9799_16073# 0
C2882 VPWR a_13243_5829# 0
C2883 a_9877_10533# VPWR 0.59881f
C2884 w_6756_13609# VGND 0.01919f
C2885 sky130_fd_sc_hd__inv_1_2.Y a_4625_15373# 0
C2886 a_12509_4593# VPWR 0.06779f
C2887 a_10639_4597# sky130_fd_sc_hd__inv_1_0.A 0
C2888 a_14297_5463# A 0.00709f
C2889 a_4576_5047# a_3229_5051# 0.08907f
C2890 a_3010_1791# VGND 0
C2891 a_16871_4938# A 0.00367f
C2892 a_8113_13753# w_9392_16287# 0.00656f
C2893 a_15672_4951# a_14325_4589# 0.03325f
C2894 a_13315_2025# a_13243_1743# 0.21146f
C2895 a_4849_11293# a_4839_12857# 0.82158f
C2896 w_6756_13609# a_6635_15235# 0
C2897 a_14255_1769# a_14066_2135# 0
C2898 w_5786_13983# a_4839_12857# 0.08124f
C2899 a_6021_13769# VPWR 0
C2900 a_6087_14735# a_6862_13645# 0
C2901 a_15255_4841# a_15227_5715# 0.00177f
C2902 sky130_fd_sc_hd__inv_1_2.A a_9877_10533# 0.22585f
C2903 a_15672_4585# sky130_fd_sc_hd__inv_1_0.A 0
C2904 a_15644_5459# VPWR 0.2042f
C2905 a_14325_4589# sky130_fd_sc_hd__mux2_1_0.A1 0.00122f
C2906 a_9811_11277# a_10937_12911# 0.18651f
C2907 a_4910_5047# a_4159_5303# 0.00682f
C2908 a_4913_13781# a_4847_14525# 0.0012f
C2909 a_13357_5719# a_14297_5463# 0.13962f
C2910 w_5484_4958# a_4159_5303# 0
C2911 VPWR w_10868_12105# 0.07869f
C2912 a_13313_4563# a_13411_5463# 0
C2913 a_12439_1773# VPWR 0.06764f
C2914 a_2175_5051# a_1950_5025# 0.00487f
C2915 a_15071_2131# a_15185_2021# 0
C2916 a_4213_5047# a_3229_5051# 0.08312f
C2917 a_7605_2145# sky130_fd_sc_hd__inv_1_0.A 0
C2918 a_3949_5413# VPWR 0
C2919 a_4627_12141# a_4839_12857# 0
C2920 a_6915_5043# VPWR 1.05198f
C2921 a_11553_1773# VGND 0.01595f
C2922 a_9599_10561# a_9685_10561# 0.00658f
C2923 a_11597_15219# a_11049_14719# 0.08954f
C2924 VPWR a_9475_14759# 0.3877f
C2925 a_9801_12841# a_9557_14759# 0
C2926 a_14136_4955# VPWR 0
C2927 sky130_fd_sc_hd__inv_1_5.VPB VPWR 0.06925f
C2928 a_9557_5837# a_9725_5837# 0
C2929 sky130_fd_sc_hd__mux2_1_0.A0 a_14297_5463# 0
C2930 a_15309_4585# w_14764_4500# 0.01092f
C2931 a_15227_5715# VGND 1.19394f
C2932 a_12924_1769# a_12976_1743# 0.1439f
C2933 a_6862_13645# a_7113_13395# 0.10945f
C2934 Y a_5584_5043# 0.0012f
C2935 a_16871_4938# sky130_fd_sc_hd__mux2_1_0.A0 0.08041f
C2936 a_9877_10533# a_12809_13987# 0
C2937 a_13271_4589# a_13313_4563# 0
C2938 VGND a_9587_15357# 0.24327f
C2939 a_9332_5445# a_9725_5471# 0.02283f
C2940 w_4430_16303# sky130_fd_sc_hd__inv_1_2.Y 0
C2941 a_9799_16073# a_9587_15357# 0
C2942 a_5975_5299# A 0.00228f
C2943 VGND a_4213_5413# 0.20073f
C2944 a_6392_5409# w_5484_4958# 0.00139f
C2945 sky130_fd_sc_hd__mux2_1_0.S w_14764_4500# 0.0011f
C2946 a_15141_4585# a_15309_4585# 0
C2947 a_11331_5467# VPWR 0.00136f
C2948 a_4513_14775# w_4440_14739# 0.06993f
C2949 a_11499_2029# sky130_fd_sc_hd__inv_1_0.A 0.00294f
C2950 w_4432_13071# a_4905_12113# 0
C2951 a_4503_16339# a_4847_14525# 0
C2952 a_4637_10577# a_4515_11543# 0.00144f
C2953 a_4637_10577# w_4442_11507# 0
C2954 a_9683_1777# w_9138_1692# 0.01092f
C2955 a_5999_1783# w_5454_1698# 0.01092f
C2956 a_4637_10577# a_4915_10549# 0.1296f
C2957 a_10611_5471# a_11541_5723# 0.21188f
C2958 a_13439_4589# w_12894_4504# 0.01092f
C2959 a_4546_2153# VPWR 0.01963f
C2960 a_11049_14719# a_10771_14747# 0.1109f
C2961 a_11427_5467# A 0
C2962 w_4538_13995# a_4505_13107# 0
C2963 a_9461_5471# a_9725_5471# 0
C2964 a_11623_4959# A 0
C2965 a_13774_5829# VPWR 0.01982f
C2966 a_4880_2153# VPWR 0
C2967 a_9332_5445# VGND 0.51815f
C2968 a_10116_4963# A 0
C2969 a_11986_4593# w_11078_4508# 0.01154f
C2970 a_4635_13809# a_5851_13769# 0
C2971 a_13802_4589# VGND 0.01131f
C2972 a_24407_14651# a_24774_14701# 0
C2973 a_14325_4589# a_14916_4559# 0.11887f
C2974 a_14975_1765# sky130_fd_sc_hd__inv_1_0.A 0
C2975 a_15071_2131# sky130_fd_sc_hd__inv_1_0.A 0
C2976 a_11553_1773# a_11385_1773# 0
C2977 VGND a_9461_5471# 0
C2978 a_9875_13765# a_11824_13629# 0
C2979 a_9699_4853# w_11078_4508# 0
C2980 a_7899_5405# A 0
C2981 sky130_fd_sc_hd__inv_1_0.Y a_2676_1791# 0.08982f
C2982 w_10748_13967# a_10937_12911# 0
C2983 a_4763_14775# VPWR 0.32009f
C2984 w_6570_15449# VGND 0.00665f
C2985 a_10569_1777# w_9138_1692# 0.02026f
C2986 Y VPWR 1.29284f
C2987 a_10088_5471# A 0
C2988 a_11178_4593# a_10639_4597# 0.0725f
C2989 a_8262_5405# VPWR 0.01999f
C2990 uio_in[6] uio_in[7] 0.03102f
C2991 a_5933_13769# a_4913_13781# 0
C2992 sky130_fd_sc_hd__inv_1_4.A VGND 0.25634f
C2993 a_9867_12097# a_11091_12911# 0
C2994 a_9683_1777# sky130_fd_sc_hd__inv_1_0.A 0
C2995 a_1950_5025# VPWR 0.30536f
C2996 a_15185_2021# a_15936_1765# 0.00682f
C2997 a_9360_4571# VPWR 0.39467f
C2998 uio_out[4] uio_out[5] 0.03102f
C2999 w_6570_15449# a_6635_15235# 0.08205f
C3000 a_13175_4589# VPWR 0.00118f
C3001 a_6029_5043# a_5861_5043# 0
C3002 a_3040_5051# VGND 0
C3003 a_3199_1791# a_2676_1791# 0
C3004 w_4440_14739# a_4839_12857# 0.00408f
C3005 a_14297_5463# a_14836_5459# 0.0725f
C3006 a_4015_2153# a_4183_2153# 0
C3007 a_12924_1769# a_13105_2135# 0
C3008 a_6003_11935# VGND 0.13487f
C3009 a_7845_5295# a_6915_5043# 0.21188f
C3010 a_13018_5437# a_13147_5829# 0.00792f
C3011 VGND sky130_fd_sc_hd__inv_1_2.VPB 0.01278f
C3012 a_4847_14525# a_6717_15235# 0.00159f
C3013 sky130_fd_sc_hd__inv_1_5.Y a_24962_14701# 0
C3014 a_7424_1779# a_5945_2039# 0
C3015 a_13732_1769# w_12824_1684# 0.01154f
C3016 a_11623_4593# a_10639_4597# 0.08312f
C3017 VPWR w_9180_5386# 0.52056f
C3018 a_6911_15235# a_7173_15235# 0
C3019 VPWR a_15602_1765# 0.2057f
C3020 a_10965_11919# w_10872_13125# 0
C3021 a_9801_12841# a_9865_15329# 0.1369f
C3022 w_14694_1680# a_15185_2021# 0.10454f
C3023 VGND a_11679_15219# 0.00151f
C3024 a_9799_16073# a_11679_15219# 0
C3025 a_5099_5047# w_3668_4962# 0.01094f
C3026 VGND a_4045_5413# 0.00231f
C3027 a_11359_4593# sky130_fd_sc_hd__inv_1_0.A 0
C3028 a_9599_10561# VGND 0.24388f
C3029 w_9500_13979# a_9475_14759# 0.0035f
C3030 a_10569_1777# sky130_fd_sc_hd__inv_1_0.A 0.00267f
C3031 a_4837_16089# a_5809_14763# 0.03093f
C3032 a_8755_1779# VPWR 1.04258f
C3033 a_9465_16323# a_9725_14759# 0
C3034 a_23731_14309# a_23511_14335# 0.0457f
C3035 a_11499_2029# a_12976_1743# 0.00492f
C3036 a_4505_13107# VPWR 0.38927f
C3037 sky130_fd_sc_hd__inv_1_2.Y VPWR 1.38991f
C3038 a_3820_5021# a_4213_5413# 0.02301f
C3039 a_7454_5039# a_5975_5299# 0
C3040 a_2676_1791# a_2313_1791# 0.00985f
C3041 a_13774_5463# a_14297_5463# 0
C3042 a_12250_1773# VPWR 0
C3043 a_4913_13781# a_6329_12927# 0.0204f
C3044 a_7476_1753# w_5454_1698# 0
C3045 a_8262_5039# VGND 0.01509f
C3046 a_9629_2033# VGND 1.19975f
C3047 a_7815_2035# w_9138_1692# 0
C3048 a_13271_4589# a_13046_4563# 0.00487f
C3049 sky130_fd_sc_hd__inv_1_0.A a_15936_1765# 0
C3050 w_11078_4508# a_10611_5471# 0
C3051 sky130_fd_sc_hd__inv_1_5.VPB sky130_fd_sc_hd__inv_1_5.A 0.05645f
C3052 a_11049_14719# a_11291_12911# 0
C3053 sky130_fd_sc_hd__inv_1_2.A sky130_fd_sc_hd__inv_1_2.Y 0.10747f
C3054 a_9671_5727# a_10088_5471# 0.03016f
C3055 a_9557_14759# a_9865_15329# 0
C3056 a_4837_16089# a_6127_13769# 0.00702f
C3057 sky130_fd_sc_hd__inv_1_5.Y a_24774_14701# 0
C3058 a_9877_10533# a_11243_11891# 0.44698f
C3059 a_13018_5437# A 0.00516f
C3060 a_10771_14747# w_9402_14723# 0
C3061 a_13046_4563# a_13313_4563# 0.11512f
C3062 a_14846_1739# a_15185_2021# 0.04737f
C3063 a_9809_14509# a_9467_13091# 0
C3064 VPWR a_9419_1777# 0.00114f
C3065 a_23511_14701# a_23511_14335# 0.00987f
C3066 ui_in[5] ui_in[4] 0.03102f
C3067 w_5906_12121# VPWR 0.07869f
C3068 a_13243_1743# w_12824_1684# 0.24672f
C3069 a_4159_5303# a_5584_5043# 0
C3070 a_9673_15357# VPWR 0.00333f
C3071 a_4183_1787# VGND 0.0153f
C3072 a_6057_12927# a_5975_12927# 0.00517f
C3073 a_8262_5405# a_7845_5295# 0.06611f
C3074 w_4432_13071# a_4849_11293# 0.00299f
C3075 w_14694_1680# sky130_fd_sc_hd__inv_1_0.A 0.02746f
C3076 a_11202_5441# A 0.00521f
C3077 a_13357_5719# a_13018_5437# 0.04737f
C3078 a_1898_5051# VPWR 0.08401f
C3079 a_7845_5295# a_9360_4571# 0
C3080 a_5735_1783# VGND 0
C3081 a_6281_11907# w_5906_12121# 0.02153f
C3082 a_3229_5051# w_3668_4962# 0.25055f
C3083 A a_23511_14335# 0.00544f
C3084 a_11243_11891# w_10868_12105# 0.02153f
C3085 a_7869_2145# VPWR 0.00911f
C3086 a_9308_4597# sky130_fd_sc_hd__inv_1_0.A 0
C3087 a_11553_2139# a_11385_2139# 0
C3088 a_7815_2035# sky130_fd_sc_hd__inv_1_0.A 0.00297f
C3089 a_14325_4589# w_14736_5374# 0.00258f
C3090 a_13385_4845# VGND 1.17207f
C3091 a_9875_13765# a_11089_13753# 0
C3092 VGND a_11906_13629# 0
C3093 a_3010_2157# VGND 0.00245f
C3094 a_11049_14719# w_11718_13593# 0
C3095 a_14297_5463# w_14764_4500# 0
C3096 sky130_fd_sc_hd__inv_1_0.Y a_3010_1791# 0
C3097 a_3768_5047# a_3949_5413# 0
C3098 a_3919_2153# VGND 0.00305f
C3099 a_9875_13765# a_9467_13091# 0
C3100 a_5945_2039# a_5873_1757# 0.21146f
C3101 a_11623_4959# a_11569_4849# 0.03622f
C3102 w_4432_13071# a_4627_12141# 0
C3103 a_12924_1769# w_11008_1688# 0.00227f
C3104 a_12135_15219# VPWR 0.55326f
C3105 a_10046_2143# VPWR 0.01966f
C3106 a_7845_5295# w_9180_5386# 0
C3107 a_15672_4585# a_14325_4589# 0.08907f
C3108 a_15281_5825# w_14736_5374# 0
C3109 a_13439_4589# VPWR 0.17476f
C3110 w_10674_14933# a_9475_14759# 0
C3111 a_5851_13769# a_5809_14763# 0
C3112 uo_out[5] uo_out[6] 0.03102f
C3113 a_10965_11919# a_10937_12911# 0
C3114 a_16006_4951# VPWR 0
C3115 a_14846_1739# sky130_fd_sc_hd__inv_1_0.A 0.00279f
C3116 w_12866_5378# a_13411_5463# 0.01092f
C3117 a_1868_1791# VGND 0.09509f
C3118 a_3820_5021# a_4045_5413# 0.00559f
C3119 a_13732_1769# a_13369_1769# 0.00985f
C3120 sky130_fd_sc_hd__inv_1_2.A a_12135_15219# 0.04463f
C3121 a_4637_10577# a_4723_10577# 0.00658f
C3122 a_10450_4597# VPWR 0
C3123 a_5945_2039# sky130_fd_sc_hd__inv_1_0.A 0.00224f
C3124 VGND ui_in[0] 0.53405f
C3125 a_4159_5303# VPWR 0.34536f
C3126 a_11767_15219# VPWR 0.00151f
C3127 a_5069_1787# VGND 0.06388f
C3128 a_9467_13091# w_9404_11491# 0
C3129 a_11595_5467# A 0
C3130 a_6362_1783# a_5945_2039# 0.03016f
C3131 a_5851_13769# a_6127_13769# 0.00119f
C3132 VGND a_13285_5437# 0.66733f
C3133 sky130_fd_sc_hd__inv_1_4.A sky130_fd_sc_hd__inv_1_4.VPB 0.05681f
C3134 a_9671_5727# a_11202_5441# 0.00446f
C3135 a_11289_2139# sky130_fd_sc_hd__inv_1_0.A 0
C3136 w_12866_5378# a_13313_4563# 0.00258f
C3137 a_6392_5409# VPWR 0.01964f
C3138 a_14916_4559# w_12894_4504# 0
C3139 a_4903_15345# a_5975_12927# 0
C3140 a_9809_14509# VPWR 0.3635f
C3141 a_11623_4593# a_11359_4593# 0
C3142 a_9801_12841# a_12075_13379# 0.00444f
C3143 a_9725_14509# a_9475_14759# 0.00723f
C3144 a_7424_1779# VGND 0.08651f
C3145 a_24962_14701# a_24234_14385# 0.1456f
C3146 a_4753_16339# a_4837_16089# 0.07445f
C3147 a_13243_5829# A 0
C3148 a_11873_15219# a_12135_15219# 0
C3149 a_4905_12113# VGND 0.43935f
C3150 a_3768_5047# Y 0.00167f
C3151 a_7669_14003# a_4915_10549# 0.07457f
C3152 a_7731_5039# VPWR 0
C3153 a_12509_4593# A 0
C3154 a_4755_12857# a_4505_13107# 0.00723f
C3155 VGND a_9717_13091# 0.02544f
C3156 a_6129_12927# a_4839_12857# 0.00312f
C3157 w_11532_15433# VGND 0.00665f
C3158 w_11532_15433# a_9799_16073# 0.09702f
C3159 a_15045_4585# a_15309_4585# 0
C3160 a_4915_10549# a_9467_13091# 0.00237f
C3161 a_13369_1769# a_13243_1743# 0.08094f
C3162 a_9811_11277# a_9877_10533# 0.00639f
C3163 a_5765_5043# a_5636_5017# 0.00758f
C3164 VPWR VPB 0.06609f
C3165 a_9801_12841# a_12631_13987# 0
C3166 Y a_4910_5413# 0
C3167 VGND a_11091_12911# 0.00291f
C3168 a_13243_5463# a_13018_5437# 0.00487f
C3169 a_24407_14651# VPWR 0.00288f
C3170 a_13357_5719# a_13243_5829# 0
C3171 a_15644_5459# A 0
C3172 a_2289_5307# a_3229_5051# 0.13962f
C3173 a_4837_16089# a_4913_13781# 0.01745f
C3174 a_9875_13765# VPWR 0.60287f
C3175 VPWR sky130_fd_sc_hd__inv_1_3.VPB 0.07652f
C3176 Y a_2343_5417# 0.0517f
C3177 a_9725_5837# VPWR 0.00613f
C3178 a_4513_14775# a_4625_15373# 0
C3179 a_2343_5417# a_1950_5025# 0.02301f
C3180 a_5099_5047# w_5484_4958# 0.0025f
C3181 a_6915_5043# A 0.00267f
C3182 uio_oe[4] uio_oe[3] 0.03102f
C3183 a_12250_2139# VGND 0.00244f
C3184 a_7815_2035# w_7324_1694# 0.10454f
C3185 a_24774_14701# a_24234_14385# 0.17579f
C3186 a_4635_13809# a_4721_13809# 0.00658f
C3187 a_4183_1787# w_3638_1702# 0.01092f
C3188 a_11499_2029# w_11008_1688# 0.10454f
C3189 a_8755_1779# a_9515_1777# 0
C3190 a_14864_4585# a_15045_4951# 0
C3191 a_9811_11277# w_10868_12105# 0.0984f
C3192 w_9394_13055# a_9717_13091# 0.01327f
C3193 a_11331_5833# VGND 0.00311f
C3194 a_15185_2021# VGND 1.19592f
C3195 a_8232_1779# a_8755_1779# 0
C3196 a_4837_16089# a_4503_16339# 0.16891f
C3197 a_11331_5467# A 0
C3198 a_9811_11277# a_9475_14759# 0.00146f
C3199 a_11230_4567# a_10639_4597# 0.11887f
C3200 a_5606_1757# a_5554_1783# 0.1439f
C3201 VPWR w_9404_11491# 0.16044f
C3202 a_15644_5459# sky130_fd_sc_hd__mux2_1_0.A0 0
C3203 a_14297_5463# a_14108_5829# 0
C3204 VGND w_9138_1692# 0.2932f
C3205 a_4576_5047# VGND 0.01333f
C3206 a_10569_1777# a_10380_2143# 0
C3207 a_15672_4951# VPWR 0.02182f
C3208 a_13774_5829# A 0.00188f
C3209 a_7669_14003# a_6389_13769# 0.00196f
C3210 a_11986_4593# a_10611_5471# 0
C3211 a_5945_2039# w_7324_1694# 0
C3212 a_13369_2135# a_13732_2135# 0.00847f
C3213 a_13369_2135# sky130_fd_sc_hd__inv_1_0.A 0
C3214 VPWR w_5910_13141# 0.0888f
C3215 a_8113_13753# a_7669_14003# 0.10318f
C3216 a_9238_1777# VPWR 0.07483f
C3217 a_15255_4841# sky130_fd_sc_hd__inv_1_0.A 0
C3218 a_11202_5441# a_11595_5833# 0.02301f
C3219 w_10748_13967# a_9877_10533# 0
C3220 a_24407_14651# ui_in[1] 0.00109f
C3221 a_4513_14775# w_4430_16303# 0
C3222 a_5873_1757# VGND 0.61194f
C3223 a_14946_4905# a_13313_4563# 0
C3224 a_9683_2143# a_8755_1779# 0.04534f
C3225 a_7635_5039# VPWR 0.00116f
C3226 a_10771_14747# w_10872_13125# 0
C3227 sky130_fd_sc_hd__mux2_1_0.A1 VPWR 0.2778f
C3228 a_15185_2021# a_15239_1765# 0.00386f
C3229 a_9699_4853# a_10611_5471# 0
C3230 w_11050_5382# a_12481_5467# 0.01094f
C3231 VGND a_7173_15235# 0.32171f
C3232 a_4213_5047# VGND 0.01521f
C3233 a_6281_11907# w_5910_13141# 0
C3234 a_14255_1769# a_15185_2021# 0.21188f
C3235 a_13357_5719# a_13774_5829# 0.06611f
C3236 a_7845_5295# a_7731_5039# 0
C3237 a_5069_1787# w_3638_1702# 0.01094f
C3238 w_6570_15449# a_4903_15345# 0
C3239 a_13046_4563# w_12866_5378# 0.00104f
C3240 a_4515_11543# VPWR 0.3853f
C3241 a_4513_14775# w_4538_13995# 0.0035f
C3242 Y A 0.11807f
C3243 VPWR w_4442_11507# 0.16044f
C3244 a_6635_15235# a_7173_15235# 0.08446f
C3245 a_4915_10549# VPWR 0.69549f
C3246 a_8262_5405# A 0
C3247 a_9477_11527# a_9877_10533# 0
C3248 a_13732_2135# VGND 0.18636f
C3249 VGND sky130_fd_sc_hd__inv_1_0.A 0.75219f
C3250 a_9360_4571# A 0
C3251 a_4913_13781# a_5851_13769# 0.0094f
C3252 sky130_fd_sc_hd__inv_1_5.Y VPWR 1.0628f
C3253 sky130_fd_sc_hd__inv_1_5.Y sky130_fd_sc_hd__mux4_1_0.VPB 0.10326f
C3254 a_12481_5467# VPWR 0.06365f
C3255 a_11986_4959# a_10639_4597# 0.03325f
C3256 a_12135_15219# a_11243_11891# 0.09936f
C3257 a_4183_1787# sky130_fd_sc_hd__inv_1_0.Y 0
C3258 a_6362_1783# VGND 0.01331f
C3259 a_9589_12125# w_10868_12105# 0
C3260 w_5712_14949# VPWR 0.0786f
C3261 a_11595_5467# a_11569_4849# 0
C3262 a_4915_10549# a_6281_11907# 0.43285f
C3263 a_11553_2139# a_11916_2139# 0.00847f
C3264 a_9865_15329# a_12075_13379# 0
C3265 w_4530_12327# VPWR 0.17848f
C3266 a_2313_2157# a_2676_2157# 0.00847f
C3267 a_9699_4853# a_9753_4963# 0.03622f
C3268 a_4837_16089# a_6717_15235# 0
C3269 w_10674_14933# a_12135_15219# 0
C3270 a_11541_5723# a_13285_5437# 0.00412f
C3271 ui_in[7] uio_in[0] 0.03102f
C3272 sky130_fd_sc_hd__inv_1_5.Y sky130_fd_sc_hd__inv_1_2.A 0.34711f
C3273 a_10569_1777# w_11008_1688# 0.25055f
C3274 a_7476_1753# a_7869_2145# 0.02301f
C3275 sky130_fd_sc_hd__inv_1_0.Y a_5735_1783# 0
C3276 a_2145_2157# VGND 0.0024f
C3277 a_9875_13765# w_9500_13979# 0.01958f
C3278 a_15239_2131# a_15185_2021# 0.03622f
C3279 A w_9180_5386# 0.0065f
C3280 a_4576_5413# a_4213_5413# 0.00847f
C3281 a_13105_1769# a_13369_1769# 0
C3282 a_12966_5463# a_13285_5437# 0.04799f
C3283 a_12881_13987# VPWR 0
C3284 a_4849_11293# VGND 1.26863f
C3285 a_7454_5039# a_6915_5043# 0.0725f
C3286 a_3199_1791# a_4183_1787# 0.08312f
C3287 a_3010_2157# sky130_fd_sc_hd__inv_1_0.Y 0
C3288 a_10046_1777# VPWR 0.20638f
C3289 w_5786_13983# VGND 0.01862f
C3290 a_10813_13753# a_11824_13629# 0
C3291 sky130_fd_sc_hd__inv_1_0.A a_15239_1765# 0
C3292 a_3919_2153# sky130_fd_sc_hd__inv_1_0.Y 0
C3293 a_8566_2145# a_8755_1779# 0
C3294 a_14916_4559# VPWR 0.31865f
C3295 a_4765_11293# a_4515_11543# 0.00723f
C3296 a_7669_14003# a_4839_12857# 0
C3297 a_14255_1769# sky130_fd_sc_hd__inv_1_0.A 0.00715f
C3298 sky130_fd_sc_hd__inv_1_5.Y a_23677_14335# 0
C3299 w_9208_4512# sky130_fd_sc_hd__mux2_1_0.S 0.00202f
C3300 sky130_fd_sc_hd__inv_1_2.A a_12881_13987# 0
C3301 sky130_fd_sc_hd__inv_1_5.A sky130_fd_sc_hd__inv_1_3.VPB 0
C3302 a_17053_4938# sky130_fd_sc_hd__mux2_1_0.S 0.00526f
C3303 a_9557_5471# a_9725_5471# 0
C3304 a_8596_5039# VGND 0
C3305 a_6029_5409# a_5765_5409# 0
C3306 a_12509_4593# a_11569_4849# 0.12975f
C3307 a_13385_4845# a_13411_5829# 0
C3308 a_10569_1777# a_11108_1773# 0.0725f
C3309 a_15978_5459# VPWR 0
C3310 ua[4] a_14975_1765# 0
C3311 a_6087_14735# sky130_fd_sc_hd__inv_1_2.Y 0.09734f
C3312 a_4910_5413# a_4159_5303# 0.00696f
C3313 a_11385_1773# sky130_fd_sc_hd__inv_1_0.A 0
C3314 a_10046_2143# a_9683_2143# 0.00847f
C3315 a_4627_12141# VGND 0.24254f
C3316 a_3010_2157# a_3199_1791# 0
C3317 a_1868_1791# sky130_fd_sc_hd__inv_1_0.Y 0.0073f
C3318 a_16006_4585# VPWR 0
C3319 a_13369_2135# a_12976_1743# 0.02301f
C3320 w_4538_13995# a_4839_12857# 0.00445f
C3321 a_2676_2157# w_1768_1706# 0.00139f
C3322 a_7701_2145# a_7815_2035# 0
C3323 sky130_fd_sc_hd__inv_1_5.Y ui_in[1] 0.02204f
C3324 a_13313_4563# sky130_fd_sc_hd__mux2_1_0.S 0.02903f
C3325 w_10674_14933# a_9809_14509# 0.00381f
C3326 a_24152_14385# a_24234_14385# 0.04662f
C3327 sky130_fd_sc_hd__inv_1_0.Y a_5069_1787# 0
C3328 a_6389_13769# VPWR 0.38708f
C3329 a_6389_13769# a_6944_13645# 0.00183f
C3330 a_9360_4571# a_9671_5727# 0
C3331 a_8113_13753# VPWR 2.11591f
C3332 a_13439_4955# VGND 0.19548f
C3333 VGND a_9557_5471# 0
C3334 a_12292_5833# VGND 0.00291f
C3335 VPWR a_14975_2131# 0
C3336 w_9502_10747# VPWR 0.166f
C3337 a_4513_14775# VPWR 0.38904f
C3338 a_11623_4959# a_11455_4959# 0
C3339 a_10771_14747# a_10937_12911# 0
C3340 a_2313_2157# VGND 0.19866f
C3341 a_9877_10533# a_12713_13987# 0
C3342 a_17339_4938# sky130_fd_sc_hd__mux2_1_0.A1 0
C3343 w_10872_13125# a_11291_12911# 0.02303f
C3344 a_4837_16089# a_4847_14525# 0.46421f
C3345 a_6389_13769# a_6281_11907# 0.00255f
C3346 a_4213_5047# a_3820_5021# 0.02283f
C3347 a_15239_2131# sky130_fd_sc_hd__inv_1_0.A 0.00137f
C3348 a_6885_1783# a_7815_2035# 0.21188f
C3349 a_4505_13107# a_4587_13107# 0.00641f
C3350 a_8113_13753# a_6281_11907# 0.00287f
C3351 a_5099_5047# a_5584_5043# 0.02709f
C3352 a_11230_4567# a_11359_4593# 0.00758f
C3353 Y a_5765_5043# 0
C3354 a_9875_13765# a_10895_13753# 0
C3355 a_8113_13753# sky130_fd_sc_hd__inv_1_2.A 0.16034f
C3356 uio_oe[5] uio_oe[6] 0.03102f
C3357 a_9280_5471# VGND 0.12844f
C3358 a_12976_1743# VGND 0.40116f
C3359 a_6029_5409# VGND 0.20237f
C3360 a_14946_4905# a_13046_4563# 0
C3361 a_9671_5727# w_9180_5386# 0.10454f
C3362 a_11178_4593# VGND 0.07994f
C3363 a_13411_5829# a_13285_5437# 0.04534f
C3364 a_4915_10549# w_9500_13979# 0.00206f
C3365 w_9392_16287# VGND 0.06272f
C3366 a_9308_4597# w_7354_4954# 0.00201f
C3367 a_5895_14763# a_4839_12857# 0
C3368 a_4597_11543# VPWR 0.02511f
C3369 w_9392_16287# a_9799_16073# 0.02445f
C3370 a_9865_15329# a_9587_15357# 0.12165f
C3371 w_10674_14933# a_9875_13765# 0
C3372 a_9559_11527# a_4915_10549# 0
C3373 a_9475_14759# a_9725_14759# 0.02504f
C3374 a_5873_1757# w_3638_1702# 0.00743f
C3375 a_10965_11919# a_9877_10533# 0
C3376 a_9809_14509# a_9725_14509# 0.00206f
C3377 a_12924_1769# VPWR 0.07454f
C3378 VGND w_7324_1694# 0.29306f
C3379 a_5735_2149# a_5606_1757# 0.00792f
C3380 a_4915_10549# a_9549_13091# 0
C3381 a_13802_4955# VGND 0.18285f
C3382 a_6885_1783# a_5945_2039# 0.13962f
C3383 a_12439_1773# w_12824_1684# 0.0025f
C3384 Y a_2079_5417# 0
C3385 a_5975_5299# a_6726_5409# 0.00696f
C3386 a_9875_13765# a_10983_13753# 0.00104f
C3387 VGND w_1768_1706# 0.29741f
C3388 a_4847_14525# a_4595_14775# 0
C3389 a_2079_5417# a_1950_5025# 0.00792f
C3390 sky130_fd_sc_hd__inv_1_5.Y sky130_fd_sc_hd__inv_1_5.A 0.15583f
C3391 a_11623_4593# VGND 0.01251f
C3392 a_16006_4951# A 0
C3393 a_6862_13645# a_4913_13781# 0
C3394 a_12135_15219# a_9811_11277# 0
C3395 a_6726_5043# VGND 0
C3396 a_9801_12841# a_11906_13629# 0
C3397 w_11050_5382# a_10639_4597# 0.00258f
C3398 a_5861_5043# VPWR 0
C3399 a_13369_2135# a_13105_2135# 0
C3400 ui_in[0] a_23677_14701# 0.0594f
C3401 a_4839_12857# VPWR 0.75065f
C3402 a_5099_5047# VPWR 0.06751f
C3403 w_4440_14739# VGND 0.07437f
C3404 a_6029_5043# VGND 0.01597f
C3405 a_10965_11919# w_10868_12105# 0.05631f
C3406 a_6944_13645# a_4839_12857# 0
C3407 a_10569_1777# a_11289_1773# 0
C3408 VGND a_4711_15373# 0.00661f
C3409 VPWR a_24234_14385# 0.22976f
C3410 a_5933_13769# a_4837_16089# 0
C3411 a_24234_14385# sky130_fd_sc_hd__mux4_1_0.VPB 0.05795f
C3412 a_10813_13753# a_11089_13753# 0.00119f
C3413 a_6281_11907# a_4839_12857# 0.02336f
C3414 VGND w_3668_4962# 0.29368f
C3415 a_14946_4905# a_15017_5825# 0
C3416 a_6392_5409# A 0
C3417 VPWR w_14736_5374# 0.5114f
C3418 a_5851_13769# a_4847_14525# 0
C3419 a_4503_16339# w_4528_15559# 0.0035f
C3420 a_10639_4597# VPWR 1.1195f
C3421 a_15185_2021# a_15071_1765# 0
C3422 a_11108_1773# a_11289_2139# 0
C3423 a_13105_2135# VGND 0.00305f
C3424 a_8113_13753# w_9500_13979# 0.00438f
C3425 a_12631_13987# a_12075_13379# 0.28206f
C3426 a_9809_14509# a_9811_11277# 0.00506f
C3427 a_15672_4585# VPWR 0.21095f
C3428 a_11291_12911# a_10937_12911# 0.09582f
C3429 a_4723_10577# VPWR 0.00176f
C3430 a_13046_4563# sky130_fd_sc_hd__mux2_1_0.S 0
C3431 a_15255_4841# a_14325_4589# 0.21188f
C3432 a_15113_5459# a_14946_4905# 0
C3433 a_14946_4905# w_12866_5378# 0
C3434 a_15017_5825# a_14888_5433# 0.00792f
C3435 a_7731_5039# A 0
C3436 sky130_fd_sc_hd__inv_1_0.Y a_5873_1757# 0.0011f
C3437 a_15644_5825# w_14736_5374# 0.00139f
C3438 VPB A 0.05211f
C3439 a_7605_1779# sky130_fd_sc_hd__inv_1_0.A 0
C3440 a_11623_4959# a_11359_4959# 0
C3441 a_4763_14775# a_4635_13809# 0
C3442 a_7605_2145# VPWR 0
C3443 a_12135_15219# w_10748_13967# 0
C3444 a_24407_14651# A 0
C3445 ua[4] a_14846_1739# 0
C3446 a_11958_5467# VGND 0.01767f
C3447 a_15255_4841# a_15281_5825# 0
C3448 a_11351_13753# a_9877_10533# 0.00262f
C3449 a_12881_13987# a_11243_11891# 0
C3450 a_15113_5459# a_14888_5433# 0.00487f
C3451 a_15113_5825# a_14946_4905# 0
C3452 w_12866_5378# a_14888_5433# 0
C3453 ui_in[0] ua[0] 0.53257f
C3454 a_10380_2143# VGND 0.00244f
C3455 a_13201_1769# sky130_fd_sc_hd__inv_1_0.A 0
C3456 VPWR a_3229_5051# 1.0518f
C3457 a_12292_5467# VPWR 0
C3458 a_14325_4589# VGND 0.07198f
C3459 a_9725_5837# A 0.0014f
C3460 a_3199_1791# a_5873_1757# 0
C3461 sky130_fd_sc_hd__inv_1_0.Y sky130_fd_sc_hd__inv_1_0.A 0.11803f
C3462 a_9717_12841# a_4915_10549# 0
C3463 a_9801_12841# a_9717_13091# 0.08134f
C3464 a_24234_14385# ui_in[1] 0.28582f
C3465 a_8113_13753# a_9715_16323# 0
C3466 a_7506_5013# a_7899_5039# 0.02283f
C3467 a_9875_13765# a_9811_11277# 0.26616f
C3468 a_11499_2029# VPWR 0.34562f
C3469 a_2079_5417# a_1898_5051# 0
C3470 a_12292_5833# a_11541_5723# 0.00696f
C3471 a_15309_4951# a_14946_4905# 0.19411f
C3472 a_4513_14775# a_4763_14525# 0.00723f
C3473 a_9801_12841# a_11091_12911# 0.00312f
C3474 a_15281_5825# VGND 0.20007f
C3475 a_4637_10577# VGND 0.2439f
C3476 a_15071_1765# sky130_fd_sc_hd__inv_1_0.A 0
C3477 sky130_fd_sc_hd__inv_1_5.Y a_23731_14309# 0.09059f
C3478 a_9725_14509# a_4915_10549# 0
C3479 a_15113_5825# a_14888_5433# 0.00559f
C3480 a_12994_4589# VGND 0.08826f
C3481 a_2145_2157# sky130_fd_sc_hd__inv_1_0.Y 0
C3482 a_5933_13769# a_5851_13769# 0.00578f
C3483 a_6057_12927# a_4849_11293# 0.00146f
C3484 a_4721_13809# a_4913_13781# 0.00222f
C3485 Y a_4045_5047# 0
C3486 a_7869_1779# a_7815_2035# 0.00386f
C3487 a_7701_2145# VGND 0.00231f
C3488 a_9419_2143# sky130_fd_sc_hd__inv_1_0.A 0
C3489 a_4635_13809# a_4505_13107# 0.00115f
C3490 a_15672_4951# A 0
C3491 a_9597_13793# w_9402_14723# 0
C3492 a_9811_11277# w_9404_11491# 0.02399f
C3493 a_14975_1765# VPWR 0.00115f
C3494 a_15071_2131# VPWR 0
C3495 w_11078_4508# sky130_fd_sc_hd__inv_1_0.A 0
C3496 a_6362_2149# w_5454_1698# 0.00139f
C3497 a_10813_13753# VPWR 0.3558f
C3498 a_3820_5021# w_3668_4962# 0.05213f
C3499 a_5735_2149# a_5554_1783# 0
C3500 w_10674_14933# a_8113_13753# 0
C3501 a_2289_5307# VGND 1.20002f
C3502 a_15113_5459# a_15281_5459# 0
C3503 a_7635_5039# A 0
C3504 sky130_fd_sc_hd__mux2_1_0.A1 A 0.01978f
C3505 a_9867_12097# a_9467_13091# 0
C3506 sky130_fd_sc_hd__inv_1_5.Y a_23511_14701# 0.09907f
C3507 a_4903_15345# a_7173_15235# 0
C3508 a_9683_1777# VPWR 0.17495f
C3509 a_6885_1783# VGND 0.67804f
C3510 a_24407_14651# a_24318_14385# 0
C3511 VGND w_11008_1688# 0.29328f
C3512 a_11455_4593# sky130_fd_sc_hd__inv_1_0.A 0
C3513 w_12866_5378# sky130_fd_sc_hd__mux2_1_0.S 0.00344f
C3514 a_9585_4963# VGND 0.00223f
C3515 a_9671_5727# a_9725_5837# 0.03622f
C3516 a_10116_4963# w_9208_4512# 0.00139f
C3517 a_9557_5837# VGND 0.00294f
C3518 a_4755_12857# a_4839_12857# 0.00208f
C3519 w_7354_4954# VGND 0.29951f
C3520 a_15141_4951# a_15309_4951# 0
C3521 a_2313_2157# sky130_fd_sc_hd__inv_1_0.Y 0.05199f
C3522 a_9875_13765# w_10748_13967# 0.00175f
C3523 sky130_fd_sc_hd__inv_1_5.Y A 0.00452f
C3524 a_24962_14701# VGND 0.18885f
C3525 a_17125_4938# VPWR 0.06504f
C3526 a_4839_12857# a_4763_14525# 0
C3527 a_12481_5467# A 0.00206f
C3528 a_5851_13769# a_6329_12927# 0
C3529 a_5999_2149# a_5873_1757# 0.04534f
C3530 a_11385_2139# sky130_fd_sc_hd__inv_1_0.A 0
C3531 a_4915_10549# a_9811_11277# 0
C3532 a_6029_5409# a_5861_5409# 0
C3533 a_11108_1773# VGND 0.08645f
C3534 sky130_fd_sc_hd__mux2_1_0.A1 sky130_fd_sc_hd__mux2_1_0.A0 0.39945f
C3535 a_13201_1769# a_12976_1743# 0.00487f
C3536 a_6087_14735# w_5712_14949# 0.02211f
C3537 a_11359_4593# VPWR 0.00133f
C3538 a_10088_5837# VPWR 0.01964f
C3539 a_14946_4905# a_14888_5433# 0.00485f
C3540 a_10569_1777# VPWR 1.05228f
C3541 a_15309_4951# sky130_fd_sc_hd__mux2_1_0.S 0
C3542 a_6129_12927# VGND 0.00291f
C3543 a_6911_15235# VPWR 0
C3544 a_4849_11293# a_4903_15345# 0.30844f
C3545 a_5999_2149# sky130_fd_sc_hd__inv_1_0.A 0
C3546 a_4903_15345# w_5786_13983# 0.07513f
C3547 a_4915_10549# a_7113_13395# 0.16058f
C3548 a_9589_12125# w_9404_11491# 0.00155f
C3549 a_9727_11527# a_9599_10561# 0
C3550 a_14916_4559# A 0
C3551 w_4432_13071# VPWR 0.16326f
C3552 VPWR a_15936_1765# 0
C3553 a_12509_4593# a_12320_4959# 0
C3554 sky130_fd_sc_hd__inv_1_0.Y w_1768_1706# 0.25031f
C3555 a_6696_1783# a_5945_2039# 0.00682f
C3556 a_11427_5833# VPWR 0
C3557 a_24774_14701# VGND 0.06373f
C3558 a_1920_1765# VGND 0.40886f
C3559 a_4576_5047# a_5903_5017# 0
C3560 VGND a_11824_13629# 0.13594f
C3561 a_6003_11935# a_5975_12927# 0
C3562 a_9809_14509# a_9725_14759# 0.07979f
C3563 a_15978_5459# A 0
C3564 a_4910_5047# VGND 0
C3565 w_12566_13951# VPWR 0.07508f
C3566 a_11824_13629# a_9799_16073# 0
C3567 a_11230_4567# VGND 0.38979f
C3568 a_7815_2035# a_8566_1779# 0.00682f
C3569 w_5484_4958# VGND 0.29342f
C3570 a_15141_4951# a_14946_4905# 0.00207f
C3571 a_9477_11527# w_9404_11491# 0.06993f
C3572 a_9865_15329# w_11532_15433# 0
C3573 a_5099_5047# a_4910_5413# 0
C3574 a_11178_4593# w_11078_4508# 0.01793f
C3575 a_11958_5467# a_11541_5723# 0.03016f
C3576 a_9629_2033# a_9515_2143# 0
C3577 a_9867_12097# VPWR 0.28921f
C3578 ua[0] sky130_fd_sc_hd__inv_1_0.A 0
C3579 ua[4] VGND 0
C3580 a_10116_4597# a_10639_4597# 0
C3581 a_3199_1791# w_1768_1706# 0.02026f
C3582 sky130_fd_sc_hd__inv_1_2.A w_12566_13951# 0.02092f
C3583 a_4129_2043# VGND 1.20051f
C3584 w_14694_1680# VPWR 0.50762f
C3585 a_13147_5463# a_13285_5437# 0
C3586 a_10813_13753# w_9500_13979# 0
C3587 a_2289_5307# a_3820_5021# 0.00446f
C3588 a_9875_13765# a_9683_13793# 0.00222f
C3589 a_15309_4585# a_14946_4905# 0.01182f
C3590 a_14794_1765# sky130_fd_sc_hd__inv_1_0.A 0.00159f
C3591 a_6087_14735# a_6389_13769# 0.00427f
C3592 a_14946_4905# a_15281_5459# 0.00242f
C3593 a_13018_5437# a_13411_5463# 0.02283f
C3594 a_9589_12125# a_4915_10549# 0.00128f
C3595 a_4513_14775# a_6087_14735# 0
C3596 a_4849_11293# a_4755_13107# 0
C3597 a_9308_4597# VPWR 0.10729f
C3598 a_14946_4905# sky130_fd_sc_hd__mux2_1_0.S 0.56407f
C3599 a_7815_2035# VPWR 0.34502f
C3600 a_15978_5459# sky130_fd_sc_hd__mux2_1_0.A0 0
C3601 a_14108_5463# VGND 0
C3602 a_23731_14309# a_24234_14385# 0.12294f
C3603 a_11623_4593# w_11078_4508# 0.01092f
C3604 a_6392_5043# VGND 0.01331f
C3605 w_7604_13967# a_7173_15235# 0.11864f
C3606 a_3738_1787# a_2259_2047# 0
C3607 a_2079_5051# VPWR 0.00123f
C3608 a_15281_5459# a_14888_5433# 0.02283f
C3609 a_10771_14747# a_9475_14759# 0
C3610 a_2313_1791# w_1768_1706# 0.01092f
C3611 a_9477_11527# a_4915_10549# 0.00232f
C3612 a_4159_5303# a_4045_5047# 0
C3613 a_6915_5043# a_6726_5409# 0
C3614 VGND w_12894_4504# 0.28722f
C3615 a_3768_5047# a_3229_5051# 0.0725f
C3616 a_10857_14747# VPWR 0
C3617 a_9585_4597# a_9360_4571# 0.00487f
C3618 a_6389_13769# a_7113_13395# 0.06159f
C3619 a_17339_4938# a_17125_4938# 0.00557f
C3620 a_11289_1773# VGND 0
C3621 a_9332_5445# a_9461_5471# 0.00758f
C3622 sky130_fd_sc_hd__inv_1_2.Y a_5809_14763# 0
C3623 a_11986_4959# VGND 0.18607f
C3624 a_14888_5433# sky130_fd_sc_hd__mux2_1_0.S 0
C3625 a_13313_4563# a_13018_5437# 0
C3626 a_4627_12141# a_4755_13107# 0
C3627 a_8113_13753# a_7113_13395# 0.02955f
C3628 a_14846_1739# VPWR 0.29469f
C3629 a_9290_1751# a_8755_1779# 0.11411f
C3630 a_1920_1765# a_2049_1791# 0.00758f
C3631 a_11623_4593# a_11455_4593# 0
C3632 a_10611_5471# a_13285_5437# 0
C3633 a_14136_4589# a_13385_4845# 0.00682f
C3634 a_11906_13629# a_12075_13379# 0
C3635 a_7476_1753# a_7605_2145# 0.00792f
C3636 VGND a_4625_15373# 0.24327f
C3637 a_13271_4955# VGND 0.00234f
C3638 a_5945_2039# VPWR 0.34533f
C3639 a_7506_5013# a_5975_5299# 0.00446f
C3640 a_9489_4963# VPWR 0
C3641 a_5831_1783# a_5945_2039# 0
C3642 a_6862_13645# a_6329_12927# 0.10646f
C3643 a_4213_5413# a_4045_5413# 0
C3644 a_4913_13781# a_6021_13769# 0.00104f
C3645 a_10965_11919# a_9875_13765# 0
C3646 a_5831_2149# a_5945_2039# 0
C3647 a_10813_13753# a_10895_13753# 0.00578f
C3648 a_4903_15345# w_4440_14739# 0.00599f
C3649 a_8596_5405# VPWR 0
C3650 a_12135_15219# a_11351_13753# 0.00152f
C3651 a_7869_1779# VGND 0.01554f
C3652 a_11289_2139# VPWR 0
C3653 a_9753_4597# VGND 0.01261f
C3654 a_10813_13753# a_11243_11891# 0
C3655 a_15113_5459# a_14297_5463# 0
C3656 w_12866_5378# a_14297_5463# 0.02026f
C3657 a_9290_1751# a_9419_1777# 0.00758f
C3658 a_4903_15345# a_4711_15373# 0.00101f
C3659 a_4915_10549# a_9683_13793# 0
C3660 a_6087_14735# a_4839_12857# 0.02474f
C3661 a_24234_14385# A 0.07599f
C3662 a_8113_13753# w_10748_13967# 0
C3663 a_11569_4849# a_12481_5467# 0
C3664 a_4837_16089# a_5851_13769# 0.08387f
C3665 a_9589_12125# w_9502_10747# 0
C3666 a_9489_4597# sky130_fd_sc_hd__inv_1_0.A 0
C3667 a_11986_4593# sky130_fd_sc_hd__inv_1_0.A 0
C3668 a_9685_10561# VPWR 0.00176f
C3669 A w_14736_5374# 0.00647f
C3670 a_9683_1777# a_9515_1777# 0
C3671 a_9465_16323# w_9490_15543# 0.0035f
C3672 a_10639_4597# A 0
C3673 a_5584_5043# a_5765_5409# 0
C3674 a_7506_5013# a_7899_5405# 0.02301f
C3675 a_7669_14003# VGND 0.24155f
C3676 w_4430_16303# VGND 0.06271f
C3677 VGND a_11089_13753# 0.00413f
C3678 a_11089_13753# a_9799_16073# 0.00702f
C3679 a_10813_13753# a_10983_13753# 0.00167f
C3680 a_9699_4853# sky130_fd_sc_hd__inv_1_0.A 0
C3681 a_15672_4951# w_14764_4500# 0.00139f
C3682 a_9675_12125# a_4915_10549# 0
C3683 a_7605_1779# a_6885_1783# 0
C3684 a_7845_5295# a_9308_4597# 0
C3685 VGND a_9467_13091# 0.29689f
C3686 a_9477_11527# w_9502_10747# 0.0035f
C3687 a_9465_16323# w_9402_14723# 0
C3688 a_7113_13395# a_4839_12857# 0.00444f
C3689 a_4880_1787# VGND 0
C3690 a_24152_14385# VGND 0.22746f
C3691 a_6029_5409# a_5903_5017# 0.04534f
C3692 a_4839_12857# a_4587_13107# 0
C3693 a_13357_5719# w_14736_5374# 0
C3694 VGND w_4538_13995# 0.11975f
C3695 sky130_fd_sc_hd__mux2_1_0.A1 w_14764_4500# 0.02202f
C3696 a_15309_4951# a_14297_5463# 0
C3697 a_9809_14509# a_11351_13753# 0
C3698 a_14864_4585# a_14916_4559# 0.1439f
C3699 a_3790_1761# VGND 0.40141f
C3700 a_6696_1783# VGND 0
C3701 a_2175_5051# VGND 0
C3702 ua[1] VNB 0.14696f
C3703 ua[2] VNB 0.14696f
C3704 ua[3] VNB 0.14696f
C3705 ua[4] VNB 0.14465f
C3706 ua[5] VNB 0.14471f
C3707 ua[6] VNB 0.14538f
C3708 ua[7] VNB 0.1455f
C3709 ena VNB 0.07038f
C3710 clk VNB 0.04288f
C3711 rst_n VNB 0.04288f
C3712 ui_in[2] VNB 0.04288f
C3713 ui_in[3] VNB 0.04288f
C3714 ui_in[4] VNB 0.04288f
C3715 ui_in[5] VNB 0.04288f
C3716 ui_in[6] VNB 0.04288f
C3717 ui_in[7] VNB 0.04288f
C3718 uio_in[0] VNB 0.04288f
C3719 uio_in[1] VNB 0.04288f
C3720 uio_in[2] VNB 0.04288f
C3721 uio_in[3] VNB 0.04288f
C3722 uio_in[4] VNB 0.04288f
C3723 uio_in[5] VNB 0.04288f
C3724 uio_in[6] VNB 0.04288f
C3725 uio_in[7] VNB 0.04288f
C3726 uo_out[0] VNB 0.04288f
C3727 uo_out[1] VNB 0.04288f
C3728 uo_out[2] VNB 0.04288f
C3729 uo_out[3] VNB 0.04288f
C3730 uo_out[4] VNB 0.04288f
C3731 uo_out[5] VNB 0.04288f
C3732 uo_out[6] VNB 0.04288f
C3733 uo_out[7] VNB 0.04288f
C3734 uio_out[0] VNB 0.04288f
C3735 uio_out[1] VNB 0.04288f
C3736 uio_out[2] VNB 0.04288f
C3737 uio_out[3] VNB 0.04288f
C3738 uio_out[4] VNB 0.04288f
C3739 uio_out[5] VNB 0.04288f
C3740 uio_out[6] VNB 0.04288f
C3741 uio_out[7] VNB 0.04288f
C3742 uio_oe[0] VNB 0.04288f
C3743 uio_oe[1] VNB 0.04288f
C3744 uio_oe[2] VNB 0.04288f
C3745 uio_oe[3] VNB 0.04288f
C3746 uio_oe[4] VNB 0.04288f
C3747 uio_oe[5] VNB 0.04288f
C3748 uio_oe[6] VNB 0.04288f
C3749 uio_oe[7] VNB 0.07038f
C3750 Y VNB 2.29089f
C3751 ua[0] VNB 9.60658f
C3752 A VNB 10.0952f
C3753 ui_in[0] VNB 8.89585f
C3754 ui_in[1] VNB 8.7197f
C3755 VPWR VNB 79.9919f
C3756 VGND VNB 90.63161f
C3757 VPB VNB 0.33898f
C3758 a_15602_1765# VNB 0.00345f
C3759 a_15239_1765# VNB 0.00484f
C3760 a_13732_1769# VNB 0.00345f
C3761 a_13369_1769# VNB 0.00484f
C3762 a_15602_2131# VNB 0.01578f
C3763 a_15239_2131# VNB 0.01584f
C3764 a_14794_1765# VNB 0.06682f
C3765 a_15185_2021# VNB 0.27343f
C3766 a_14846_1739# VNB 0.13081f
C3767 a_14255_1769# VNB 0.55211f
C3768 a_11916_1773# VNB 0.00345f
C3769 a_11553_1773# VNB 0.00484f
C3770 a_13732_2135# VNB 0.01578f
C3771 a_13369_2135# VNB 0.01584f
C3772 a_12924_1769# VNB 0.06298f
C3773 a_13315_2025# VNB 0.26543f
C3774 a_13243_1743# VNB 0.46761f
C3775 a_12976_1743# VNB 0.13025f
C3776 a_12439_1773# VNB 0.05657f
C3777 a_10046_1777# VNB 0.00345f
C3778 a_9683_1777# VNB 0.00484f
C3779 a_11916_2139# VNB 0.01578f
C3780 a_11553_2139# VNB 0.01584f
C3781 a_11108_1773# VNB 0.06682f
C3782 a_11499_2029# VNB 0.26466f
C3783 a_11160_1747# VNB 0.13081f
C3784 a_10569_1777# VNB 0.55211f
C3785 a_8232_1779# VNB 0.00345f
C3786 a_7869_1779# VNB 0.00484f
C3787 a_10046_2143# VNB 0.01578f
C3788 a_9683_2143# VNB 0.01584f
C3789 a_9238_1777# VNB 0.06285f
C3790 a_9629_2033# VNB 0.26543f
C3791 a_9290_1751# VNB 0.13016f
C3792 a_8755_1779# VNB 0.52093f
C3793 a_6362_1783# VNB 0.00345f
C3794 a_5999_1783# VNB 0.00484f
C3795 a_8232_2145# VNB 0.01578f
C3796 a_7869_2145# VNB 0.01584f
C3797 a_7424_1779# VNB 0.06682f
C3798 a_7815_2035# VNB 0.26452f
C3799 a_7476_1753# VNB 0.13081f
C3800 a_6885_1783# VNB 0.55211f
C3801 a_4546_1787# VNB 0.00345f
C3802 a_4183_1787# VNB 0.00484f
C3803 a_6362_2149# VNB 0.01578f
C3804 a_5999_2149# VNB 0.01584f
C3805 a_5554_1783# VNB 0.06298f
C3806 a_5945_2039# VNB 0.26543f
C3807 a_5873_1757# VNB 0.46708f
C3808 a_5606_1757# VNB 0.13025f
C3809 a_5069_1787# VNB 0.05657f
C3810 a_2676_1791# VNB 0.00345f
C3811 a_2313_1791# VNB 0.00484f
C3812 a_4546_2153# VNB 0.01578f
C3813 a_4183_2153# VNB 0.01584f
C3814 a_3738_1787# VNB 0.06682f
C3815 a_4129_2043# VNB 0.26466f
C3816 a_3790_1761# VNB 0.13081f
C3817 a_3199_1791# VNB 0.55211f
C3818 a_2676_2157# VNB 0.01578f
C3819 a_2313_2157# VNB 0.01584f
C3820 a_1868_1791# VNB 0.10031f
C3821 a_2259_2047# VNB 0.26543f
C3822 a_1920_1765# VNB 0.1359f
C3823 sky130_fd_sc_hd__inv_1_0.Y VNB 2.28963f
C3824 a_15672_4585# VNB 0.00345f
C3825 a_15309_4585# VNB 0.00484f
C3826 a_13802_4589# VNB 0.00345f
C3827 a_13439_4589# VNB 0.00484f
C3828 a_15672_4951# VNB 0.01578f
C3829 a_15309_4951# VNB 0.01584f
C3830 a_14864_4585# VNB 0.06682f
C3831 a_15255_4841# VNB 0.26397f
C3832 a_14946_4905# VNB 1.04897f
C3833 a_14916_4559# VNB 0.12906f
C3834 a_14325_4589# VNB 0.51247f
C3835 a_11986_4593# VNB 0.00345f
C3836 a_11623_4593# VNB 0.00484f
C3837 a_13802_4955# VNB 0.01578f
C3838 a_13439_4955# VNB 0.01584f
C3839 a_12994_4589# VNB 0.06298f
C3840 a_13385_4845# VNB 0.26214f
C3841 a_13313_4563# VNB 0.43239f
C3842 a_13046_4563# VNB 0.12849f
C3843 a_12509_4593# VNB 0.05657f
C3844 a_10116_4597# VNB 0.00345f
C3845 a_9753_4597# VNB 0.00484f
C3846 a_11986_4959# VNB 0.01578f
C3847 a_11623_4959# VNB 0.01584f
C3848 a_11178_4593# VNB 0.06682f
C3849 a_11569_4849# VNB 0.26136f
C3850 a_11230_4567# VNB 0.12906f
C3851 a_10639_4597# VNB 0.51206f
C3852 a_10116_4963# VNB 0.01578f
C3853 a_9753_4963# VNB 0.01584f
C3854 a_9308_4597# VNB 0.09346f
C3855 a_9699_4853# VNB 0.26214f
C3856 a_9360_4571# VNB 0.13349f
C3857 a_8262_5039# VNB 0.00345f
C3858 a_7899_5039# VNB 0.00484f
C3859 a_17125_4938# VNB 0.13914f
C3860 sky130_fd_sc_hd__mux2_1_0.A1 VNB 0.44799f
C3861 a_16871_4938# VNB 0.23758f
C3862 a_15644_5459# VNB 0.00345f
C3863 a_15281_5459# VNB 0.00484f
C3864 sky130_fd_sc_hd__mux2_1_0.A0 VNB 0.5186f
C3865 a_13774_5463# VNB 0.00345f
C3866 a_13411_5463# VNB 0.00484f
C3867 a_15644_5825# VNB 0.01578f
C3868 a_15281_5825# VNB 0.01584f
C3869 a_14836_5459# VNB 0.06682f
C3870 a_15227_5715# VNB 0.27134f
C3871 a_14888_5433# VNB 0.12984f
C3872 a_14297_5463# VNB 0.50345f
C3873 a_11958_5467# VNB 0.00345f
C3874 a_11595_5467# VNB 0.00484f
C3875 a_13774_5829# VNB 0.01578f
C3876 a_13411_5829# VNB 0.01584f
C3877 a_12966_5463# VNB 0.06298f
C3878 a_13357_5719# VNB 0.26335f
C3879 a_13285_5437# VNB 0.42555f
C3880 a_13018_5437# VNB 0.12928f
C3881 a_12481_5467# VNB 0.05657f
C3882 a_10088_5471# VNB 0.00345f
C3883 a_9725_5471# VNB 0.00484f
C3884 a_11958_5833# VNB 0.01578f
C3885 a_11595_5833# VNB 0.01584f
C3886 a_11150_5467# VNB 0.06682f
C3887 a_11541_5723# VNB 0.26257f
C3888 a_11202_5441# VNB 0.12984f
C3889 a_10611_5471# VNB 0.50409f
C3890 sky130_fd_sc_hd__mux2_1_0.S VNB 1.40108f
C3891 a_6392_5043# VNB 0.00345f
C3892 a_6029_5043# VNB 0.00484f
C3893 a_8262_5405# VNB 0.01578f
C3894 a_7899_5405# VNB 0.01584f
C3895 a_7454_5039# VNB 0.06682f
C3896 a_7845_5295# VNB 0.27171f
C3897 a_7506_5013# VNB 0.13081f
C3898 a_6915_5043# VNB 0.55211f
C3899 a_4576_5047# VNB 0.00345f
C3900 a_4213_5047# VNB 0.00484f
C3901 a_6392_5409# VNB 0.01578f
C3902 a_6029_5409# VNB 0.01584f
C3903 a_5584_5043# VNB 0.06298f
C3904 a_5975_5299# VNB 0.26543f
C3905 a_5903_5017# VNB 0.46708f
C3906 a_5636_5017# VNB 0.13025f
C3907 a_5099_5047# VNB 0.05657f
C3908 a_2706_5051# VNB 0.00345f
C3909 a_2343_5051# VNB 0.00484f
C3910 a_4576_5413# VNB 0.01578f
C3911 a_4213_5413# VNB 0.01584f
C3912 a_3768_5047# VNB 0.06682f
C3913 a_4159_5303# VNB 0.26466f
C3914 a_3820_5021# VNB 0.13081f
C3915 a_3229_5051# VNB 0.55211f
C3916 a_2706_5417# VNB 0.01578f
C3917 a_2343_5417# VNB 0.01584f
C3918 a_1898_5051# VNB 0.10031f
C3919 a_2289_5307# VNB 0.26543f
C3920 a_1950_5025# VNB 0.1359f
C3921 a_10088_5837# VNB 0.01578f
C3922 a_9725_5837# VNB 0.01584f
C3923 a_9280_5471# VNB 0.09442f
C3924 a_9671_5727# VNB 0.26335f
C3925 a_9332_5445# VNB 0.13493f
C3926 a_9599_10561# VNB 0.1752f
C3927 a_4637_10577# VNB 0.1752f
C3928 a_9727_11527# VNB 0.00137f
C3929 a_9477_11527# VNB 0.24712f
C3930 a_4765_11543# VNB 0.00137f
C3931 a_4515_11543# VNB 0.24712f
C3932 a_10965_11919# VNB 0.1732f
C3933 a_9867_12097# VNB 0.54635f
C3934 a_6003_11935# VNB 0.1732f
C3935 a_9589_12125# VNB 0.17114f
C3936 a_4905_12113# VNB 0.55094f
C3937 a_4627_12141# VNB 0.17114f
C3938 a_9717_13091# VNB 0.00137f
C3939 a_9467_13091# VNB 0.24424f
C3940 a_10937_12911# VNB 0.16539f
C3941 a_4755_13107# VNB 0.00137f
C3942 a_4505_13107# VNB 0.24424f
C3943 a_5975_12927# VNB 0.16539f
C3944 a_11291_12911# VNB 0.46058f
C3945 a_11824_13629# VNB 0.1516f
C3946 a_12075_13379# VNB 0.40216f
C3947 a_11243_11891# VNB 1.12822f
C3948 a_9877_10533# VNB 3.44942f
C3949 a_12631_13987# VNB 0.15779f
C3950 a_11351_13753# VNB 0.31965f
C3951 a_10813_13753# VNB 0.16387f
C3952 a_9875_13765# VNB 0.45251f
C3953 a_6329_12927# VNB 0.46058f
C3954 a_6862_13645# VNB 0.1516f
C3955 a_7113_13395# VNB 0.39872f
C3956 a_6281_11907# VNB 1.1397f
C3957 a_4915_10549# VNB 3.27518f
C3958 a_9597_13793# VNB 0.16601f
C3959 a_7669_14003# VNB 0.1564f
C3960 a_6389_13769# VNB 0.31965f
C3961 a_5851_13769# VNB 0.16387f
C3962 a_4913_13781# VNB 0.45689f
C3963 a_4635_13809# VNB 0.17003f
C3964 a_24318_14385# VNB 0.02499f
C3965 a_24152_14385# VNB 0.02039f
C3966 a_23511_14335# VNB 0.04207f
C3967 a_24962_14701# VNB 0.16413f
C3968 a_24774_14701# VNB 0.2179f
C3969 a_24234_14385# VNB 0.03874f
C3970 a_24241_14651# VNB 0.00666f
C3971 sky130_fd_sc_hd__inv_1_0.A VNB 11.8725f
C3972 a_23731_14309# VNB 0.33779f
C3973 a_23677_14701# VNB 0.00373f
C3974 a_23511_14701# VNB 0.02865f
C3975 a_9725_14759# VNB 0.00137f
C3976 a_9475_14759# VNB 0.24496f
C3977 a_9801_12841# VNB 1.33033f
C3978 a_9811_11277# VNB 2.17869f
C3979 a_10771_14747# VNB 0.1671f
C3980 a_4763_14775# VNB 0.00137f
C3981 a_4513_14775# VNB 0.24496f
C3982 a_4839_12857# VNB 1.33478f
C3983 a_4849_11293# VNB 2.17869f
C3984 a_5809_14763# VNB 0.1671f
C3985 a_12135_15219# VNB 0.75127f
C3986 a_11597_15219# VNB 0.17279f
C3987 a_11049_14719# VNB 0.33714f
C3988 a_9809_14509# VNB 0.62284f
C3989 a_8113_13753# VNB 3.07869f
C3990 a_9865_15329# VNB 0.69482f
C3991 a_7173_15235# VNB 0.79677f
C3992 a_6635_15235# VNB 0.17279f
C3993 a_6087_14735# VNB 0.33714f
C3994 a_4847_14525# VNB 0.63122f
C3995 a_9587_15357# VNB 0.17275f
C3996 a_4903_15345# VNB 0.69937f
C3997 a_4625_15373# VNB 0.17275f
C3998 sky130_fd_sc_hd__inv_1_5.A VNB 0.45825f
C3999 sky130_fd_sc_hd__inv_1_4.A VNB 0.40476f
C4000 a_9799_16073# VNB 1.62449f
C4001 a_9715_16323# VNB 0.00137f
C4002 a_9465_16323# VNB 0.24845f
C4003 a_4837_16089# VNB 1.72323f
C4004 a_4753_16339# VNB 0.00137f
C4005 a_4503_16339# VNB 0.24845f
C4006 sky130_fd_sc_hd__inv_1_5.Y VNB 4.18678f
C4007 sky130_fd_sc_hd__inv_1_2.Y VNB 2.47775f
C4008 sky130_fd_sc_hd__inv_1_2.A VNB 8.34761f
C4009 w_14694_1680# VNB 1.49072f
C4010 w_12824_1684# VNB 1.49072f
C4011 w_11008_1688# VNB 1.49072f
C4012 w_9138_1692# VNB 1.49072f
C4013 w_7324_1694# VNB 1.49072f
C4014 w_5454_1698# VNB 1.49072f
C4015 w_3638_1702# VNB 1.49072f
C4016 w_1768_1706# VNB 1.49072f
C4017 sky130_fd_sc_hd__inv_1_0.VPB VNB 0.33898f
C4018 sky130_fd_sc_hd__mux2_1_0.VPB VNB 0.87055f
C4019 w_14764_4500# VNB 1.49072f
C4020 w_12894_4504# VNB 1.49072f
C4021 w_11078_4508# VNB 1.49072f
C4022 w_9208_4512# VNB 1.49072f
C4023 w_7354_4954# VNB 1.49072f
C4024 w_5484_4958# VNB 1.49072f
C4025 w_3668_4962# VNB 1.49072f
C4026 w_1798_4966# VNB 1.49072f
C4027 w_14736_5374# VNB 1.49072f
C4028 w_12866_5378# VNB 1.49072f
C4029 w_11050_5382# VNB 1.49072f
C4030 w_9180_5386# VNB 1.49072f
C4031 w_9502_10747# VNB 0.51617f
C4032 w_4540_10763# VNB 0.51617f
C4033 w_9404_11491# VNB 0.69336f
C4034 w_4442_11507# VNB 0.69336f
C4035 w_10868_12105# VNB 0.51617f
C4036 w_9492_12311# VNB 0.51617f
C4037 w_5906_12121# VNB 0.51617f
C4038 w_4530_12327# VNB 0.51617f
C4039 w_10872_13125# VNB 0.51617f
C4040 w_9394_13055# VNB 0.69336f
C4041 w_5910_13141# VNB 0.51617f
C4042 w_4432_13071# VNB 0.69336f
C4043 w_11718_13593# VNB 0.51617f
C4044 w_6756_13609# VNB 0.51617f
C4045 w_12566_13951# VNB 0.60476f
C4046 w_10748_13967# VNB 0.69336f
C4047 w_9500_13979# VNB 0.51617f
C4048 w_7604_13967# VNB 0.60476f
C4049 w_5786_13983# VNB 0.69336f
C4050 w_4538_13995# VNB 0.51617f
C4051 sky130_fd_sc_hd__mux4_1_0.VPB VNB 1.9337f
C4052 w_10674_14933# VNB 0.51617f
C4053 w_9402_14723# VNB 0.69336f
C4054 w_5712_14949# VNB 0.51617f
C4055 w_4440_14739# VNB 0.69336f
C4056 w_11532_15433# VNB 0.69336f
C4057 w_9490_15543# VNB 0.51617f
C4058 w_6570_15449# VNB 0.69336f
C4059 w_4528_15559# VNB 0.51617f
C4060 sky130_fd_sc_hd__inv_1_5.VPB VNB 0.33898f
C4061 sky130_fd_sc_hd__inv_1_4.VPB VNB 0.33898f
C4062 sky130_fd_sc_hd__inv_1_3.VPB VNB 0.33898f
C4063 w_9392_16287# VNB 0.69336f
C4064 w_4430_16303# VNB 0.69336f
C4065 sky130_fd_sc_hd__inv_1_2.VPB VNB 0.33898f
.ends

