magic
tech sky130A
magscale 1 2
timestamp 1754940301
<< error_s >>
rect -138 1011 582 1332
rect -65 797 -13 927
rect 17 797 71 927
rect 101 797 155 927
rect 185 797 239 927
rect 269 797 423 927
rect 453 797 517 927
rect -40 267 496 588
rect 253 165 305 183
rect 57 81 113 165
rect 143 81 197 165
rect 227 81 305 165
rect 253 53 305 81
rect 335 53 391 183
rect 2002 157 2722 478
rect 2482 27 2575 73
rect -128 -553 592 -232
rect 1144 -343 1680 -22
rect 2067 -57 2119 27
rect 2149 -57 2207 27
rect 2237 -57 2313 27
rect 2343 -57 2409 27
rect 2439 -57 2575 27
rect 2605 -57 2657 73
rect 1437 -445 1489 -427
rect 1241 -529 1297 -445
rect 1327 -529 1381 -445
rect 1411 -529 1489 -445
rect 1437 -557 1489 -529
rect 1519 -557 1575 -427
rect -55 -767 -3 -637
rect 27 -767 81 -637
rect 111 -767 165 -637
rect 195 -767 249 -637
rect 279 -767 433 -637
rect 463 -767 527 -637
rect -30 -1297 506 -976
rect 1218 -1309 1938 -988
rect 3116 -1325 3744 -1004
rect 263 -1399 315 -1381
rect 67 -1483 123 -1399
rect 153 -1483 207 -1399
rect 237 -1483 315 -1399
rect 263 -1511 315 -1483
rect 345 -1511 401 -1381
rect 1698 -1439 1791 -1393
rect 1283 -1523 1335 -1439
rect 1365 -1523 1423 -1439
rect 1453 -1523 1529 -1439
rect 1559 -1523 1625 -1439
rect 1655 -1523 1791 -1439
rect 1821 -1523 1873 -1393
rect 2188 -1683 2724 -1362
rect 3542 -1449 3595 -1409
rect 3181 -1533 3233 -1449
rect 3263 -1533 3329 -1449
rect 3359 -1533 3413 -1449
rect 3443 -1533 3497 -1449
rect 3527 -1533 3595 -1449
rect 3542 -1539 3595 -1533
rect 3625 -1539 3679 -1409
rect 2463 -1813 2515 -1767
rect -136 -2221 584 -1900
rect 1342 -2151 1878 -1830
rect 2282 -1897 2334 -1813
rect 2364 -1897 2418 -1813
rect 2448 -1897 2515 -1813
rect 2545 -1897 2597 -1767
rect 1681 -2281 1731 -2235
rect -63 -2435 -11 -2305
rect 19 -2435 73 -2305
rect 103 -2435 157 -2305
rect 187 -2435 241 -2305
rect 271 -2435 425 -2305
rect 455 -2435 519 -2305
rect 1407 -2365 1459 -2281
rect 1489 -2365 1531 -2281
rect 1561 -2365 1603 -2281
rect 1633 -2365 1731 -2281
rect 1761 -2365 1813 -2235
rect -38 -2965 498 -2644
rect 255 -3067 307 -3049
rect 59 -3151 115 -3067
rect 145 -3151 199 -3067
rect 229 -3151 307 -3067
rect 255 -3179 307 -3151
rect 337 -3179 393 -3049
rect 1338 -3171 1874 -2850
rect 1631 -3273 1683 -3255
rect 1435 -3357 1491 -3273
rect 1521 -3357 1575 -3273
rect 1605 -3357 1683 -3273
rect 1631 -3385 1683 -3357
rect 1713 -3385 1769 -3255
rect -126 -3785 594 -3464
rect -53 -3999 -1 -3869
rect 29 -3999 83 -3869
rect 113 -3999 167 -3869
rect 197 -3999 251 -3869
rect 281 -3999 435 -3869
rect 465 -3999 529 -3869
rect -28 -4529 508 -4208
rect 265 -4631 317 -4613
rect 69 -4715 125 -4631
rect 155 -4715 209 -4631
rect 239 -4715 317 -4631
rect 265 -4743 317 -4715
rect 347 -4743 403 -4613
<< nwell >>
rect -128 -553 592 -232
rect -30 -1297 506 -976
rect -136 -2221 584 -1900
rect -38 -2965 498 -2644
rect -126 -3785 594 -3464
rect -28 -4529 508 -4208
<< pwell >>
rect -81 -793 553 -611
rect -61 -831 -27 -793
rect 237 -1373 427 -1355
rect 41 -1537 427 -1373
rect 41 -1541 71 -1537
rect 37 -1575 71 -1541
rect -89 -2461 545 -2279
rect -69 -2499 -35 -2461
rect 229 -3041 419 -3023
rect 33 -3205 419 -3041
rect 33 -3209 63 -3205
rect 29 -3243 63 -3209
rect -79 -4025 555 -3843
rect -59 -4063 -25 -4025
rect 239 -4605 429 -4587
rect 43 -4769 429 -4605
rect 43 -4773 73 -4769
rect 39 -4807 73 -4773
<< ndiff >>
rect -55 -719 -3 -637
rect -55 -753 -47 -719
rect -13 -753 -3 -719
rect -55 -767 -3 -753
rect 27 -697 81 -637
rect 27 -731 37 -697
rect 71 -731 81 -697
rect 27 -767 81 -731
rect 111 -719 165 -637
rect 111 -753 121 -719
rect 155 -753 165 -719
rect 111 -767 165 -753
rect 195 -767 249 -637
rect 279 -717 433 -637
rect 279 -751 289 -717
rect 323 -751 389 -717
rect 423 -751 433 -717
rect 279 -767 433 -751
rect 463 -646 527 -637
rect 463 -680 479 -646
rect 513 -680 527 -646
rect 463 -714 527 -680
rect 463 -748 479 -714
rect 513 -748 527 -714
rect 463 -767 527 -748
rect 263 -1399 315 -1381
rect 67 -1437 123 -1399
rect 67 -1471 79 -1437
rect 113 -1471 123 -1437
rect 67 -1483 123 -1471
rect 153 -1483 207 -1399
rect 237 -1465 315 -1399
rect 237 -1483 271 -1465
rect 263 -1499 271 -1483
rect 305 -1499 315 -1465
rect 263 -1511 315 -1499
rect 345 -1465 401 -1381
rect 345 -1499 355 -1465
rect 389 -1499 401 -1465
rect 345 -1511 401 -1499
rect -63 -2387 -11 -2305
rect -63 -2421 -55 -2387
rect -21 -2421 -11 -2387
rect -63 -2435 -11 -2421
rect 19 -2365 73 -2305
rect 19 -2399 29 -2365
rect 63 -2399 73 -2365
rect 19 -2435 73 -2399
rect 103 -2387 157 -2305
rect 103 -2421 113 -2387
rect 147 -2421 157 -2387
rect 103 -2435 157 -2421
rect 187 -2435 241 -2305
rect 271 -2385 425 -2305
rect 271 -2419 281 -2385
rect 315 -2419 381 -2385
rect 415 -2419 425 -2385
rect 271 -2435 425 -2419
rect 455 -2314 519 -2305
rect 455 -2348 471 -2314
rect 505 -2348 519 -2314
rect 455 -2382 519 -2348
rect 455 -2416 471 -2382
rect 505 -2416 519 -2382
rect 455 -2435 519 -2416
rect 255 -3067 307 -3049
rect 59 -3105 115 -3067
rect 59 -3139 71 -3105
rect 105 -3139 115 -3105
rect 59 -3151 115 -3139
rect 145 -3151 199 -3067
rect 229 -3133 307 -3067
rect 229 -3151 263 -3133
rect 255 -3167 263 -3151
rect 297 -3167 307 -3133
rect 255 -3179 307 -3167
rect 337 -3133 393 -3049
rect 337 -3167 347 -3133
rect 381 -3167 393 -3133
rect 337 -3179 393 -3167
rect -53 -3951 -1 -3869
rect -53 -3985 -45 -3951
rect -11 -3985 -1 -3951
rect -53 -3999 -1 -3985
rect 29 -3929 83 -3869
rect 29 -3963 39 -3929
rect 73 -3963 83 -3929
rect 29 -3999 83 -3963
rect 113 -3951 167 -3869
rect 113 -3985 123 -3951
rect 157 -3985 167 -3951
rect 113 -3999 167 -3985
rect 197 -3999 251 -3869
rect 281 -3949 435 -3869
rect 281 -3983 291 -3949
rect 325 -3983 391 -3949
rect 425 -3983 435 -3949
rect 281 -3999 435 -3983
rect 465 -3878 529 -3869
rect 465 -3912 481 -3878
rect 515 -3912 529 -3878
rect 465 -3946 529 -3912
rect 465 -3980 481 -3946
rect 515 -3980 529 -3946
rect 465 -3999 529 -3980
rect 265 -4631 317 -4613
rect 69 -4669 125 -4631
rect 69 -4703 81 -4669
rect 115 -4703 125 -4669
rect 69 -4715 125 -4703
rect 155 -4715 209 -4631
rect 239 -4697 317 -4631
rect 239 -4715 273 -4697
rect 265 -4731 273 -4715
rect 307 -4731 317 -4697
rect 265 -4743 317 -4731
rect 347 -4697 403 -4613
rect 347 -4731 357 -4697
rect 391 -4731 403 -4697
rect 347 -4743 403 -4731
<< pdiff >>
rect -55 -329 -3 -317
rect -55 -363 -47 -329
rect -13 -363 -3 -329
rect -55 -397 -3 -363
rect -55 -431 -47 -397
rect -13 -431 -3 -397
rect -55 -517 -3 -431
rect 27 -517 81 -317
rect 111 -339 165 -317
rect 111 -373 121 -339
rect 155 -373 165 -339
rect 111 -407 165 -373
rect 111 -441 121 -407
rect 155 -441 165 -407
rect 111 -517 165 -441
rect 195 -339 249 -317
rect 195 -373 205 -339
rect 239 -373 249 -339
rect 195 -407 249 -373
rect 195 -441 205 -407
rect 239 -441 249 -407
rect 195 -517 249 -441
rect 279 -339 331 -317
rect 279 -373 289 -339
rect 323 -373 331 -339
rect 279 -517 331 -373
rect 385 -339 437 -317
rect 385 -373 393 -339
rect 427 -373 437 -339
rect 385 -407 437 -373
rect 385 -441 393 -407
rect 427 -441 437 -407
rect 385 -517 437 -441
rect 467 -337 527 -317
rect 467 -371 477 -337
rect 511 -371 527 -337
rect 467 -405 527 -371
rect 467 -439 477 -405
rect 511 -439 527 -405
rect 467 -473 527 -439
rect 467 -507 477 -473
rect 511 -507 527 -473
rect 467 -517 527 -507
rect 263 -1073 315 -1061
rect 263 -1103 271 -1073
rect 67 -1115 123 -1103
rect 67 -1149 79 -1115
rect 113 -1149 123 -1115
rect 67 -1187 123 -1149
rect 153 -1115 207 -1103
rect 153 -1149 163 -1115
rect 197 -1149 207 -1115
rect 153 -1187 207 -1149
rect 237 -1107 271 -1103
rect 305 -1107 315 -1073
rect 237 -1141 315 -1107
rect 237 -1175 271 -1141
rect 305 -1175 315 -1141
rect 237 -1187 315 -1175
rect 253 -1261 315 -1187
rect 345 -1073 440 -1061
rect 345 -1107 375 -1073
rect 409 -1107 440 -1073
rect 345 -1141 440 -1107
rect 345 -1175 375 -1141
rect 409 -1175 440 -1141
rect 345 -1261 440 -1175
rect -63 -1997 -11 -1985
rect -63 -2031 -55 -1997
rect -21 -2031 -11 -1997
rect -63 -2065 -11 -2031
rect -63 -2099 -55 -2065
rect -21 -2099 -11 -2065
rect -63 -2185 -11 -2099
rect 19 -2185 73 -1985
rect 103 -2007 157 -1985
rect 103 -2041 113 -2007
rect 147 -2041 157 -2007
rect 103 -2075 157 -2041
rect 103 -2109 113 -2075
rect 147 -2109 157 -2075
rect 103 -2185 157 -2109
rect 187 -2007 241 -1985
rect 187 -2041 197 -2007
rect 231 -2041 241 -2007
rect 187 -2075 241 -2041
rect 187 -2109 197 -2075
rect 231 -2109 241 -2075
rect 187 -2185 241 -2109
rect 271 -2007 323 -1985
rect 271 -2041 281 -2007
rect 315 -2041 323 -2007
rect 271 -2185 323 -2041
rect 377 -2007 429 -1985
rect 377 -2041 385 -2007
rect 419 -2041 429 -2007
rect 377 -2075 429 -2041
rect 377 -2109 385 -2075
rect 419 -2109 429 -2075
rect 377 -2185 429 -2109
rect 459 -2005 519 -1985
rect 459 -2039 469 -2005
rect 503 -2039 519 -2005
rect 459 -2073 519 -2039
rect 459 -2107 469 -2073
rect 503 -2107 519 -2073
rect 459 -2141 519 -2107
rect 459 -2175 469 -2141
rect 503 -2175 519 -2141
rect 459 -2185 519 -2175
rect 255 -2741 307 -2729
rect 255 -2771 263 -2741
rect 59 -2783 115 -2771
rect 59 -2817 71 -2783
rect 105 -2817 115 -2783
rect 59 -2855 115 -2817
rect 145 -2783 199 -2771
rect 145 -2817 155 -2783
rect 189 -2817 199 -2783
rect 145 -2855 199 -2817
rect 229 -2775 263 -2771
rect 297 -2775 307 -2741
rect 229 -2809 307 -2775
rect 229 -2843 263 -2809
rect 297 -2843 307 -2809
rect 229 -2855 307 -2843
rect 245 -2929 307 -2855
rect 337 -2741 432 -2729
rect 337 -2775 367 -2741
rect 401 -2775 432 -2741
rect 337 -2809 432 -2775
rect 337 -2843 367 -2809
rect 401 -2843 432 -2809
rect 337 -2929 432 -2843
rect -53 -3561 -1 -3549
rect -53 -3595 -45 -3561
rect -11 -3595 -1 -3561
rect -53 -3629 -1 -3595
rect -53 -3663 -45 -3629
rect -11 -3663 -1 -3629
rect -53 -3749 -1 -3663
rect 29 -3749 83 -3549
rect 113 -3571 167 -3549
rect 113 -3605 123 -3571
rect 157 -3605 167 -3571
rect 113 -3639 167 -3605
rect 113 -3673 123 -3639
rect 157 -3673 167 -3639
rect 113 -3749 167 -3673
rect 197 -3571 251 -3549
rect 197 -3605 207 -3571
rect 241 -3605 251 -3571
rect 197 -3639 251 -3605
rect 197 -3673 207 -3639
rect 241 -3673 251 -3639
rect 197 -3749 251 -3673
rect 281 -3571 333 -3549
rect 281 -3605 291 -3571
rect 325 -3605 333 -3571
rect 281 -3749 333 -3605
rect 387 -3571 439 -3549
rect 387 -3605 395 -3571
rect 429 -3605 439 -3571
rect 387 -3639 439 -3605
rect 387 -3673 395 -3639
rect 429 -3673 439 -3639
rect 387 -3749 439 -3673
rect 469 -3569 529 -3549
rect 469 -3603 479 -3569
rect 513 -3603 529 -3569
rect 469 -3637 529 -3603
rect 469 -3671 479 -3637
rect 513 -3671 529 -3637
rect 469 -3705 529 -3671
rect 469 -3739 479 -3705
rect 513 -3739 529 -3705
rect 469 -3749 529 -3739
rect 265 -4305 317 -4293
rect 265 -4335 273 -4305
rect 69 -4347 125 -4335
rect 69 -4381 81 -4347
rect 115 -4381 125 -4347
rect 69 -4419 125 -4381
rect 155 -4347 209 -4335
rect 155 -4381 165 -4347
rect 199 -4381 209 -4347
rect 155 -4419 209 -4381
rect 239 -4339 273 -4335
rect 307 -4339 317 -4305
rect 239 -4373 317 -4339
rect 239 -4407 273 -4373
rect 307 -4407 317 -4373
rect 239 -4419 317 -4407
rect 255 -4493 317 -4419
rect 347 -4305 442 -4293
rect 347 -4339 377 -4305
rect 411 -4339 442 -4305
rect 347 -4373 442 -4339
rect 347 -4407 377 -4373
rect 411 -4407 442 -4373
rect 347 -4493 442 -4407
<< ndiffc >>
rect -47 -753 -13 -719
rect 37 -731 71 -697
rect 121 -753 155 -719
rect 289 -751 323 -717
rect 389 -751 423 -717
rect 479 -680 513 -646
rect 479 -748 513 -714
rect 79 -1471 113 -1437
rect 271 -1499 305 -1465
rect 355 -1499 389 -1465
rect -55 -2421 -21 -2387
rect 29 -2399 63 -2365
rect 113 -2421 147 -2387
rect 281 -2419 315 -2385
rect 381 -2419 415 -2385
rect 471 -2348 505 -2314
rect 471 -2416 505 -2382
rect 71 -3139 105 -3105
rect 263 -3167 297 -3133
rect 347 -3167 381 -3133
rect -45 -3985 -11 -3951
rect 39 -3963 73 -3929
rect 123 -3985 157 -3951
rect 291 -3983 325 -3949
rect 391 -3983 425 -3949
rect 481 -3912 515 -3878
rect 481 -3980 515 -3946
rect 81 -4703 115 -4669
rect 273 -4731 307 -4697
rect 357 -4731 391 -4697
<< pdiffc >>
rect -47 -363 -13 -329
rect -47 -431 -13 -397
rect 121 -373 155 -339
rect 121 -441 155 -407
rect 205 -373 239 -339
rect 205 -441 239 -407
rect 289 -373 323 -339
rect 393 -373 427 -339
rect 393 -441 427 -407
rect 477 -371 511 -337
rect 477 -439 511 -405
rect 477 -507 511 -473
rect 79 -1149 113 -1115
rect 163 -1149 197 -1115
rect 271 -1107 305 -1073
rect 271 -1175 305 -1141
rect 375 -1107 409 -1073
rect 375 -1175 409 -1141
rect -55 -2031 -21 -1997
rect -55 -2099 -21 -2065
rect 113 -2041 147 -2007
rect 113 -2109 147 -2075
rect 197 -2041 231 -2007
rect 197 -2109 231 -2075
rect 281 -2041 315 -2007
rect 385 -2041 419 -2007
rect 385 -2109 419 -2075
rect 469 -2039 503 -2005
rect 469 -2107 503 -2073
rect 469 -2175 503 -2141
rect 71 -2817 105 -2783
rect 155 -2817 189 -2783
rect 263 -2775 297 -2741
rect 263 -2843 297 -2809
rect 367 -2775 401 -2741
rect 367 -2843 401 -2809
rect -45 -3595 -11 -3561
rect -45 -3663 -11 -3629
rect 123 -3605 157 -3571
rect 123 -3673 157 -3639
rect 207 -3605 241 -3571
rect 207 -3673 241 -3639
rect 291 -3605 325 -3571
rect 395 -3605 429 -3571
rect 395 -3673 429 -3639
rect 479 -3603 513 -3569
rect 479 -3671 513 -3637
rect 479 -3739 513 -3705
rect 81 -4381 115 -4347
rect 165 -4381 199 -4347
rect 273 -4339 307 -4305
rect 273 -4407 307 -4373
rect 377 -4339 411 -4305
rect 377 -4407 411 -4373
<< poly >>
rect -3 -317 27 -291
rect 81 -317 111 -291
rect 165 -317 195 -291
rect 249 -317 279 -291
rect 437 -317 467 -291
rect -3 -549 27 -517
rect 81 -549 111 -517
rect 165 -549 195 -517
rect 249 -549 279 -517
rect 437 -549 467 -517
rect -15 -565 39 -549
rect -15 -599 -5 -565
rect 29 -599 39 -565
rect -15 -615 39 -599
rect 81 -565 195 -549
rect 81 -599 112 -565
rect 146 -599 195 -565
rect 81 -615 195 -599
rect 237 -565 291 -549
rect 237 -599 247 -565
rect 281 -599 291 -565
rect 237 -615 291 -599
rect 333 -565 467 -549
rect 333 -599 343 -565
rect 377 -582 467 -565
rect 377 -599 463 -582
rect 333 -615 463 -599
rect -3 -637 27 -615
rect 81 -637 111 -615
rect 165 -637 195 -615
rect 249 -637 279 -615
rect 433 -637 463 -615
rect -3 -793 27 -767
rect 81 -793 111 -767
rect 165 -793 195 -767
rect 249 -793 279 -767
rect 433 -793 463 -767
rect 315 -1061 345 -1035
rect 123 -1103 153 -1077
rect 207 -1103 237 -1077
rect 123 -1293 153 -1187
rect 66 -1309 153 -1293
rect 66 -1343 82 -1309
rect 116 -1343 153 -1309
rect 66 -1359 153 -1343
rect 123 -1399 153 -1359
rect 207 -1293 237 -1187
rect 315 -1293 345 -1261
rect 207 -1309 273 -1293
rect 207 -1343 223 -1309
rect 257 -1343 273 -1309
rect 207 -1359 273 -1343
rect 315 -1309 381 -1293
rect 315 -1343 331 -1309
rect 365 -1343 381 -1309
rect 315 -1359 381 -1343
rect 207 -1399 237 -1359
rect 315 -1381 345 -1359
rect 123 -1509 153 -1483
rect 207 -1509 237 -1483
rect 315 -1537 345 -1511
rect -11 -1985 19 -1959
rect 73 -1985 103 -1959
rect 157 -1985 187 -1959
rect 241 -1985 271 -1959
rect 429 -1985 459 -1959
rect -11 -2217 19 -2185
rect 73 -2217 103 -2185
rect 157 -2217 187 -2185
rect 241 -2217 271 -2185
rect 429 -2217 459 -2185
rect -23 -2233 31 -2217
rect -23 -2267 -13 -2233
rect 21 -2267 31 -2233
rect -23 -2283 31 -2267
rect 73 -2233 187 -2217
rect 73 -2267 104 -2233
rect 138 -2267 187 -2233
rect 73 -2283 187 -2267
rect 229 -2233 283 -2217
rect 229 -2267 239 -2233
rect 273 -2267 283 -2233
rect 229 -2283 283 -2267
rect 325 -2233 459 -2217
rect 325 -2267 335 -2233
rect 369 -2250 459 -2233
rect 369 -2267 455 -2250
rect 325 -2283 455 -2267
rect -11 -2305 19 -2283
rect 73 -2305 103 -2283
rect 157 -2305 187 -2283
rect 241 -2305 271 -2283
rect 425 -2305 455 -2283
rect -11 -2461 19 -2435
rect 73 -2461 103 -2435
rect 157 -2461 187 -2435
rect 241 -2461 271 -2435
rect 425 -2461 455 -2435
rect 307 -2729 337 -2703
rect 115 -2771 145 -2745
rect 199 -2771 229 -2745
rect 115 -2961 145 -2855
rect 58 -2977 145 -2961
rect 58 -3011 74 -2977
rect 108 -3011 145 -2977
rect 58 -3027 145 -3011
rect 115 -3067 145 -3027
rect 199 -2961 229 -2855
rect 307 -2961 337 -2929
rect 199 -2977 265 -2961
rect 199 -3011 215 -2977
rect 249 -3011 265 -2977
rect 199 -3027 265 -3011
rect 307 -2977 373 -2961
rect 307 -3011 323 -2977
rect 357 -3011 373 -2977
rect 307 -3027 373 -3011
rect 199 -3067 229 -3027
rect 307 -3049 337 -3027
rect 115 -3177 145 -3151
rect 199 -3177 229 -3151
rect 307 -3205 337 -3179
rect 1446 -3233 1462 -3208
rect -1 -3549 29 -3523
rect 83 -3549 113 -3523
rect 167 -3549 197 -3523
rect 251 -3549 281 -3523
rect 439 -3549 469 -3523
rect -1 -3781 29 -3749
rect 83 -3781 113 -3749
rect 167 -3781 197 -3749
rect 251 -3781 281 -3749
rect 439 -3781 469 -3749
rect -13 -3797 41 -3781
rect -13 -3831 -3 -3797
rect 31 -3831 41 -3797
rect -13 -3847 41 -3831
rect 83 -3797 197 -3781
rect 83 -3831 114 -3797
rect 148 -3831 197 -3797
rect 83 -3847 197 -3831
rect 239 -3797 293 -3781
rect 239 -3831 249 -3797
rect 283 -3831 293 -3797
rect 239 -3847 293 -3831
rect 335 -3797 469 -3781
rect 335 -3831 345 -3797
rect 379 -3814 469 -3797
rect 379 -3831 465 -3814
rect 335 -3847 465 -3831
rect -1 -3869 29 -3847
rect 83 -3869 113 -3847
rect 167 -3869 197 -3847
rect 251 -3869 281 -3847
rect 435 -3869 465 -3847
rect -1 -4025 29 -3999
rect 83 -4025 113 -3999
rect 167 -4025 197 -3999
rect 251 -4025 281 -3999
rect 435 -4025 465 -3999
rect 317 -4293 347 -4267
rect 125 -4335 155 -4309
rect 209 -4335 239 -4309
rect 125 -4525 155 -4419
rect 68 -4541 155 -4525
rect 68 -4575 84 -4541
rect 118 -4575 155 -4541
rect 68 -4591 155 -4575
rect 125 -4631 155 -4591
rect 209 -4525 239 -4419
rect 317 -4525 347 -4493
rect 209 -4541 275 -4525
rect 209 -4575 225 -4541
rect 259 -4575 275 -4541
rect 209 -4591 275 -4575
rect 317 -4541 383 -4525
rect 317 -4575 333 -4541
rect 367 -4575 383 -4541
rect 317 -4591 383 -4575
rect 209 -4631 239 -4591
rect 317 -4613 347 -4591
rect 125 -4741 155 -4715
rect 209 -4741 239 -4715
rect 317 -4769 347 -4743
<< polycont >>
rect -5 -599 29 -565
rect 112 -599 146 -565
rect 247 -599 281 -565
rect 343 -599 377 -565
rect 82 -1343 116 -1309
rect 223 -1343 257 -1309
rect 331 -1343 365 -1309
rect -13 -2267 21 -2233
rect 104 -2267 138 -2233
rect 239 -2267 273 -2233
rect 335 -2267 369 -2233
rect 74 -3011 108 -2977
rect 215 -3011 249 -2977
rect 323 -3011 357 -2977
rect -3 -3831 31 -3797
rect 114 -3831 148 -3797
rect 249 -3831 283 -3797
rect 345 -3831 379 -3797
rect 84 -4575 118 -4541
rect 225 -4575 259 -4541
rect 333 -4575 367 -4541
<< locali >>
rect -90 -287 -61 -253
rect -27 -287 31 -253
rect 65 -287 123 -253
rect 157 -287 215 -253
rect 249 -287 307 -253
rect 341 -287 399 -253
rect 433 -287 491 -253
rect 525 -287 554 -253
rect -73 -329 3 -321
rect -73 -363 -47 -329
rect -13 -363 3 -329
rect -73 -397 3 -363
rect -73 -431 -47 -397
rect -13 -431 3 -397
rect -73 -457 3 -431
rect 121 -339 155 -287
rect 121 -407 155 -373
rect 121 -457 155 -441
rect 189 -339 255 -321
rect 189 -373 205 -339
rect 239 -373 255 -339
rect 189 -407 255 -373
rect 289 -339 323 -287
rect 289 -389 323 -373
rect 357 -339 437 -321
rect 357 -373 393 -339
rect 427 -373 437 -339
rect 189 -441 205 -407
rect 239 -423 255 -407
rect 357 -407 437 -373
rect 357 -423 393 -407
rect 239 -441 393 -423
rect 427 -441 437 -407
rect 189 -457 437 -441
rect 473 -337 537 -321
rect 473 -371 477 -337
rect 511 -362 537 -337
rect 473 -396 488 -371
rect 522 -396 537 -362
rect 473 -405 537 -396
rect 473 -439 477 -405
rect 511 -439 537 -405
rect -73 -649 -39 -457
rect 473 -473 537 -439
rect -5 -525 256 -491
rect 473 -507 477 -473
rect 511 -507 537 -473
rect -5 -564 44 -525
rect -5 -565 -4 -564
rect 30 -598 44 -564
rect 29 -599 44 -598
rect 78 -562 188 -559
rect 78 -565 116 -562
rect 78 -599 112 -565
rect 150 -596 188 -562
rect 146 -599 188 -596
rect 222 -565 256 -525
rect 411 -541 537 -507
rect 331 -565 377 -549
rect 222 -599 247 -565
rect 281 -599 297 -565
rect 331 -599 343 -565
rect -5 -615 44 -599
rect 331 -649 377 -599
rect -73 -683 377 -649
rect 37 -697 71 -683
rect -63 -753 -47 -719
rect -13 -753 3 -719
rect 411 -717 445 -541
rect 37 -747 71 -731
rect -63 -797 3 -753
rect 105 -753 121 -719
rect 155 -753 171 -719
rect 254 -751 289 -717
rect 323 -751 389 -717
rect 423 -751 445 -717
rect 479 -646 537 -630
rect 513 -680 537 -646
rect 479 -714 537 -680
rect 513 -748 537 -714
rect 105 -797 171 -753
rect 479 -797 537 -748
rect -90 -831 -61 -797
rect -27 -831 31 -797
rect 65 -831 123 -797
rect 157 -831 215 -797
rect 249 -831 307 -797
rect 341 -831 399 -797
rect 433 -831 491 -797
rect 525 -831 554 -797
rect 8 -1031 37 -997
rect 71 -1031 129 -997
rect 163 -1031 221 -997
rect 255 -1031 313 -997
rect 347 -1031 405 -997
rect 439 -1031 468 -997
rect 65 -1115 121 -1031
rect 255 -1073 321 -1031
rect 65 -1149 79 -1115
rect 113 -1149 121 -1115
rect 65 -1165 121 -1149
rect 155 -1115 215 -1099
rect 155 -1149 163 -1115
rect 197 -1149 215 -1115
rect 155 -1209 215 -1149
rect 255 -1107 271 -1073
rect 305 -1107 321 -1073
rect 255 -1141 321 -1107
rect 255 -1175 271 -1141
rect 305 -1175 321 -1141
rect 359 -1073 451 -1065
rect 359 -1107 375 -1073
rect 409 -1107 451 -1073
rect 359 -1141 451 -1107
rect 359 -1175 375 -1141
rect 409 -1175 451 -1141
rect 28 -1286 81 -1221
rect 155 -1243 343 -1209
rect 28 -1326 30 -1286
rect 72 -1293 81 -1286
rect 309 -1293 343 -1243
rect 72 -1309 163 -1293
rect 72 -1326 82 -1309
rect 28 -1343 82 -1326
rect 116 -1343 163 -1309
rect 207 -1296 275 -1293
rect 207 -1336 220 -1296
rect 262 -1336 275 -1296
rect 207 -1343 223 -1336
rect 257 -1343 275 -1336
rect 309 -1309 367 -1293
rect 309 -1343 331 -1309
rect 365 -1343 367 -1309
rect 309 -1359 367 -1343
rect 309 -1377 343 -1359
rect 65 -1415 343 -1377
rect 401 -1408 451 -1175
rect 65 -1437 131 -1415
rect 65 -1471 79 -1437
rect 113 -1471 131 -1437
rect 401 -1442 410 -1408
rect 446 -1442 451 -1408
rect 401 -1449 451 -1442
rect 65 -1487 131 -1471
rect 255 -1465 305 -1449
rect 255 -1499 271 -1465
rect 255 -1541 305 -1499
rect 339 -1465 451 -1449
rect 339 -1499 355 -1465
rect 389 -1499 451 -1465
rect 339 -1507 451 -1499
rect 8 -1575 37 -1541
rect 71 -1575 129 -1541
rect 163 -1575 221 -1541
rect 255 -1575 313 -1541
rect 347 -1575 405 -1541
rect 439 -1575 468 -1541
rect -98 -1955 -69 -1921
rect -35 -1955 23 -1921
rect 57 -1955 115 -1921
rect 149 -1955 207 -1921
rect 241 -1955 299 -1921
rect 333 -1955 391 -1921
rect 425 -1955 483 -1921
rect 517 -1955 546 -1921
rect -81 -1997 -5 -1989
rect -81 -2031 -55 -1997
rect -21 -2031 -5 -1997
rect -81 -2065 -5 -2031
rect -81 -2099 -55 -2065
rect -21 -2099 -5 -2065
rect -81 -2125 -5 -2099
rect 113 -2007 147 -1955
rect 113 -2075 147 -2041
rect 113 -2125 147 -2109
rect 181 -2007 247 -1989
rect 181 -2041 197 -2007
rect 231 -2041 247 -2007
rect 181 -2075 247 -2041
rect 281 -2007 315 -1955
rect 281 -2057 315 -2041
rect 349 -2007 429 -1989
rect 349 -2041 385 -2007
rect 419 -2041 429 -2007
rect 181 -2109 197 -2075
rect 231 -2091 247 -2075
rect 349 -2075 429 -2041
rect 349 -2091 385 -2075
rect 231 -2109 385 -2091
rect 419 -2109 429 -2075
rect 181 -2125 429 -2109
rect 465 -2005 529 -1989
rect 465 -2039 469 -2005
rect 503 -2039 529 -2005
rect 465 -2072 529 -2039
rect 465 -2073 480 -2072
rect 465 -2107 469 -2073
rect 514 -2106 529 -2072
rect 503 -2107 529 -2106
rect -81 -2317 -47 -2125
rect 465 -2141 529 -2107
rect -13 -2193 248 -2159
rect 465 -2175 469 -2141
rect 503 -2175 529 -2141
rect -13 -2232 36 -2193
rect -13 -2233 -12 -2232
rect 22 -2266 36 -2232
rect 21 -2267 36 -2266
rect 70 -2230 180 -2227
rect 70 -2233 108 -2230
rect 70 -2267 104 -2233
rect 142 -2264 180 -2230
rect 138 -2267 180 -2264
rect 214 -2233 248 -2193
rect 403 -2209 529 -2175
rect 323 -2233 369 -2217
rect 214 -2267 239 -2233
rect 273 -2267 289 -2233
rect 323 -2267 335 -2233
rect -13 -2283 36 -2267
rect 323 -2317 369 -2267
rect -81 -2351 369 -2317
rect 29 -2365 63 -2351
rect -71 -2421 -55 -2387
rect -21 -2421 -5 -2387
rect 403 -2385 437 -2209
rect 29 -2415 63 -2399
rect -71 -2465 -5 -2421
rect 97 -2421 113 -2387
rect 147 -2421 163 -2387
rect 246 -2419 281 -2385
rect 315 -2419 381 -2385
rect 415 -2419 437 -2385
rect 471 -2314 529 -2298
rect 505 -2348 529 -2314
rect 471 -2382 529 -2348
rect 505 -2416 529 -2382
rect 97 -2465 163 -2421
rect 471 -2465 529 -2416
rect -98 -2499 -69 -2465
rect -35 -2499 23 -2465
rect 57 -2499 115 -2465
rect 149 -2499 207 -2465
rect 241 -2499 299 -2465
rect 333 -2499 391 -2465
rect 425 -2499 483 -2465
rect 517 -2499 546 -2465
rect 0 -2699 29 -2665
rect 63 -2699 121 -2665
rect 155 -2699 213 -2665
rect 247 -2699 305 -2665
rect 339 -2699 397 -2665
rect 431 -2699 460 -2665
rect 57 -2783 113 -2699
rect 247 -2741 313 -2699
rect 57 -2817 71 -2783
rect 105 -2817 113 -2783
rect 57 -2833 113 -2817
rect 147 -2783 207 -2767
rect 147 -2817 155 -2783
rect 189 -2817 207 -2783
rect 147 -2877 207 -2817
rect 247 -2775 263 -2741
rect 297 -2775 313 -2741
rect 247 -2809 313 -2775
rect 247 -2843 263 -2809
rect 297 -2843 313 -2809
rect 351 -2741 443 -2733
rect 351 -2775 367 -2741
rect 401 -2775 443 -2741
rect 351 -2809 443 -2775
rect 351 -2843 367 -2809
rect 401 -2843 443 -2809
rect 20 -2954 73 -2889
rect 147 -2911 335 -2877
rect 20 -2994 22 -2954
rect 64 -2961 73 -2954
rect 301 -2961 335 -2911
rect 393 -2922 443 -2843
rect 393 -2956 402 -2922
rect 438 -2956 443 -2922
rect 64 -2977 155 -2961
rect 64 -2994 74 -2977
rect 20 -3011 74 -2994
rect 108 -3011 155 -2977
rect 199 -2964 267 -2961
rect 199 -3004 212 -2964
rect 254 -3004 267 -2964
rect 199 -3011 215 -3004
rect 249 -3011 267 -3004
rect 301 -2977 359 -2961
rect 301 -3011 323 -2977
rect 357 -3011 359 -2977
rect 301 -3027 359 -3011
rect 301 -3045 335 -3027
rect 57 -3083 335 -3045
rect 57 -3105 123 -3083
rect 57 -3139 71 -3105
rect 105 -3139 123 -3105
rect 393 -3117 443 -2956
rect 57 -3155 123 -3139
rect 247 -3133 297 -3117
rect 247 -3167 263 -3133
rect 247 -3209 297 -3167
rect 331 -3133 443 -3117
rect 331 -3167 347 -3133
rect 381 -3167 443 -3133
rect 331 -3175 443 -3167
rect 0 -3243 29 -3209
rect 63 -3243 121 -3209
rect 155 -3243 213 -3209
rect 247 -3243 305 -3209
rect 339 -3243 397 -3209
rect 431 -3243 460 -3209
rect -88 -3519 -59 -3485
rect -25 -3519 33 -3485
rect 67 -3519 125 -3485
rect 159 -3519 217 -3485
rect 251 -3519 309 -3485
rect 343 -3519 401 -3485
rect 435 -3519 493 -3485
rect 527 -3519 556 -3485
rect -71 -3561 5 -3553
rect -71 -3595 -45 -3561
rect -11 -3595 5 -3561
rect -71 -3629 5 -3595
rect -71 -3663 -45 -3629
rect -11 -3663 5 -3629
rect -71 -3689 5 -3663
rect 123 -3571 157 -3519
rect 123 -3639 157 -3605
rect 123 -3689 157 -3673
rect 191 -3571 257 -3553
rect 191 -3605 207 -3571
rect 241 -3605 257 -3571
rect 191 -3639 257 -3605
rect 291 -3571 325 -3519
rect 291 -3621 325 -3605
rect 359 -3571 439 -3553
rect 359 -3605 395 -3571
rect 429 -3605 439 -3571
rect 191 -3673 207 -3639
rect 241 -3655 257 -3639
rect 359 -3639 439 -3605
rect 359 -3655 395 -3639
rect 241 -3673 395 -3655
rect 429 -3673 439 -3639
rect 191 -3689 439 -3673
rect 475 -3569 539 -3553
rect 475 -3603 479 -3569
rect 513 -3603 539 -3569
rect 475 -3636 539 -3603
rect 475 -3637 480 -3636
rect 475 -3671 479 -3637
rect 516 -3670 539 -3636
rect 513 -3671 539 -3670
rect -71 -3881 -37 -3689
rect 475 -3705 539 -3671
rect -3 -3757 258 -3723
rect 475 -3739 479 -3705
rect 513 -3739 539 -3705
rect -3 -3796 46 -3757
rect -3 -3797 -2 -3796
rect 32 -3830 46 -3796
rect 31 -3831 46 -3830
rect 80 -3794 190 -3791
rect 80 -3797 118 -3794
rect 80 -3831 114 -3797
rect 152 -3828 190 -3794
rect 148 -3831 190 -3828
rect 224 -3797 258 -3757
rect 413 -3773 539 -3739
rect 333 -3797 379 -3781
rect 224 -3831 249 -3797
rect 283 -3831 299 -3797
rect 333 -3831 345 -3797
rect -3 -3847 46 -3831
rect 333 -3881 379 -3831
rect -71 -3915 379 -3881
rect 39 -3929 73 -3915
rect -61 -3985 -45 -3951
rect -11 -3985 5 -3951
rect 413 -3949 447 -3773
rect 39 -3979 73 -3963
rect -61 -4029 5 -3985
rect 107 -3985 123 -3951
rect 157 -3985 173 -3951
rect 256 -3983 291 -3949
rect 325 -3983 391 -3949
rect 425 -3983 447 -3949
rect 481 -3878 539 -3862
rect 515 -3912 539 -3878
rect 481 -3946 539 -3912
rect 515 -3980 539 -3946
rect 107 -4029 173 -3985
rect 481 -4029 539 -3980
rect -88 -4063 -59 -4029
rect -25 -4063 33 -4029
rect 67 -4063 125 -4029
rect 159 -4063 217 -4029
rect 251 -4063 309 -4029
rect 343 -4063 401 -4029
rect 435 -4063 493 -4029
rect 527 -4063 556 -4029
rect 10 -4263 39 -4229
rect 73 -4263 131 -4229
rect 165 -4263 223 -4229
rect 257 -4263 315 -4229
rect 349 -4263 407 -4229
rect 441 -4263 470 -4229
rect 67 -4347 123 -4263
rect 257 -4305 323 -4263
rect 67 -4381 81 -4347
rect 115 -4381 123 -4347
rect 67 -4397 123 -4381
rect 157 -4347 217 -4331
rect 157 -4381 165 -4347
rect 199 -4381 217 -4347
rect 157 -4441 217 -4381
rect 257 -4339 273 -4305
rect 307 -4339 323 -4305
rect 257 -4373 323 -4339
rect 257 -4407 273 -4373
rect 307 -4407 323 -4373
rect 361 -4305 453 -4297
rect 361 -4339 377 -4305
rect 411 -4339 453 -4305
rect 361 -4373 453 -4339
rect 361 -4407 377 -4373
rect 411 -4407 453 -4373
rect 30 -4518 83 -4453
rect 157 -4475 345 -4441
rect 30 -4558 32 -4518
rect 74 -4525 83 -4518
rect 311 -4525 345 -4475
rect 74 -4541 165 -4525
rect 74 -4558 84 -4541
rect 30 -4575 84 -4558
rect 118 -4575 165 -4541
rect 209 -4528 277 -4525
rect 209 -4568 222 -4528
rect 264 -4568 277 -4528
rect 209 -4575 225 -4568
rect 259 -4575 277 -4568
rect 311 -4541 369 -4525
rect 311 -4575 333 -4541
rect 367 -4575 369 -4541
rect 311 -4591 369 -4575
rect 311 -4609 345 -4591
rect 67 -4647 345 -4609
rect 67 -4669 133 -4647
rect 67 -4703 81 -4669
rect 115 -4703 133 -4669
rect 403 -4681 453 -4407
rect 67 -4719 133 -4703
rect 257 -4697 307 -4681
rect 257 -4731 273 -4697
rect 257 -4773 307 -4731
rect 341 -4697 453 -4681
rect 341 -4731 357 -4697
rect 391 -4731 453 -4697
rect 341 -4739 453 -4731
rect 10 -4807 39 -4773
rect 73 -4807 131 -4773
rect 165 -4807 223 -4773
rect 257 -4807 315 -4773
rect 349 -4807 407 -4773
rect 441 -4807 470 -4773
<< viali >>
rect 476 1060 510 1098
rect -14 966 20 1000
rect 106 968 140 1002
rect 20 238 62 278
rect 210 228 252 268
rect 402 164 438 198
rect 2064 72 2100 108
rect 2236 106 2270 142
rect 2622 106 2656 140
rect 2430 52 2464 88
rect 2334 -16 2368 18
rect 1576 -180 1616 -144
rect -61 -287 -27 -253
rect 31 -287 65 -253
rect 123 -287 157 -253
rect 215 -287 249 -253
rect 307 -287 341 -253
rect 399 -287 433 -253
rect 491 -287 525 -253
rect 488 -371 511 -362
rect 511 -371 522 -362
rect 488 -396 522 -371
rect 1256 -388 1290 -354
rect 1396 -388 1432 -354
rect -4 -565 30 -564
rect -4 -598 29 -565
rect 29 -598 30 -565
rect 116 -565 150 -562
rect 116 -596 146 -565
rect 146 -596 150 -565
rect -61 -831 -27 -797
rect 31 -831 65 -797
rect 123 -831 157 -797
rect 215 -831 249 -797
rect 307 -831 341 -797
rect 399 -831 433 -797
rect 491 -831 525 -797
rect 37 -1031 71 -997
rect 129 -1031 163 -997
rect 221 -1031 255 -997
rect 313 -1031 347 -997
rect 405 -1031 439 -997
rect 3328 -1160 3364 -1126
rect 30 -1326 72 -1286
rect 220 -1309 262 -1296
rect 220 -1336 223 -1309
rect 223 -1336 257 -1309
rect 257 -1336 262 -1309
rect 1282 -1350 1316 -1316
rect 1644 -1360 1680 -1322
rect 1550 -1406 1584 -1372
rect 3312 -1374 3362 -1332
rect 3484 -1372 3522 -1336
rect 410 -1442 446 -1408
rect 1452 -1446 1486 -1412
rect 1826 -1478 1864 -1440
rect 37 -1575 71 -1541
rect 129 -1575 163 -1541
rect 221 -1575 255 -1541
rect 313 -1575 347 -1541
rect 405 -1575 439 -1541
rect 2594 -1562 2628 -1528
rect 2444 -1722 2478 -1688
rect 2266 -1772 2300 -1738
rect -69 -1955 -35 -1921
rect 23 -1955 57 -1921
rect 115 -1955 149 -1921
rect 207 -1955 241 -1921
rect 299 -1955 333 -1921
rect 391 -1955 425 -1921
rect 483 -1955 517 -1921
rect 1578 -1994 1614 -1958
rect 1774 -2052 1812 -2014
rect 480 -2073 514 -2072
rect 480 -2106 503 -2073
rect 503 -2106 514 -2073
rect -12 -2233 22 -2232
rect -12 -2266 21 -2233
rect 21 -2266 22 -2233
rect 108 -2233 142 -2230
rect 108 -2264 138 -2233
rect 138 -2264 142 -2233
rect 1426 -2266 1460 -2232
rect 1628 -2260 1664 -2226
rect -69 -2499 -35 -2465
rect 23 -2499 57 -2465
rect 115 -2499 149 -2465
rect 207 -2499 241 -2465
rect 299 -2499 333 -2465
rect 391 -2499 425 -2465
rect 483 -2499 517 -2465
rect 29 -2699 63 -2665
rect 121 -2699 155 -2665
rect 213 -2699 247 -2665
rect 305 -2699 339 -2665
rect 397 -2699 431 -2665
rect 22 -2994 64 -2954
rect 402 -2956 438 -2922
rect 212 -2977 254 -2964
rect 212 -3004 215 -2977
rect 215 -3004 249 -2977
rect 249 -3004 254 -2977
rect 1778 -3130 1812 -3096
rect 29 -3243 63 -3209
rect 121 -3243 155 -3209
rect 213 -3243 247 -3209
rect 305 -3243 339 -3209
rect 397 -3243 431 -3209
rect 1450 -3214 1486 -3180
rect 1590 -3216 1626 -3182
rect -59 -3519 -25 -3485
rect 33 -3519 67 -3485
rect 125 -3519 159 -3485
rect 217 -3519 251 -3485
rect 309 -3519 343 -3485
rect 401 -3519 435 -3485
rect 493 -3519 527 -3485
rect 480 -3637 516 -3636
rect 480 -3670 513 -3637
rect 513 -3670 516 -3637
rect -2 -3797 32 -3796
rect -2 -3830 31 -3797
rect 31 -3830 32 -3797
rect 118 -3797 152 -3794
rect 118 -3828 148 -3797
rect 148 -3828 152 -3797
rect -59 -4063 -25 -4029
rect 33 -4063 67 -4029
rect 125 -4063 159 -4029
rect 217 -4063 251 -4029
rect 309 -4063 343 -4029
rect 401 -4063 435 -4029
rect 493 -4063 527 -4029
rect 39 -4263 73 -4229
rect 131 -4263 165 -4229
rect 223 -4263 257 -4229
rect 315 -4263 349 -4229
rect 407 -4263 441 -4229
rect 32 -4558 74 -4518
rect 222 -4541 264 -4528
rect 222 -4568 225 -4541
rect 225 -4568 259 -4541
rect 259 -4568 264 -4541
rect 39 -4807 73 -4773
rect 131 -4807 165 -4773
rect 223 -4807 257 -4773
rect 315 -4807 349 -4773
rect 407 -4807 441 -4773
<< metal1 >>
rect -22 1000 38 1276
rect 1378 1114 1580 1146
rect 1378 1112 1438 1114
rect 464 1098 1438 1112
rect 464 1060 476 1098
rect 510 1060 1438 1098
rect 464 1048 1438 1060
rect 1508 1112 1580 1114
rect 1508 1048 1691 1112
rect 464 1046 1691 1048
rect 1378 1020 1580 1046
rect -22 966 -14 1000
rect 20 966 38 1000
rect -22 946 38 966
rect 68 1002 178 1016
rect 68 968 106 1002
rect 140 968 178 1002
rect 68 960 178 968
rect 102 702 133 960
rect 6 502 82 516
rect 6 278 82 294
rect 208 278 262 524
rect 1625 341 1691 1046
rect 6 238 20 278
rect 62 238 82 278
rect 6 222 82 238
rect 198 268 266 278
rect 1625 275 2479 341
rect 2223 272 2289 275
rect 198 228 210 268
rect 252 228 266 268
rect 16 36 70 222
rect 198 216 266 228
rect 390 210 476 218
rect 390 198 408 210
rect 390 164 402 198
rect 390 156 408 164
rect 462 156 476 210
rect 390 144 476 156
rect 626 166 2288 224
rect 626 160 2289 166
rect 198 -8 266 56
rect -90 -253 554 -222
rect -90 -287 -61 -253
rect -27 -287 31 -253
rect 65 -287 123 -253
rect 157 -287 215 -253
rect 249 -287 307 -253
rect 341 -287 399 -253
rect 433 -287 491 -253
rect 525 -287 554 -253
rect -90 -318 554 -287
rect -12 -564 48 -318
rect 626 -350 690 160
rect 2223 142 2289 160
rect 2046 108 2114 132
rect 2046 72 2064 108
rect 2100 72 2114 108
rect 2223 106 2236 142
rect 2270 106 2289 142
rect 2223 98 2289 106
rect 2046 50 2114 72
rect 2413 88 2479 275
rect 2610 148 2666 152
rect 2610 140 2832 148
rect 2610 106 2622 140
rect 2656 106 2832 140
rect 2610 98 2832 106
rect 2610 94 2666 98
rect 2413 52 2430 88
rect 2464 52 2479 88
rect 2322 22 2380 38
rect 1780 18 2380 22
rect 1780 -16 2334 18
rect 2368 -16 2380 18
rect 1780 -22 2380 -16
rect 1782 -136 1862 -22
rect 2322 -28 2380 -22
rect 2413 -26 2479 52
rect 1536 -144 1862 -136
rect 472 -362 690 -350
rect 472 -396 488 -362
rect 522 -396 690 -362
rect 472 -414 690 -396
rect 722 -212 1452 -160
rect 1536 -180 1576 -144
rect 1616 -180 1862 -144
rect 1536 -194 1862 -180
rect -12 -598 -4 -564
rect 30 -598 48 -564
rect -12 -618 48 -598
rect 78 -562 188 -548
rect 78 -596 116 -562
rect 150 -596 188 -562
rect 78 -604 188 -596
rect 112 -766 143 -604
rect -90 -797 554 -766
rect -90 -831 -61 -797
rect -27 -831 31 -797
rect 65 -831 123 -797
rect 157 -831 215 -797
rect 249 -831 307 -797
rect 341 -831 399 -797
rect 433 -831 491 -797
rect 525 -831 554 -797
rect -90 -862 554 -831
rect 8 -997 468 -966
rect 8 -1031 37 -997
rect 71 -1031 129 -997
rect 163 -1031 221 -997
rect 255 -1031 313 -997
rect 347 -1031 405 -997
rect 439 -1031 468 -997
rect 8 -1062 468 -1031
rect 16 -1286 92 -1268
rect 220 -1286 266 -1062
rect 16 -1326 30 -1286
rect 72 -1326 92 -1286
rect 16 -1342 92 -1326
rect 208 -1296 276 -1286
rect 208 -1336 220 -1296
rect 262 -1336 276 -1296
rect 24 -1510 78 -1342
rect 208 -1348 276 -1336
rect 398 -1392 570 -1378
rect 398 -1408 462 -1392
rect 398 -1442 410 -1408
rect 446 -1442 462 -1408
rect 398 -1454 462 -1442
rect 522 -1454 570 -1392
rect 398 -1472 570 -1454
rect 8 -1541 468 -1510
rect 8 -1575 37 -1541
rect 71 -1575 129 -1541
rect 163 -1575 221 -1541
rect 255 -1575 313 -1541
rect 347 -1575 405 -1541
rect 439 -1575 468 -1541
rect 8 -1606 468 -1575
rect -98 -1921 546 -1890
rect -98 -1955 -69 -1921
rect -35 -1955 23 -1921
rect 57 -1955 115 -1921
rect 149 -1955 207 -1921
rect 241 -1955 299 -1921
rect 333 -1955 391 -1921
rect 425 -1955 483 -1921
rect 517 -1955 546 -1921
rect -98 -1986 546 -1955
rect 722 -1926 774 -212
rect 1400 -336 1452 -212
rect 1202 -341 1338 -340
rect 994 -354 1338 -341
rect 994 -388 1256 -354
rect 1290 -388 1338 -354
rect 994 -414 1338 -388
rect 1372 -354 1452 -336
rect 1372 -388 1396 -354
rect 1432 -388 1452 -354
rect 1372 -402 1452 -388
rect 994 -419 1277 -414
rect 994 -1321 1072 -419
rect 2779 -1115 2829 98
rect 2779 -1120 2830 -1115
rect 2779 -1126 3506 -1120
rect 2779 -1160 3328 -1126
rect 3364 -1160 3506 -1126
rect 2779 -1167 3506 -1160
rect 2822 -1168 3506 -1167
rect 2878 -1262 3546 -1202
rect 1255 -1316 1333 -1263
rect 2878 -1274 2952 -1262
rect 1255 -1321 1282 -1316
rect 994 -1350 1282 -1321
rect 1316 -1350 1333 -1316
rect 994 -1399 1333 -1350
rect 722 -1936 808 -1926
rect -20 -2232 40 -1986
rect 722 -1988 730 -1936
rect 792 -1988 808 -1936
rect 722 -1996 808 -1988
rect 722 -2064 774 -1996
rect 468 -2072 774 -2064
rect 468 -2106 480 -2072
rect 514 -2106 774 -2072
rect 468 -2116 774 -2106
rect 994 -2207 1072 -1399
rect 1434 -1402 1504 -1356
rect 1434 -1454 1444 -1402
rect 1496 -1454 1504 -1402
rect 1434 -1494 1504 -1454
rect 1532 -1362 1600 -1306
rect 1532 -1414 1542 -1362
rect 1594 -1414 1600 -1362
rect 1532 -1492 1600 -1414
rect 1634 -1322 1706 -1304
rect 1634 -1360 1644 -1322
rect 1680 -1360 1706 -1322
rect 1634 -1406 1706 -1360
rect 1634 -1462 1640 -1406
rect 1692 -1462 1706 -1406
rect 2878 -1362 2950 -1274
rect 3268 -1312 3408 -1300
rect 1634 -1488 1706 -1462
rect 1812 -1440 2098 -1420
rect 1812 -1478 1826 -1440
rect 1864 -1478 2098 -1440
rect 1812 -1494 2098 -1478
rect 2017 -1507 2098 -1494
rect 2878 -1506 2948 -1362
rect 3268 -1388 3298 -1312
rect 3378 -1334 3408 -1312
rect 3474 -1320 3546 -1262
rect 3378 -1388 3406 -1334
rect 3452 -1336 3546 -1320
rect 3452 -1372 3484 -1336
rect 3522 -1372 3546 -1336
rect 3452 -1388 3546 -1372
rect 3268 -1402 3406 -1388
rect 2017 -1581 2495 -1507
rect 2552 -1528 2948 -1506
rect 2552 -1562 2594 -1528
rect 2628 -1562 2948 -1528
rect 2552 -1578 2948 -1562
rect 2421 -1688 2495 -1581
rect 1976 -1738 2325 -1715
rect 1976 -1772 2266 -1738
rect 2300 -1772 2325 -1738
rect 1976 -1789 2325 -1772
rect 2421 -1722 2444 -1688
rect 2478 -1722 2495 -1688
rect 1552 -1954 1650 -1948
rect 1552 -2006 1572 -1954
rect 1626 -2006 1650 -1954
rect 1976 -1994 2050 -1789
rect 2421 -1803 2495 -1722
rect 1552 -2024 1650 -2006
rect 1764 -2014 2050 -1994
rect 1764 -2052 1774 -2014
rect 1812 -2052 2050 -2014
rect 1764 -2068 2050 -2052
rect -20 -2266 -12 -2232
rect 22 -2266 40 -2232
rect -20 -2286 40 -2266
rect 70 -2230 180 -2216
rect 70 -2264 108 -2230
rect 142 -2264 180 -2230
rect 70 -2272 180 -2264
rect 994 -2232 1513 -2207
rect 994 -2266 1426 -2232
rect 1460 -2266 1513 -2232
rect 104 -2434 135 -2272
rect 994 -2285 1513 -2266
rect 1608 -2210 1690 -2138
rect 1608 -2264 1628 -2210
rect 1680 -2264 1690 -2210
rect -98 -2465 546 -2434
rect -98 -2499 -69 -2465
rect -35 -2499 23 -2465
rect 57 -2499 115 -2465
rect 149 -2499 207 -2465
rect 241 -2499 299 -2465
rect 333 -2499 391 -2465
rect 425 -2499 483 -2465
rect 517 -2499 546 -2465
rect -98 -2530 546 -2499
rect 0 -2665 460 -2634
rect 0 -2699 29 -2665
rect 63 -2699 121 -2665
rect 155 -2699 213 -2665
rect 247 -2699 305 -2665
rect 339 -2699 397 -2665
rect 431 -2699 460 -2665
rect 0 -2730 460 -2699
rect 8 -2954 84 -2928
rect 208 -2954 258 -2730
rect 392 -2902 542 -2888
rect 392 -2922 438 -2902
rect 8 -2994 22 -2954
rect 64 -2994 84 -2954
rect 8 -3010 84 -2994
rect 200 -2964 268 -2954
rect 200 -3004 212 -2964
rect 254 -3004 268 -2964
rect 392 -2956 402 -2922
rect 392 -2970 438 -2956
rect 500 -2970 542 -2902
rect 392 -2986 542 -2970
rect 22 -3178 74 -3010
rect 200 -3016 268 -3004
rect 994 -3171 1072 -2285
rect 1608 -2322 1690 -2264
rect 1766 -3084 1834 -3074
rect 1766 -3136 1772 -3084
rect 1824 -3136 1834 -3084
rect 1766 -3142 1834 -3136
rect 0 -3209 460 -3178
rect 0 -3243 29 -3209
rect 63 -3243 121 -3209
rect 155 -3243 213 -3209
rect 247 -3243 305 -3209
rect 339 -3243 397 -3209
rect 431 -3243 460 -3209
rect 0 -3274 460 -3243
rect 994 -3180 1527 -3171
rect 994 -3214 1450 -3180
rect 1486 -3214 1527 -3180
rect 994 -3249 1527 -3214
rect 1574 -3174 1644 -3166
rect 1574 -3226 1582 -3174
rect 1634 -3226 1644 -3174
rect 1574 -3232 1644 -3226
rect -88 -3485 556 -3454
rect -88 -3519 -59 -3485
rect -25 -3519 33 -3485
rect 67 -3519 125 -3485
rect 159 -3519 217 -3485
rect 251 -3519 309 -3485
rect 343 -3519 401 -3485
rect 435 -3519 493 -3485
rect 527 -3519 556 -3485
rect -88 -3550 556 -3519
rect -10 -3796 50 -3550
rect 994 -3622 1072 -3249
rect 474 -3636 1072 -3622
rect 474 -3670 480 -3636
rect 516 -3670 1072 -3636
rect 474 -3700 1072 -3670
rect -10 -3830 -2 -3796
rect 32 -3830 50 -3796
rect -10 -3850 50 -3830
rect 80 -3794 190 -3780
rect 80 -3828 118 -3794
rect 152 -3828 190 -3794
rect 80 -3836 190 -3828
rect 114 -3998 145 -3836
rect -88 -4029 556 -3998
rect -88 -4063 -59 -4029
rect -25 -4063 33 -4029
rect 67 -4063 125 -4029
rect 159 -4063 217 -4029
rect 251 -4063 309 -4029
rect 343 -4063 401 -4029
rect 435 -4063 493 -4029
rect 527 -4063 556 -4029
rect -88 -4094 556 -4063
rect 10 -4229 470 -4198
rect 10 -4263 39 -4229
rect 73 -4263 131 -4229
rect 165 -4263 223 -4229
rect 257 -4263 315 -4229
rect 349 -4263 407 -4229
rect 441 -4263 470 -4229
rect 10 -4294 470 -4263
rect 18 -4518 94 -4506
rect 18 -4558 32 -4518
rect 74 -4558 94 -4518
rect 18 -4574 94 -4558
rect 208 -4528 280 -4294
rect 208 -4562 222 -4528
rect 210 -4568 222 -4562
rect 264 -4562 280 -4528
rect 264 -4568 278 -4562
rect 38 -4742 88 -4574
rect 210 -4584 278 -4568
rect 210 -4742 278 -4738
rect 10 -4773 470 -4742
rect 10 -4807 39 -4773
rect 73 -4807 131 -4773
rect 165 -4807 223 -4773
rect 257 -4807 315 -4773
rect 349 -4807 407 -4773
rect 441 -4807 470 -4773
rect 10 -4838 470 -4807
<< via1 >>
rect 1438 1048 1508 1114
rect 408 198 462 210
rect 408 164 438 198
rect 438 164 462 198
rect 408 156 462 164
rect 462 -1454 522 -1392
rect 730 -1988 792 -1936
rect 1444 -1412 1496 -1402
rect 1444 -1446 1452 -1412
rect 1452 -1446 1486 -1412
rect 1486 -1446 1496 -1412
rect 1444 -1454 1496 -1446
rect 1542 -1372 1594 -1362
rect 1542 -1406 1550 -1372
rect 1550 -1406 1584 -1372
rect 1584 -1406 1594 -1372
rect 1542 -1414 1594 -1406
rect 1640 -1462 1692 -1406
rect 3298 -1332 3378 -1312
rect 3298 -1374 3312 -1332
rect 3312 -1374 3362 -1332
rect 3362 -1374 3378 -1332
rect 3298 -1388 3378 -1374
rect 1572 -1958 1626 -1954
rect 1572 -1994 1578 -1958
rect 1578 -1994 1614 -1958
rect 1614 -1994 1626 -1958
rect 1572 -2006 1626 -1994
rect 1628 -2226 1680 -2210
rect 1628 -2260 1664 -2226
rect 1664 -2260 1680 -2226
rect 1628 -2264 1680 -2260
rect 438 -2970 500 -2902
rect 1772 -3096 1824 -3084
rect 1772 -3130 1778 -3096
rect 1778 -3130 1812 -3096
rect 1812 -3130 1824 -3096
rect 1772 -3136 1824 -3130
rect 1582 -3182 1634 -3174
rect 1582 -3216 1590 -3182
rect 1590 -3216 1626 -3182
rect 1626 -3216 1634 -3182
rect 1582 -3226 1634 -3216
<< metal2 >>
rect 1378 1114 1580 1146
rect 1378 1048 1438 1114
rect 1508 1048 1580 1114
rect 1378 1020 1580 1048
rect 390 210 498 218
rect 390 156 408 210
rect 462 180 498 210
rect 462 156 890 180
rect 390 144 890 156
rect 854 -1194 890 144
rect 1442 -782 1510 1020
rect 1442 -850 1600 -782
rect 854 -1230 1464 -1194
rect 1428 -1356 1464 -1230
rect 400 -1392 570 -1380
rect 400 -1454 462 -1392
rect 522 -1412 570 -1392
rect 1428 -1402 1504 -1356
rect 1428 -1412 1444 -1402
rect 522 -1454 1146 -1412
rect 400 -1460 1146 -1454
rect 1426 -1454 1444 -1412
rect 1496 -1454 1504 -1402
rect 1426 -1460 1504 -1454
rect 400 -1474 570 -1460
rect 1096 -1700 1144 -1460
rect 1434 -1498 1504 -1460
rect 1532 -1362 1600 -850
rect 1532 -1414 1542 -1362
rect 1594 -1414 1600 -1362
rect 1532 -1500 1600 -1414
rect 1633 -1406 1707 -1307
rect 3270 -1312 3408 -1300
rect 3270 -1388 3298 -1312
rect 3378 -1388 3408 -1312
rect 3270 -1402 3408 -1388
rect 1633 -1462 1640 -1406
rect 1692 -1462 1707 -1406
rect 1633 -1491 1707 -1462
rect 1633 -1565 1775 -1491
rect 1096 -1748 1606 -1700
rect 1558 -1920 1606 -1748
rect 792 -1926 1198 -1924
rect 722 -1936 1198 -1926
rect 722 -1988 730 -1936
rect 792 -1988 1198 -1936
rect 722 -1996 1198 -1988
rect 1126 -2122 1198 -1996
rect 1552 -1954 1650 -1920
rect 1552 -2006 1572 -1954
rect 1626 -2006 1650 -1954
rect 1552 -2024 1650 -2006
rect 1701 -2120 1775 -1565
rect 3290 -1636 3358 -1402
rect 3270 -1638 3358 -1636
rect 1572 -2122 1775 -2120
rect 1126 -2194 1775 -2122
rect 3210 -1706 3358 -1638
rect 1618 -2210 1690 -2194
rect 1618 -2264 1628 -2210
rect 1680 -2264 1690 -2210
rect 1618 -2348 1690 -2264
rect 392 -2902 542 -2888
rect 392 -2970 438 -2902
rect 500 -2954 542 -2902
rect 500 -2970 1622 -2954
rect 392 -2986 1622 -2970
rect 1590 -3166 1622 -2986
rect 3210 -3074 3278 -1706
rect 1766 -3084 3278 -3074
rect 1766 -3136 1772 -3084
rect 1824 -3136 3278 -3084
rect 1766 -3142 3278 -3136
rect 1574 -3174 1644 -3166
rect 1574 -3226 1582 -3174
rect 1634 -3226 1644 -3174
rect 1574 -3232 1644 -3226
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1754938408
transform 1 0 -2 0 1 6
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_1
timestamp 1754938408
transform 1 0 8 0 1 -1558
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_2
timestamp 1754938408
transform 1 0 10 0 1 -4790
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_3
timestamp 1754938408
transform 1 0 0 0 1 -3226
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_4
timestamp 1754938408
transform 1 0 1376 0 1 -3432
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_5
timestamp 1754938408
transform 1 0 1182 0 1 -604
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  sky130_fd_sc_hd__and3_1_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1754938408
transform 1 0 1380 0 1 -2412
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  sky130_fd_sc_hd__and4_1_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1754938408
transform 1 0 1256 0 1 -1570
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  sky130_fd_sc_hd__and4_1_1
timestamp 1754938408
transform 1 0 2040 0 1 -104
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  sky130_fd_sc_hd__or2_1_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1754938408
transform 1 0 2226 0 1 -1944
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  sky130_fd_sc_hd__or4_1_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1754938408
transform 1 0 3154 0 1 -1586
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1754938408
transform 1 0 -100 0 1 750
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_1
timestamp 1754938408
transform 1 0 -90 0 1 -814
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_2
timestamp 1754938408
transform 1 0 -88 0 1 -4046
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_3
timestamp 1754938408
transform 1 0 -98 0 1 -2482
box -38 -48 682 592
<< labels >>
rlabel metal1 s -90 -318 554 -222 1 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s -90 -862 554 -766 1 VGND
port 3 nsew ground bidirectional abutment
rlabel comment s -90 -814 -90 -814 4 xor2_1
flabel metal1 s -61 -831 -27 -797 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s -61 -287 -27 -253 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel nwell s -61 -287 -27 -253 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s -61 -831 -27 -797 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel locali s 123 -593 157 -559 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 491 -525 525 -491 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 31 -525 65 -491 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
rlabel metal1 s 8 -1062 468 -966 1 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 8 -1606 468 -1510 1 VGND
port 3 nsew ground bidirectional abutment
rlabel comment s 8 -1558 8 -1558 4 and2_1
flabel pwell s 37 -1575 71 -1541 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 37 -1031 71 -997 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel locali s 37 -1337 71 -1303 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 129 -1337 163 -1303 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 221 -1337 255 -1303 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 405 -1133 439 -1099 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 405 -1201 439 -1167 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 405 -1269 439 -1235 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 405 -1337 439 -1303 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 405 -1473 439 -1439 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 405 -1405 439 -1371 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel metal1 s 37 -1575 71 -1541 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 37 -1031 71 -997 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s -98 -1986 546 -1890 1 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s -98 -2530 546 -2434 1 VGND
port 3 nsew ground bidirectional abutment
rlabel comment s -98 -2482 -98 -2482 4 xor2_1
flabel metal1 s -69 -2499 -35 -2465 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s -69 -1955 -35 -1921 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel nwell s -69 -1955 -35 -1921 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s -69 -2499 -35 -2465 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel locali s 115 -2261 149 -2227 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 483 -2193 517 -2159 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 23 -2193 57 -2159 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
rlabel metal1 s 0 -2730 460 -2634 1 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 -3274 460 -3178 1 VGND
port 3 nsew ground bidirectional abutment
rlabel comment s 0 -3226 0 -3226 4 and2_1
flabel pwell s 29 -3243 63 -3209 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 29 -2699 63 -2665 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel locali s 29 -3005 63 -2971 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 121 -3005 155 -2971 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 213 -3005 247 -2971 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 397 -2801 431 -2767 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 397 -2869 431 -2835 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 397 -2937 431 -2903 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 397 -3005 431 -2971 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 397 -3141 431 -3107 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 397 -3073 431 -3039 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel metal1 s 29 -3243 63 -3209 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 29 -2699 63 -2665 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s -88 -3550 556 -3454 1 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s -88 -4094 556 -3998 1 VGND
port 3 nsew ground bidirectional abutment
rlabel comment s -88 -4046 -88 -4046 4 xor2_1
flabel metal1 s -59 -4063 -25 -4029 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s -59 -3519 -25 -3485 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel nwell s -59 -3519 -25 -3485 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s -59 -4063 -25 -4029 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel locali s 125 -3825 159 -3791 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 493 -3757 527 -3723 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 33 -3757 67 -3723 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
rlabel metal1 s 10 -4294 470 -4198 1 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 10 -4838 470 -4742 1 VGND
port 3 nsew ground bidirectional abutment
rlabel comment s 10 -4790 10 -4790 4 and2_1
flabel pwell s 39 -4807 73 -4773 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 39 -4263 73 -4229 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel locali s 39 -4569 73 -4535 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 131 -4569 165 -4535 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 223 -4569 257 -4535 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 407 -4365 441 -4331 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 407 -4433 441 -4399 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 407 -4501 441 -4467 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 407 -4569 441 -4535 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 407 -4705 441 -4671 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 407 -4637 441 -4603 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel metal1 s 39 -4807 73 -4773 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 39 -4263 73 -4229 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
<< end >>
