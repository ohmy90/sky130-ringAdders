* NGSPICE file created from tt_um_ohmy90_adders.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
.ends

.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X a_277_47#
X0 a_277_47# a_247_21# a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X1 VGND S0 a_247_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08138 pd=0.96719 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X2 a_834_97# a_247_21# a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=0.10858 pd=1.36 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=4318,272
X3 VGND A3 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0.08138 pd=0.96719 as=0.10855 ps=1.36 w=0.42 l=0.15
**devattr s=4316,272 d=2268,138
X4 a_1290_413# S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.08399 ps=0.95455 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X5 a_834_97# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10858 pd=1.36 as=0.08138 ps=0.96719 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X6 a_750_97# S0 a_757_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1274 pd=1.16667 as=0.10855 ps=1.36 w=0.42 l=0.15
**devattr s=4316,272 d=2268,138
X7 a_27_47# S0 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.09322 ps=1.07 w=0.42 l=0.15
**devattr s=3409,185 d=4368,272
X8 X a_1478_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12594 ps=1.49685 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X9 VPWR A1 a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.08399 pd=0.95455 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X10 VPWR S0 a_247_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.08399 pd=0.95455 as=0.1083 ps=1.36 w=0.42 l=0.15
**devattr s=4332,272 d=4316,272
X11 X a_1478_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.19997 ps=2.27273 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X12 a_193_47# A0 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.08138 ps=0.96719 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X13 a_750_97# a_1290_413# a_1478_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1274 pd=1.16667 as=0.09209 ps=0.99 w=0.42 l=0.15
**devattr s=3683,198 d=10752,424
X14 a_1478_413# S1 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09209 pd=0.99 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=3683,198
X15 a_1290_413# S1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.08138 ps=0.96719 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X16 a_277_47# a_247_21# a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.09322 pd=1.07 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3409,185
X17 a_750_97# S0 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.10855 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X18 a_923_363# a_247_21# a_750_97# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09013 pd=0.995 as=0.1274 ps=1.16667 w=0.42 l=0.15
**devattr s=2268,138 d=3605,199
X19 a_757_363# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.36 as=0.08399 ps=0.95455 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X20 VPWR A3 a_923_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.08399 pd=0.95455 as=0.09013 ps=0.995 w=0.42 l=0.15
**devattr s=3605,199 d=2268,138
X21 a_277_47# a_1290_413# a_1478_413# VNB sky130_fd_pr__nfet_01v8 ad=0.09322 pd=1.07 as=0.15102 ps=1.285 w=0.42 l=0.15
**devattr s=6041,257 d=4368,272
X22 a_193_413# A0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.36 as=0.08399 ps=0.95455 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X23 a_193_413# S0 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.36 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=4316,272
X24 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08138 pd=0.96719 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X25 a_1478_413# S1 a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=0.15102 pd=1.285 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=6041,257
.ends

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X a_117_297# a_285_297# a_285_47#
+ a_35_297#
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13813 ps=1.4 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.13813 pd=1.4 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.13813 pd=1.4 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13813 ps=1.4 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X a_145_75# a_59_75#
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.10288 pd=0.95413 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.24495 ps=2.27174 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.08777 pd=0.81645 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.10288 ps=0.95413 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.13583 ps=1.26355 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
.ends

.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X a_150_297# a_68_297#
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0873 pd=0.93866 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4010,197
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0873 ps=0.93866 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1351 ps=1.45268 w=0.65 l=0.15
**devattr s=4010,197 d=6760,364
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.08622 pd=0.78972 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5830,267
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.20528 ps=1.88028 w=1 l=0.15
**devattr s=5830,267 d=13600,536
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
.ends

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X a_109_47# a_197_47# a_303_47#
+ a_27_47#
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1394 ps=0.98731 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3319 ps=2.35075 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1394 ps=0.98731 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1394 pd=0.98731 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.15409 pd=1.04411 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1394 pd=0.98731 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.23846 ps=1.61589 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
.ends

.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X a_277_297# a_205_297# a_27_297#
+ a_109_297#
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.07685 ps=0.85082 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.07685 ps=0.85082 w=0.42 l=0.15
**devattr s=4368,272 d=2772,150
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0877 pd=0.79268 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=5930,268
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.11894 ps=1.31674 w=0.65 l=0.15
**devattr s=4075,198 d=7020,368
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.2088 ps=1.88732 w=1 l=0.15
**devattr s=5930,268 d=10800,508
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.07685 pd=0.85082 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2772,150 d=2268,138
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2772,150
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.07685 pd=0.85082 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2268,138 d=4075,198
.ends

.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X a_181_47# a_109_47# a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07394 pd=0.75265 as=0.0805 ps=0.94333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07394 pd=0.75265 as=0.0805 ps=0.94333 w=0.42 l=0.15
**devattr s=2646,147 d=5689,267
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=1764,126
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10335 pd=0.89495 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5266,228
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0805 pd=0.94333 as=0.07394 ps=0.75265 w=0.42 l=0.15
**devattr s=2268,138 d=2646,147
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.17604 ps=1.79204 w=1 l=0.15
**devattr s=5689,267 d=10400,504
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.15995 ps=1.38505 w=0.65 l=0.15
**devattr s=5266,228 d=6760,364
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
.ends

.subckt CLA VNB sky130_fd_sc_hd__and4_1_1/a_303_47# sky130_fd_sc_hd__and4_1_0/VPB
+ sky130_fd_sc_hd__xor2_1_0/VPB sky130_fd_sc_hd__and2_1_5/VPB a_n63_n2185# a_187_n2185#
+ sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__or4_1_0/D sky130_fd_sc_hd__or2_1_0/a_150_297#
+ a_n55_n517# sky130_fd_sc_hd__and2_1_5/a_59_75# sky130_fd_sc_hd__and4_1_1/VGND sky130_fd_sc_hd__and3_1_0/a_109_47#
+ sky130_fd_sc_hd__or4_1_0/VPWR sky130_fd_sc_hd__and3_1_0/a_181_47# sky130_fd_sc_hd__xor2_1_0/a_285_297#
+ sky130_fd_sc_hd__and2_1_0/B sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__or4_1_0/a_109_297#
+ sky130_fd_sc_hd__and2_1_4/VPWR sky130_fd_sc_hd__and2_1_0/A sky130_fd_sc_hd__or2_1_0/VPB
+ sky130_fd_sc_hd__and3_1_0/a_27_47# a_187_n2435# sky130_fd_sc_hd__and3_1_0/VPWR sky130_fd_sc_hd__and4_1_1/VPB
+ sky130_fd_sc_hd__xor2_1_0/a_285_47# a_19_n2185# sky130_fd_sc_hd__xor2_1_0/a_35_297#
+ sky130_fd_sc_hd__and2_1_4/a_145_75# sky130_fd_sc_hd__and2_1_0/a_145_75# sky130_fd_sc_hd__and4_1_1/a_27_47#
+ a_155_n4715# sky130_fd_sc_hd__or4_1_0/VGND sky130_fd_sc_hd__or4_1_0/A sky130_fd_sc_hd__and2_1_4/VGND
+ sky130_fd_sc_hd__or2_1_0/a_68_297# sky130_fd_sc_hd__and2_1_0/VPB a_195_n517# a_197_n3749#
+ sky130_fd_sc_hd__or4_1_0/X sky130_fd_sc_hd__and4_1_0/a_109_47# a_195_n767# a_197_n3999#
+ sky130_fd_sc_hd__and2_1_5/VPWR sky130_fd_sc_hd__and3_1_0/VGND sky130_fd_sc_hd__or2_1_0/VPWR
+ sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and2_1_5/a_145_75# sky130_fd_sc_hd__and2_1_0/a_59_75#
+ sky130_fd_sc_hd__and4_1_0/VPWR a_153_n1483# a_27_n517# a_69_n4715# sky130_fd_sc_hd__or2_1_0/B
+ sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__or4_1_0/a_277_297# sky130_fd_sc_hd__and4_1_0/a_197_47#
+ sky130_fd_sc_hd__and2_1_4/VPB sky130_fd_sc_hd__xor2_1_0/a_117_297# sky130_fd_sc_hd__and3_1_0/VPB
+ sky130_fd_sc_hd__and4_1_0/a_303_47# sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and4_1_1/a_109_47#
+ sky130_fd_sc_hd__or4_1_0/VPB sky130_fd_sc_hd__or4_1_0/a_27_297# a_29_n3749# sky130_fd_sc_hd__and2_1_5/VGND
+ sky130_fd_sc_hd__or4_1_0/a_205_297# sky130_fd_sc_hd__and2_1_4/a_59_75# sky130_fd_sc_hd__or2_1_0/VGND
+ a_n53_n3749# sky130_fd_sc_hd__and4_1_1/A sky130_fd_sc_hd__xor2_1_0/B sky130_fd_sc_hd__and4_1_0/VGND
+ sky130_fd_sc_hd__xor2_1_0/A sky130_fd_sc_hd__or4_1_0/C a_67_n1483# sky130_fd_sc_hd__and4_1_1/VPWR
+ a_59_n3151# sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and4_1_1/a_197_47# VPB
+ X B a_145_n3151# A
Xsky130_fd_sc_hd__xor2_1_3 A B A VNB VPB B X a_19_n2185# a_187_n2185# a_187_n2435#
+ a_n63_n2185# sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__and2_1_0 sky130_fd_sc_hd__and2_1_0/A sky130_fd_sc_hd__and2_1_0/B
+ sky130_fd_sc_hd__and2_1_0/A VNB sky130_fd_sc_hd__and2_1_0/VPB sky130_fd_sc_hd__and2_1_0/B
+ sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and2_1_0/a_145_75# sky130_fd_sc_hd__and2_1_0/a_59_75#
+ sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_1 A B A VNB VPB B X a_153_n1483# a_67_n1483# sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_3 A B A VNB VPB B X a_145_n3151# a_59_n3151# sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_2 A B A VNB VPB B X a_155_n4715# a_69_n4715# sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_4 X X sky130_fd_sc_hd__and2_1_4/VGND VNB sky130_fd_sc_hd__and2_1_4/VPB
+ sky130_fd_sc_hd__and2_1_4/VPWR sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__and2_1_4/a_145_75#
+ sky130_fd_sc_hd__and2_1_4/a_59_75# sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_5 X X sky130_fd_sc_hd__and2_1_5/VGND VNB sky130_fd_sc_hd__and2_1_5/VPB
+ sky130_fd_sc_hd__and2_1_5/VPWR sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and2_1_5/a_145_75#
+ sky130_fd_sc_hd__and2_1_5/a_59_75# sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__or2_1_0 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__or2_1_0/VGND
+ VNB sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__or2_1_0/VPWR sky130_fd_sc_hd__or4_1_0/A
+ sky130_fd_sc_hd__or2_1_0/a_150_297# sky130_fd_sc_hd__or2_1_0/a_68_297# sky130_fd_sc_hd__or2_1
Xsky130_fd_sc_hd__and4_1_0 X sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__xor2_1_0/X
+ X sky130_fd_sc_hd__and4_1_0/VGND VNB sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__and4_1_0/VPWR
+ sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__and4_1_0/a_109_47# sky130_fd_sc_hd__and4_1_0/a_197_47#
+ sky130_fd_sc_hd__and4_1_0/a_303_47# sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__and4_1
Xsky130_fd_sc_hd__and4_1_1 sky130_fd_sc_hd__and4_1_1/A X sky130_fd_sc_hd__and4_1_1/C
+ sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and4_1_1/VGND VNB sky130_fd_sc_hd__and4_1_1/VPB
+ sky130_fd_sc_hd__and4_1_1/VPWR sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__and4_1_1/a_109_47#
+ sky130_fd_sc_hd__and4_1_1/a_197_47# sky130_fd_sc_hd__and4_1_1/a_303_47# sky130_fd_sc_hd__and4_1_1/a_27_47#
+ sky130_fd_sc_hd__and4_1
Xsky130_fd_sc_hd__or4_1_0 sky130_fd_sc_hd__or4_1_0/A sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__or4_1_0/C
+ sky130_fd_sc_hd__or4_1_0/D sky130_fd_sc_hd__or4_1_0/VGND VNB sky130_fd_sc_hd__or4_1_0/VPB
+ sky130_fd_sc_hd__or4_1_0/VPWR sky130_fd_sc_hd__or4_1_0/X sky130_fd_sc_hd__or4_1_0/a_277_297#
+ sky130_fd_sc_hd__or4_1_0/a_205_297# sky130_fd_sc_hd__or4_1_0/a_27_297# sky130_fd_sc_hd__or4_1_0/a_109_297#
+ sky130_fd_sc_hd__or4_1
Xsky130_fd_sc_hd__and3_1_0 X X X sky130_fd_sc_hd__and3_1_0/VGND VNB sky130_fd_sc_hd__and3_1_0/VPB
+ sky130_fd_sc_hd__and3_1_0/VPWR sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__and3_1_0/a_181_47#
+ sky130_fd_sc_hd__and3_1_0/a_109_47# sky130_fd_sc_hd__and3_1_0/a_27_47# sky130_fd_sc_hd__and3_1
Xsky130_fd_sc_hd__xor2_1_0 sky130_fd_sc_hd__xor2_1_0/A sky130_fd_sc_hd__xor2_1_0/B
+ sky130_fd_sc_hd__xor2_1_0/A VNB sky130_fd_sc_hd__xor2_1_0/VPB sky130_fd_sc_hd__xor2_1_0/B
+ sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__xor2_1_0/a_117_297# sky130_fd_sc_hd__xor2_1_0/a_285_297#
+ sky130_fd_sc_hd__xor2_1_0/a_285_47# sky130_fd_sc_hd__xor2_1_0/a_35_297# sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_1 A B A VNB VPB B X a_27_n517# a_195_n517# a_195_n767# a_n55_n517#
+ sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_2 A B A VNB VPB B X a_29_n3749# a_197_n3749# a_197_n3999#
+ a_n53_n3749# sky130_fd_sc_hd__xor2_1
.ends

.subckt sky130_fd_sc_hd__fa_1 A B CIN VGND VNB VPB VPWR COUT SUM a_1163_413# a_738_413#
+ a_1163_47# a_208_47# a_382_413# a_738_47# a_995_47# a_1091_47# a_76_199# a_1091_413#
+ a_382_47# a_208_413#
X0 a_76_199# B a_208_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=2268,138
X1 VGND A a_382_47# VNB sky130_fd_pr__nfet_01v8 ad=0.07384 pd=0.80236 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X2 a_738_413# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.07885 ps=0.80769 w=0.42 l=0.15
**devattr s=2268,138 d=2478,143
X3 a_1091_47# CIN a_995_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X4 VPWR CIN a_738_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07885 pd=0.80769 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X5 a_382_413# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.07885 ps=0.80769 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X6 a_1163_47# B a_1091_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X7 VPWR A a_382_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07885 pd=0.80769 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X8 a_995_47# a_76_199# a_738_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2772,150
X9 a_382_413# CIN a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X10 SUM a_995_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11427 ps=1.24175 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X11 a_208_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.07384 ps=0.80236 w=0.42 l=0.15
**devattr s=4094,199 d=2520,144
X12 VGND CIN a_738_47# VNB sky130_fd_pr__nfet_01v8 ad=0.07384 pd=0.80236 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X13 a_76_199# B a_208_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=2268,138
X14 a_208_413# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.07885 ps=0.80769 w=0.42 l=0.15
**devattr s=5914,269 d=2520,144
X15 a_738_413# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.07885 ps=0.80769 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X16 VGND A a_1163_47# VNB sky130_fd_pr__nfet_01v8 ad=0.07384 pd=0.80236 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=4094,199
X17 a_738_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.07384 ps=0.80236 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X18 a_738_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.07384 ps=0.80236 w=0.42 l=0.15
**devattr s=2268,138 d=2478,143
X19 a_1163_413# B a_1091_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X20 VPWR A a_1163_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07885 pd=0.80769 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=5914,269
X21 a_382_47# CIN a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X22 a_382_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.07384 ps=0.80236 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X23 SUM a_995_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.18773 ps=1.92308 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X24 a_995_47# a_76_199# a_738_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2772,150
X25 VPWR a_76_199# COUT VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18773 pd=1.92308 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X26 a_1091_413# CIN a_995_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X27 VGND a_76_199# COUT VNB sky130_fd_pr__nfet_01v8 ad=0.11427 pd=1.24175 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
.ends

.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.08461 pd=0.79726 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.08461 ps=0.79726 w=0.42 l=0.15
**devattr s=2772,150 d=4704,280
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.08461 ps=0.79726 w=0.42 l=0.15
**devattr s=6334,279 d=3066,157
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11336 pd=0.94775 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=5796,222
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7728,268
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.11336 ps=0.94775 w=0.42 l=0.15
**devattr s=5796,222 d=4368,272
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
**devattr s=3990,179 d=2772,150
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
**devattr s=7728,268 d=1764,126
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=3990,179
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11336 ps=0.94775 w=0.42 l=0.15
**devattr s=4514,209 d=2772,150
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.20146 pd=1.89823 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=6334,279
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.17543 pd=1.46675 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4514,209
.ends

.subckt tt_um_ohmy90_adders clk ena rst_n ua[0] ua[1] ua[2] ua[3] VGND ua[5] ua[6]
+ ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0]
+ uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0]
+ uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0]
+ uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0]
+ uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
Xsky130_fd_sc_hd__inv_1_4 sky130_fd_sc_hd__inv_1_4/A VGND VNB sky130_fd_sc_hd__inv_1_4/VPB
+ VGND sky130_fd_sc_hd__inv_1_5/A sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_5 sky130_fd_sc_hd__inv_1_5/A VGND VNB sky130_fd_sc_hd__inv_1_5/VPB
+ VGND sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__mux4_1_0 sky130_fd_sc_hd__inv_1_5/Y VGND VGND VGND ui_in[1] ui_in[0]
+ VGND VNB sky130_fd_sc_hd__mux4_1_0/VPB VGND ua[0] ui_in[0] sky130_fd_sc_hd__mux4_1
XCLA_0 VNB CLA_0/sky130_fd_sc_hd__and4_1_1/a_303_47# CLA_0/sky130_fd_sc_hd__and4_1_0/VPB
+ CLA_0/sky130_fd_sc_hd__xor2_1_0/VPB CLA_0/sky130_fd_sc_hd__and2_1_5/VPB CLA_0/a_n63_n2185#
+ CLA_0/a_187_n2185# CLA_0/sky130_fd_sc_hd__and4_1_0/a_27_47# CLA_0/X CLA_0/sky130_fd_sc_hd__or2_1_0/a_150_297#
+ CLA_0/a_n55_n517# CLA_0/sky130_fd_sc_hd__and2_1_5/a_59_75# VGND CLA_0/sky130_fd_sc_hd__and3_1_0/a_109_47#
+ VGND CLA_0/sky130_fd_sc_hd__and3_1_0/a_181_47# CLA_0/sky130_fd_sc_hd__xor2_1_0/a_285_297#
+ VGND CLA_0/sky130_fd_sc_hd__or4_1_0/B CLA_0/sky130_fd_sc_hd__or4_1_0/a_109_297#
+ VGND VGND CLA_0/sky130_fd_sc_hd__or2_1_0/VPB CLA_0/sky130_fd_sc_hd__and3_1_0/a_27_47#
+ CLA_0/a_187_n2435# VGND CLA_0/sky130_fd_sc_hd__and4_1_1/VPB CLA_0/sky130_fd_sc_hd__xor2_1_0/a_285_47#
+ CLA_0/a_19_n2185# CLA_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# CLA_0/sky130_fd_sc_hd__and2_1_4/a_145_75#
+ CLA_0/sky130_fd_sc_hd__and2_1_0/a_145_75# CLA_0/sky130_fd_sc_hd__and4_1_1/a_27_47#
+ CLA_0/a_155_n4715# VGND CLA_0/sky130_fd_sc_hd__or4_1_0/A VGND CLA_0/sky130_fd_sc_hd__or2_1_0/a_68_297#
+ CLA_0/sky130_fd_sc_hd__and2_1_0/VPB CLA_0/a_195_n517# CLA_0/a_197_n3749# VGND CLA_0/sky130_fd_sc_hd__and4_1_0/a_109_47#
+ CLA_0/a_195_n767# CLA_0/a_197_n3999# VGND VGND VGND CLA_0/sky130_fd_sc_hd__and4_1_0/B
+ CLA_0/sky130_fd_sc_hd__and2_1_5/a_145_75# CLA_0/sky130_fd_sc_hd__and2_1_0/a_59_75#
+ VGND CLA_0/a_153_n1483# CLA_0/a_27_n517# CLA_0/a_69_n4715# CLA_0/sky130_fd_sc_hd__or2_1_0/B
+ CLA_0/sky130_fd_sc_hd__or2_1_0/A CLA_0/sky130_fd_sc_hd__or4_1_0/a_277_297# CLA_0/sky130_fd_sc_hd__and4_1_0/a_197_47#
+ CLA_0/sky130_fd_sc_hd__and2_1_4/VPB CLA_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# CLA_0/sky130_fd_sc_hd__and3_1_0/VPB
+ CLA_0/sky130_fd_sc_hd__and4_1_0/a_303_47# CLA_0/sky130_fd_sc_hd__and4_1_1/C CLA_0/sky130_fd_sc_hd__and4_1_1/a_109_47#
+ CLA_0/sky130_fd_sc_hd__or4_1_0/VPB CLA_0/sky130_fd_sc_hd__or4_1_0/a_27_297# CLA_0/a_29_n3749#
+ VGND CLA_0/sky130_fd_sc_hd__or4_1_0/a_205_297# CLA_0/sky130_fd_sc_hd__and2_1_4/a_59_75#
+ VGND CLA_0/a_n53_n3749# sky130_fd_sc_hd__inv_1_2/Y VGND VGND VGND CLA_0/sky130_fd_sc_hd__or4_1_0/C
+ CLA_0/a_67_n1483# VGND CLA_0/a_59_n3151# CLA_0/sky130_fd_sc_hd__xor2_1_0/X CLA_0/sky130_fd_sc_hd__and4_1_1/a_197_47#
+ CLA_0/VPB CLA_0/X VGND CLA_0/a_145_n3151# VGND CLA
XCLA_1 VNB a_11873_15219# VPB VPB VPB a_9959_13291# a_9717_13091# a_11321_14203# VGND
+ a_11906_13629# a_9967_14959# a_11019_15169# VGND a_11019_12911# VGND a_11091_12911#
+ a_9715_16323# VGND VGND a_12713_13987# VGND VGND VPB a_11261_13361# a_9717_12841#
+ VGND VPB a_9715_16073# a_9549_13091# a_9957_16523# a_11051_11919# a_9673_15357#
+ a_12105_15669# a_9685_10561# VGND VGND VGND a_12045_13829# VPB a_9725_14759# a_9727_11527#
+ VGND a_10895_13753# a_9725_14509# a_9727_11277# VGND VGND VGND VGND a_10857_14747#
+ a_9835_15779# VGND a_9683_13793# a_9557_14759# a_9847_10983# VGND VGND a_12881_13987#
+ a_10983_13753# VPB a_9547_16323# VPB a_11089_13753# VGND a_11679_15219# VPB a_13045_14187#
+ a_9559_11527# VGND a_12809_13987# a_11213_12341# VGND a_9969_11727# VGND VGND VGND
+ VGND VGND a_9845_14215# VGND a_9837_12547# VGND a_11767_15219# VPB VGND VGND a_9675_12125#
+ VGND CLA
Xsky130_fd_sc_hd__fa_1_10 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_2079_5051# a_2343_5051#
+ a_2079_5417# a_3040_5417# a_2706_5051# a_2343_5417# a_1950_5501# a_2175_5417# a_3199_5501#
+ a_2175_5051# a_2706_5417# a_3040_5051# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_0 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_2049_1791# a_2313_1791#
+ a_2049_2157# a_3010_2157# a_2676_1791# a_2313_2157# a_1920_2241# a_2145_2157# a_3169_2241#
+ a_2145_1791# a_2676_2157# a_3010_1791# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_11 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_3949_5047# a_4213_5047#
+ a_3949_5413# a_4910_5413# a_4576_5047# a_4213_5413# a_3820_5497# a_4045_5413# a_5069_5497#
+ a_4045_5047# a_4576_5413# a_4910_5047# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_1 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_3919_1787# a_4183_1787#
+ a_3919_2153# a_4880_2153# a_4546_1787# a_4183_2153# a_3790_2237# a_4015_2153# a_5039_2237#
+ a_4015_1787# a_4546_2153# a_4880_1787# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_12 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_11331_5467#
+ a_11595_5467# a_11331_5833# a_12292_5833# a_11958_5467# a_11595_5833# a_11202_5917#
+ a_11427_5833# a_12451_5917# a_11427_5467# a_11958_5833# a_12292_5467# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_3 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_7605_1779# a_7869_1779#
+ a_7605_2145# a_8566_2145# a_8232_1779# a_7869_2145# a_7476_2229# a_7701_2145# a_8725_2229#
+ a_7701_1779# a_8232_2145# a_8566_1779# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_2 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_5735_1783# a_5999_1783#
+ a_5735_2149# a_6696_2149# a_6362_1783# a_5999_2149# a_5606_2233# a_5831_2149# a_6855_2233#
+ a_5831_1783# a_6362_2149# a_6696_1783# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_4 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_14975_1765# a_15239_1765#
+ a_14975_2131# a_15936_2131# a_15602_1765# a_15239_2131# a_14846_2215# a_15071_2131#
+ a_16095_2215# a_15071_1765# a_15602_2131# a_15936_1765# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_13 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_9461_5471# a_9725_5471#
+ a_9461_5837# a_10422_5837# a_10088_5471# a_9725_5837# a_9332_5921# a_9557_5837#
+ a_9695_5921# a_9557_5471# a_10088_5837# a_10422_5471# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_15 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_15017_5459#
+ a_15281_5459# a_15017_5825# a_15978_5825# a_15644_5459# a_15281_5825# a_14888_5909#
+ a_15113_5825# a_16137_5909# a_15113_5459# a_15644_5825# a_15978_5459# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_14 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_13147_5463#
+ a_13411_5463# a_13147_5829# a_14108_5829# a_13774_5463# a_13411_5829# a_13018_5913#
+ a_13243_5829# a_14267_5913# a_13243_5463# a_13774_5829# a_14108_5463# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_5 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_13105_1769# a_13369_1769#
+ a_13105_2135# a_14066_2135# a_13732_1769# a_13369_2135# a_12976_2219# a_13201_2135#
+ a_14225_2219# a_13201_1769# a_13732_2135# a_14066_1769# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_16 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_11359_4593#
+ a_11623_4593# a_11359_4959# a_12320_4959# a_11986_4593# a_11623_4959# a_11230_5043#
+ a_11455_4959# a_12479_5043# a_11455_4593# a_11986_4959# a_12320_4593# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_6 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_9419_1777# a_9683_1777#
+ a_9419_2143# a_10380_2143# a_10046_1777# a_9683_2143# a_9290_2227# a_9515_2143#
+ a_9653_2227# a_9515_1777# a_10046_2143# a_10380_1777# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_7 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_11289_1773# a_11553_1773#
+ a_11289_2139# a_12250_2139# a_11916_1773# a_11553_2139# a_11160_2223# a_11385_2139#
+ a_12409_2223# a_11385_1773# a_11916_2139# a_12250_1773# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_17 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_9489_4597# a_9753_4597#
+ a_9489_4963# a_10450_4963# a_10116_4597# a_9753_4963# a_9360_5047# a_9585_4963#
+ a_9723_5047# a_9585_4597# a_10116_4963# a_10450_4597# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__mux2_1_0 VGND VGND VGND VGND VNB sky130_fd_sc_hd__mux2_1_0/VPB VGND
+ VGND sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__fa_1_18 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_13175_4589#
+ a_13439_4589# a_13175_4955# a_14136_4955# a_13802_4589# a_13439_4955# a_13046_5039#
+ a_13271_4955# a_14295_5039# a_13271_4589# a_13802_4955# a_14136_4589# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__inv_1_1 VGND VGND VNB VPB VGND VGND sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_0 VGND VGND VNB sky130_fd_sc_hd__inv_1_0/VPB VGND VGND sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__fa_1_8 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_7635_5039# a_7899_5039#
+ a_7635_5405# a_8596_5405# a_8262_5039# a_7899_5405# a_7506_5489# a_7731_5405# a_8755_5489#
+ a_7731_5039# a_8262_5405# a_8596_5039# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__inv_1_2 VGND VGND VNB sky130_fd_sc_hd__inv_1_2/VPB VGND sky130_fd_sc_hd__inv_1_2/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__fa_1_19 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_15045_4585#
+ a_15309_4585# a_15045_4951# a_16006_4951# a_15672_4585# a_15309_4951# a_14916_5035#
+ a_15141_4951# a_16165_5035# a_15141_4585# a_15672_4951# a_16006_4585# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_9 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_5765_5043# a_6029_5043#
+ a_5765_5409# a_6726_5409# a_6392_5043# a_6029_5409# a_5636_5493# a_5861_5409# a_6885_5493#
+ a_5861_5043# a_6392_5409# a_6726_5043# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__inv_1_3 sky130_fd_sc_hd__inv_1_5/Y VGND VNB sky130_fd_sc_hd__inv_1_3/VPB
+ VGND sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__inv_1
.ends

