* NGSPICE file created from tt_um_ohmy90_flat_adders.ext - technology: sky130A

.subckt tt_um_ohmy90_flat_adders clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5]
+ ua[6] ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7]
+ uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
+ uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
+ uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
+ VDPWR VGND
X0 a_4183_1787# a_4129_2043# a_3790_1761# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X1 a_15255_4841# a_14325_4589# a_15672_4585# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X2 a_24234_14385# ui_in[1] a_24152_14385# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.10855 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X3 VGND a_14888_5433# a_14836_5459# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X4 a_15113_5825# VDPWR a_15017_5825# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X5 a_13732_1769# VGND VDPWR w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X6 a_4711_15373# VGND a_4625_15373# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X7 a_11202_5441# a_10611_5471# a_11427_5467# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X8 VDPWR VGND a_2313_1791# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X9 VGND a_5636_5017# a_5584_5043# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X10 a_9865_15329# a_9587_15357# VDPWR w_9490_15543# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X11 a_1950_5025# a_2217_5025# a_2175_5051# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X12 VDPWR VDPWR a_15644_5459# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X13 a_5999_1783# a_5069_1787# VDPWR w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X14 VDPWR VDPWR a_9587_15357# w_9490_15543# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X15 a_4513_14775# VDPWR VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X16 a_6129_12927# a_4913_13781# a_6057_12927# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=1764,126
X17 VDPWR VDPWR a_6392_5043# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X18 a_11623_4959# a_11569_4849# a_11230_4567# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X19 VDPWR VDPWR a_11595_5467# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X20 sky130_fd_sc_hd__mux4_1_0.A3 a_17125_4938# VDPWR w_16764_4814# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=6334,279 d=10400,504
X21 a_13802_4955# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X22 a_7113_13395# a_6862_13645# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4010,197 d=6760,364
X23 VDPWR VGND a_15239_1765# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X24 a_3820_5021# a_3229_5051# a_4045_5413# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X25 VDPWR VGND a_4587_13107# w_4432_13071# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X26 a_13439_4955# a_12509_4593# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X27 a_15045_4951# a_14946_4905# a_14946_4905# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.07384 ps=0.80236 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X28 a_22274_16171# a_21506_16181# VDPWR w_22086_16385# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X29 a_2175_5417# VDPWR a_2079_5417# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X30 a_6089_11935# a_4849_11293# a_6003_11935# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X31 VDPWR VGND a_4597_11543# w_4442_11507# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X32 VDPWR a_9867_12097# a_10965_11919# w_10868_12105# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X33 a_14946_4905# a_14946_4905# a_15309_4951# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.07384 pd=0.80236 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X34 a_17346_5265# a_16195_4585# a_17125_4938# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
**devattr s=3990,179 d=2772,150
X35 VGND VGND a_9467_13091# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X36 a_15936_2131# VDPWR a_15185_2021# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X37 VGND VDPWR a_4213_5413# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X38 a_9671_5727# VGND a_10088_5471# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X39 a_11553_1773# a_11499_2029# a_11160_1747# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X40 a_13774_5463# VGND VDPWR w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X41 a_3949_5047# VGND VDPWR w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X42 VGND VGND a_8566_2145# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X43 a_9715_16323# VGND VDPWR w_9392_16287# sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X44 a_9725_14509# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X45 VGND a_1920_1765# a_1868_1791# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X46 VDPWR a_12075_13379# a_12881_13987# w_12566_13951# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=5930,268
X47 a_10422_5837# VDPWR a_9671_5727# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X48 VDPWR sky130_fd_sc_hd__mux4_1_0.A1 a_6629_15387# w_9392_17212# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X49 VDPWR VDPWR a_4753_16339# w_4430_16303# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X50 a_9332_5445# VGND a_9557_5837# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X51 VDPWR a_5606_1757# a_5554_1783# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X52 VDPWR a_12976_1743# a_12924_1769# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X53 a_4880_1787# VDPWR a_4129_2043# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X54 a_5945_2039# a_5069_1787# a_6362_2149# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X55 a_12509_4593# a_11569_4849# VDPWR w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X56 a_11359_4959# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X57 VGND VDPWR a_4546_2153# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X58 a_4903_15345# a_4625_15373# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X59 a_11541_5723# a_10611_5471# a_11958_5833# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X60 a_11230_4567# a_10639_4597# a_11455_4593# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X61 a_15644_5825# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X62 a_7476_1753# a_6885_1783# a_7701_2145# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X63 VDPWR VDPWR a_4763_14775# w_4440_14739# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X64 a_11291_12911# a_10937_12911# VDPWR w_10872_13125# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5689,267 d=10400,504
X65 a_8232_2145# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X66 a_7869_1779# a_7815_2035# a_7476_1753# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X67 a_5831_2149# VDPWR a_5735_2149# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X68 a_4913_13781# a_4635_13809# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X69 a_10813_13753# a_9799_16073# VDPWR w_10748_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X70 a_5735_1783# VGND VDPWR w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X71 VGND VDPWR a_9725_5837# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X72 VDPWR a_11202_5441# a_11150_5467# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X73 a_11499_2029# a_10569_1777# a_11916_2139# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X74 a_11986_4593# VGND VDPWR w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X75 VDPWR VDPWR a_9727_11527# w_9404_11491# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X76 a_9753_4597# VDPWR VDPWR w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X77 a_4723_10577# VGND a_4637_10577# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X78 VDPWR VDPWR a_11623_4593# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X79 a_4587_13107# VDPWR a_4505_13107# w_4432_13071# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X80 a_2079_5051# VGND VDPWR w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X81 VGND a_9360_4571# a_9308_4597# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X82 VDPWR VDPWR a_9599_10561# w_9502_10747# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X83 a_11331_5467# VGND VDPWR w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X84 a_4597_11543# VDPWR a_4515_11543# w_4442_11507# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X85 a_6944_13645# a_6329_12927# a_6862_13645# w_6756_13609# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X86 a_7669_14003# a_7173_15235# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X87 a_9467_13091# VDPWR VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X88 a_16195_4585# a_15255_4841# a_14946_4905# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11427 ps=1.24175 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X89 VDPWR VGND a_11595_5467# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X90 a_4635_13809# VGND VDPWR w_4538_13995# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X91 a_2706_5417# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X92 VDPWR VGND a_2343_5051# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X93 a_15281_5459# a_14297_5463# VDPWR w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X94 VGND a_4513_14775# a_4847_14525# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X95 a_5975_5299# a_5099_5047# a_6392_5409# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X96 VGND a_4503_16339# a_4837_16089# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X97 VGND a_9475_14759# a_9809_14509# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X98 a_13315_2025# a_12439_1773# a_13732_2135# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X99 VGND VDPWR a_4576_5413# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X100 VGND VGND a_10422_5837# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X101 a_6029_5043# a_5975_5299# a_5636_5017# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X102 a_12135_15219# a_11597_15219# VDPWR w_11532_15433# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X103 a_15602_2131# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X104 VDPWR VGND a_4880_1787# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X105 VGND a_8785_5039# a_16871_4938# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=5796,222
X106 a_11385_1773# VDPWR a_11289_1773# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X107 VGND sky130_fd_sc_hd__mux4_1_0.A1 a_23511_14335# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X108 VGND VGND a_4213_5413# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X109 VDPWR VGND a_14136_4589# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X110 VGND VGND a_15978_5825# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X111 a_6805_15235# a_4847_14525# a_6717_15235# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X112 a_7899_5405# a_6915_5043# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X113 VDPWR VDPWR a_13411_5463# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X114 a_15239_2131# a_14255_1769# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X115 a_9727_11527# VGND VDPWR w_9404_11491# sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X116 a_1920_1765# a_2187_1765# a_2145_2157# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X117 a_14325_4589# a_13385_4845# VDPWR w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X118 VDPWR a_11230_4567# a_11178_4593# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X119 VGND VDPWR a_9753_4963# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X120 a_16486_16197# sky130_fd_sc_hd__mux4_1_0.A0 VDPWR w_16298_16411# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X121 a_4546_1787# VGND VDPWR w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X122 a_23677_14701# ui_in[1] ui_in[0] sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.36 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=4316,272
X123 a_4905_12113# a_4627_12141# VDPWR w_4530_12327# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X124 a_4915_10549# a_4637_10577# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X125 a_9461_5837# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X126 a_14888_5433# a_14297_5463# a_15113_5825# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X127 a_7815_2035# a_6885_1783# a_8232_1779# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X128 a_7605_2145# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X129 VDPWR a_9809_14509# a_11597_15219# w_11532_15433# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X130 a_6087_14735# a_5809_14763# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X131 VGND a_6281_11907# a_7669_14003# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2772,150 d=2268,138
X132 VGND VDPWR a_2313_2157# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X133 VGND VDPWR a_11958_5833# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X134 a_13243_5829# VDPWR a_13147_5829# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X135 a_9683_2143# a_9629_2033# a_9290_1751# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X136 VGND VGND a_9725_5837# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X137 a_15672_4585# a_14946_4905# VDPWR w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X138 a_13411_5463# a_13357_5719# a_13018_5437# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X139 VDPWR VGND a_3010_1791# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X140 a_4183_2153# a_3199_1791# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X141 a_5099_5047# a_4159_5303# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X142 a_11553_2139# a_10569_1777# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X143 VDPWR VGND a_11623_4593# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X144 a_4763_14525# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X145 a_15309_4585# a_14325_4589# VDPWR w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X146 a_24962_14701# ui_in[0] a_24234_14385# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.15102 pd=1.285 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=6041,257
X147 a_4045_5047# VDPWR a_3949_5047# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X148 a_2259_2047# a_2187_1765# a_2676_1791# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X149 VDPWR VGND a_13369_1769# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X150 a_6696_1783# VDPWR a_5945_2039# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X151 VDPWR a_9290_1751# a_9238_1777# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X152 a_1950_5025# a_2217_5025# a_2175_5417# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X153 a_12631_13987# a_9877_10533# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4368,272 d=2772,150
X154 a_9589_12125# VGND VDPWR w_9492_12311# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X155 a_11906_13629# a_11291_12911# a_11824_13629# w_11718_13593# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X156 VGND VDPWR a_6392_5409# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X157 sky130_fd_sc_hd__mux4_1_0.A2 a_15185_2021# VDPWR w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X158 a_9753_4597# a_9699_4853# a_9360_4571# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X159 VDPWR a_13018_5437# a_12966_5463# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X160 VGND VDPWR a_13732_2135# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X161 a_6915_5043# a_5975_5299# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X162 a_7635_5405# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X163 a_12292_5467# VDPWR a_11541_5723# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X164 a_14946_4905# a_14946_4905# a_16006_4951# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.07384 pd=0.80236 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X165 a_14975_2131# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X166 a_15185_2021# a_14255_1769# a_15602_1765# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X167 VDPWR VGND a_9547_16323# w_9392_16287# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X168 a_3040_5051# VDPWR a_2289_5307# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X169 a_13201_1769# VDPWR a_13105_1769# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X170 a_8755_1779# a_7815_2035# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X171 a_5895_14763# a_4849_11293# a_5809_14763# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X172 VGND VGND a_9475_14759# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X173 VGND VGND a_7899_5405# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X174 VDPWR a_3790_1761# a_3738_1787# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X175 VGND VDPWR a_4711_15373# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X176 VDPWR a_9801_12841# a_10771_14747# w_10674_14933# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X177 a_5861_5043# VDPWR a_5765_5043# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X178 a_13147_5463# VGND VDPWR w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X179 VDPWR a_9799_16073# a_11597_15219# w_11532_15433# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X180 a_14916_4559# a_14325_4589# a_15141_4951# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X181 a_5069_1787# a_4129_2043# VDPWR w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X182 a_10639_4597# a_9699_4853# VDPWR w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X183 VGND VDPWR a_2676_2157# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X184 a_13271_4955# VDPWR a_13175_4955# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X185 VGND VGND a_4513_14775# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X186 a_9671_5727# VGND a_10088_5837# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X187 VDPWR a_14916_4559# a_14864_4585# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X188 a_11051_11919# a_9811_11277# a_10965_11919# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X189 a_13774_5829# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X190 a_3790_1761# a_3199_1791# a_4015_1787# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X191 VDPWR VDPWR a_13802_4589# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X192 VDPWR VDPWR a_8232_1779# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X193 a_11351_13753# a_10813_13753# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X194 VGND VGND a_2313_2157# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X195 VDPWR a_11351_13753# a_11906_13629# w_11718_13593# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5830,267
X196 a_9515_2143# VDPWR a_9419_2143# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X197 ua[0] a_24962_14701# VDPWR sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X198 a_4755_13107# VGND VDPWR w_4432_13071# sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X199 VDPWR VGND a_6696_1783# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X200 a_5999_2149# a_5069_1787# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X201 VDPWR VDPWR a_4183_1787# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X202 a_5933_13769# a_4849_11293# a_5851_13769# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
X203 a_9673_15357# VGND a_9587_15357# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X204 a_4576_5047# VGND VDPWR w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X205 VGND VGND a_15281_5825# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X206 VGND a_11160_1747# a_11108_1773# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X207 a_11230_4567# a_10639_4597# a_11455_4959# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X208 a_11597_15219# a_8113_13753# VDPWR w_11532_15433# sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X209 a_4765_11543# VGND VDPWR w_4442_11507# sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X210 a_21506_16181# a_20384_16179# VDPWR w_21318_16395# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X211 a_6885_1783# a_5945_2039# VDPWR w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X212 a_9683_13793# VGND a_9597_13793# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X213 VDPWR VGND a_12292_5467# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X214 a_9547_16323# VDPWR a_9465_16323# w_9392_16287# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X215 a_4503_16339# VDPWR VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X216 a_5606_1757# a_5069_1787# a_5831_1783# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X217 a_11986_4959# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X218 a_9475_14759# VDPWR VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X219 a_4015_2153# VDPWR a_3919_2153# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X220 a_17339_4938# a_16167_5459# a_17125_4938# w_16764_4814# sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
**devattr s=7728,268 d=3066,157
X221 VDPWR VGND a_3040_5051# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X222 a_11595_5833# a_11541_5723# a_11202_5441# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X223 a_6362_1783# VGND VDPWR w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X224 a_12320_4593# VDPWR a_11569_4849# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X225 VGND VDPWR a_11623_4959# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X226 VDPWR VDPWR a_9715_16323# w_9392_16287# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X227 a_10771_14747# a_9811_11277# VDPWR w_10674_14933# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X228 a_9809_14509# VDPWR a_9725_14509# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X229 a_2079_5417# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X230 a_3229_5051# a_2289_5307# VDPWR w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X231 a_9629_2033# a_8755_1779# a_10046_1777# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X232 VGND sky130_fd_sc_hd__mux4_1_0.A3 a_2217_5025# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X233 a_12481_5467# a_11541_5723# VDPWR w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X234 a_12439_1773# a_11499_2029# VDPWR w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X235 a_15309_4585# a_15255_4841# a_14916_4559# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X236 a_9585_4597# VDPWR a_9489_4597# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X237 a_11553_2139# a_11499_2029# a_11160_1747# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X238 a_11160_1747# a_10569_1777# a_11385_1773# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X239 a_14066_1769# VDPWR a_13315_2025# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X240 VGND a_7476_1753# a_7424_1779# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X241 a_2289_5307# a_2217_5025# a_2706_5051# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X242 a_15978_5459# VDPWR a_15227_5715# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X243 ui_in[0] a_23731_14309# a_23677_14335# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.09322 pd=1.07 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3409,185
X244 a_6389_13769# a_5851_13769# VDPWR w_5786_13983# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X245 a_11958_5467# VGND VDPWR w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X246 VDPWR a_4903_15345# a_5851_13769# w_5786_13983# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X247 VGND VGND a_2343_5417# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X248 VDPWR VDPWR a_15602_1765# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X249 a_7751_14003# a_4915_10549# a_7669_14003# w_7604_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2772,150
X250 VDPWR VGND a_9559_11527# w_9404_11491# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X251 a_16167_5459# a_15227_5715# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X252 VDPWR VDPWR a_2343_5051# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X253 a_9683_1777# a_8755_1779# VDPWR w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X254 a_9699_4853# VDPWR a_10116_4963# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X255 VGND VDPWR a_4723_10577# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X256 a_13369_2135# a_12439_1773# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X257 a_4625_15373# VGND VDPWR w_4528_15559# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X258 a_14136_4955# VDPWR a_13385_4845# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X259 a_19510_16177# a_18742_16187# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X260 a_11049_14719# a_10771_14747# VDPWR w_10674_14933# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X261 a_4159_5303# a_3229_5051# a_4576_5413# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X262 a_6029_5409# a_5975_5299# a_5636_5017# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X263 a_14946_4905# VDPWR a_15672_4951# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.07384 pd=0.80236 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X264 a_8596_5405# VDPWR a_7845_5295# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X265 a_5735_2149# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X266 a_24774_14701# ui_in[0] VDPWR sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X267 VDPWR a_3820_5021# a_3768_5047# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X268 a_18742_16187# a_18128_16189# VDPWR w_18554_16401# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X269 a_9865_15329# a_9587_15357# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X270 VDPWR VDPWR a_4635_13809# w_4538_13995# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X271 VGND VDPWR a_13411_5829# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X272 a_14108_5463# VDPWR a_13357_5719# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X273 a_9875_13765# a_9597_13793# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X274 a_10569_1777# a_9629_2033# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X275 VDPWR VGND a_4183_1787# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X276 a_17125_4938# a_16195_4585# a_17053_4938# w_16764_4814# sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=7728,268
X277 VDPWR VGND a_12320_4593# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X278 a_11291_12911# a_10937_12911# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=5266,228 d=6760,364
X279 VGND a_7506_5013# a_7454_5039# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X280 VDPWR sky130_fd_sc_hd__mux4_1_0.A1 a_23511_14701# sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X281 a_8113_13753# a_7669_14003# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4075,198 d=7020,368
X282 VGND a_14846_1739# a_14794_1765# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X283 a_15071_2131# VDPWR a_14975_2131# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X284 VDPWR sky130_fd_sc_hd__mux4_1_0.A2 a_2187_1765# w_6044_2758# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X285 VGND a_13046_4563# a_12994_4589# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X286 sky130_fd_sc_hd__mux4_1_0.A0 a_22274_16171# VDPWR w_22960_16387# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X287 ui_in[0] a_24774_14701# a_24962_14701# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.09322 pd=1.07 as=0.15102 ps=1.285 w=0.42 l=0.15
**devattr s=6041,257 d=4368,272
X288 a_6057_12927# a_4849_11293# a_5975_12927# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X289 a_9725_5471# VGND VDPWR w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X290 a_7869_1779# a_6885_1783# VDPWR w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X291 a_3199_1791# a_2259_2047# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X292 VDPWR VDPWR a_8262_5039# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X293 a_23677_14335# sky130_fd_sc_hd__mux4_1_0.A0 VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X294 VDPWR VGND a_14066_1769# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X295 a_13411_5829# a_13357_5719# a_13018_5437# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X296 VGND a_6389_13769# a_6862_13645# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4010,197
X297 a_9559_11527# VDPWR a_9477_11527# w_9404_11491# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X298 a_11427_5833# VDPWR a_11331_5833# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X299 a_16006_4585# VDPWR a_15255_4841# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X300 VGND VGND a_11623_4959# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X301 a_7919_14003# a_7173_15235# a_7847_14003# w_7604_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X302 a_14255_1769# a_13315_2025# VDPWR w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X303 a_11243_11891# a_10965_11919# VDPWR w_10868_12105# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X304 VDPWR VDPWR a_10046_1777# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X305 a_12976_1743# a_12439_1773# a_13201_1769# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X306 a_2313_1791# a_2187_1765# VDPWR w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X307 a_5975_12927# a_4913_13781# VDPWR w_5910_13141# sky130_fd_pr__pfet_01v8_hvt ad=0.0805 pd=0.94333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2646,147
X308 a_11385_2139# VDPWR a_11289_2139# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X309 VDPWR VDPWR a_2706_5051# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X310 a_11289_1773# VGND VDPWR w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X311 a_4213_5047# a_4159_5303# a_3820_5021# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X312 a_5636_5017# a_5099_5047# a_5861_5043# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X313 VDPWR VDPWR a_5999_1783# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X314 VDPWR VDPWR a_13369_1769# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X315 a_15141_4585# VDPWR a_15045_4585# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X316 VGND VGND a_8596_5405# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X317 a_6392_5043# VGND VDPWR w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X318 VGND a_4837_16089# a_6911_15235# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X319 VGND VGND a_15936_2131# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X320 VGND VDPWR a_10116_4963# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X321 a_13046_4563# a_12509_4593# a_13271_4955# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X322 VDPWR VGND a_11553_1773# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X323 VDPWR VGND a_14108_5463# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X324 a_4847_14525# VDPWR a_4763_14525# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X325 a_6029_5043# a_5099_5047# VDPWR w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X326 VGND VDPWR a_13439_4955# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X327 a_3040_5417# VDPWR a_2289_5307# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X328 a_7506_5013# a_6915_5043# a_7731_5405# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X329 a_8262_5405# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X330 a_10380_2143# VDPWR a_9629_2033# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X331 a_13147_5829# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X332 a_9290_1751# a_8755_1779# a_9515_2143# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X333 a_4713_12141# VGND a_4627_12141# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X334 a_5861_5409# VDPWR a_5765_5409# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X335 a_14297_5463# a_13357_5719# VDPWR w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X336 a_10983_13753# a_9865_15329# a_10895_13753# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X337 a_11089_13753# a_9799_16073# a_10983_13753# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X338 a_13018_5437# a_12481_5467# a_13243_5463# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X339 a_13369_2135# a_13315_2025# a_12976_1743# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X340 VGND VGND a_3010_2157# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X341 a_9867_12097# a_9589_12125# VDPWR w_9492_12311# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X342 a_6717_15235# a_6629_15387# a_6635_15235# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
X343 a_4837_16089# a_4503_16339# a_4753_16339# w_4430_16303# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X344 VDPWR VDPWR a_9589_12125# w_9492_12311# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X345 VDPWR VDPWR a_10088_5471# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X346 a_9877_10533# a_9599_10561# VDPWR w_9502_10747# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X347 VDPWR VGND a_7869_1779# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X348 VGND VDPWR a_9683_2143# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X349 a_2259_2047# a_2187_1765# a_2676_2157# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X350 a_4753_16089# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X351 VDPWR a_4849_11293# a_5975_12927# w_5910_13141# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0805 ps=0.94333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X352 VGND a_4839_12857# a_5895_14763# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X353 a_6696_2149# VDPWR a_5945_2039# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X354 a_15227_5715# a_14297_5463# a_15644_5825# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X355 a_10450_4597# VDPWR a_9699_4853# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X356 VDPWR a_14888_5433# a_14836_5459# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X357 a_9360_4571# VDPWR a_9585_4597# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X358 a_18128_16189# a_17254_16187# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X359 VDPWR a_5636_5017# a_5584_5043# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X360 a_7701_1779# VDPWR a_7605_1779# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X361 a_12135_15219# a_11597_15219# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X362 a_4910_5047# VDPWR a_4159_5303# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X363 a_13439_4589# a_13385_4845# a_13046_4563# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X364 a_11569_4849# a_10639_4597# a_11986_4593# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X365 VGND a_9867_12097# a_11051_11919# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X366 a_13105_1769# VGND VDPWR w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X367 VGND VDPWR a_7869_2145# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X368 a_17125_4938# a_16167_5459# a_17125_5265# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=3990,179
X369 a_15017_5459# VGND VDPWR w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X370 VGND sky130_fd_sc_hd__mux4_1_0.A1 a_6629_15387# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X371 VGND VGND a_3040_5417# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X372 VDPWR VGND a_5999_1783# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X373 a_7899_5039# a_7845_5295# a_7506_5013# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X374 a_11873_15219# a_11049_14719# a_11767_15219# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X375 VDPWR a_9801_12841# a_10813_13753# w_10748_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X376 a_5765_5043# VGND VDPWR w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X377 a_12509_4593# a_11569_4849# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X378 a_12320_4959# VDPWR a_11569_4849# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X379 VGND VGND a_10380_2143# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X380 VGND a_4505_13107# a_4839_12857# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X381 VDPWR VDPWR a_4755_13107# w_4432_13071# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X382 sky130_fd_sc_hd__mux4_1_0.A3 a_17125_4938# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4514,209 d=6760,364
X383 a_10937_12911# a_9875_13765# VDPWR w_10872_13125# sky130_fd_pr__pfet_01v8_hvt ad=0.0805 pd=0.94333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2646,147
X384 a_11595_5467# a_10611_5471# VDPWR w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X385 a_13175_4955# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X386 a_4905_12113# a_4627_12141# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X387 a_2289_5307# a_2217_5025# a_2706_5417# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X388 VDPWR VDPWR a_15281_5459# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X389 VGND VDPWR a_9673_15357# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X390 VDPWR sky130_fd_sc_hd__mux4_1_0.A3 a_24407_14651# sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.09013 ps=0.995 w=0.42 l=0.15
**devattr s=3605,199 d=2268,138
X391 VDPWR VDPWR a_4765_11543# w_4442_11507# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X392 VDPWR a_7113_13395# a_7919_14003# w_7604_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=5930,268
X393 VGND VGND a_13439_4955# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X394 VGND VDPWR a_9683_13793# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X395 a_10046_2143# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X396 VGND VGND a_4503_16339# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X397 VGND VDPWR a_2343_5417# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X398 a_9419_2143# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X399 a_12075_13379# a_11824_13629# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4010,197 d=6760,364
X400 VGND VGND a_6696_2149# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X401 sky130_fd_sc_hd__mux4_1_0.A1 a_12631_13987# VDPWR w_12566_13951# sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5930,268 d=10800,508
X402 a_12250_1773# VDPWR a_11499_2029# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X403 a_4213_5413# a_3229_5051# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X404 a_14846_1739# a_14255_1769# a_15071_2131# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X405 VDPWR VGND a_10450_4597# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X406 VDPWR VDPWR a_13774_5463# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X407 a_15239_1765# a_15185_2021# a_14846_1739# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X408 a_15281_5459# a_15227_5715# a_14888_5433# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X409 a_20384_16179# a_19510_16177# VDPWR w_20196_16393# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X410 VGND VDPWR a_7899_5405# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X411 VGND VDPWR a_15239_2131# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X412 VGND VGND a_9683_2143# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X413 a_15255_4841# a_14325_4589# a_15672_4951# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X414 a_17254_16187# a_16486_16197# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X415 a_6862_13645# a_6329_12927# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X416 VDPWR VGND a_4910_5047# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X417 VDPWR VGND a_13411_5463# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X418 a_5606_1757# a_5069_1787# a_5831_2149# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X419 a_11202_5441# a_10611_5471# a_11427_5833# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X420 a_14108_5829# VDPWR a_13357_5719# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X421 a_6362_2149# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X422 VGND a_5606_1757# a_5554_1783# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X423 a_3919_2153# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X424 a_4129_2043# a_3199_1791# a_4546_1787# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X425 a_5851_13769# a_4849_11293# VDPWR w_5786_13983# sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X426 a_4721_13809# VGND a_4635_13809# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X427 VDPWR a_9865_15329# a_10813_13753# w_10748_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X428 VDPWR a_4847_14525# a_6635_15235# w_6570_15449# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X429 VGND VDPWR a_15644_5825# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X430 a_8566_1779# VDPWR a_7815_2035# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X431 a_10116_4597# VGND VDPWR w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X432 VGND VGND a_12320_4959# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X433 VGND a_9801_12841# a_11089_13753# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X434 a_9489_4597# VGND VDPWR w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X435 VDPWR VDPWR a_4625_15373# w_4528_15559# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X436 a_12631_13987# a_12135_15219# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X437 a_9725_5837# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X438 a_11160_1747# a_10569_1777# a_11385_2139# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X439 a_13385_4845# a_12509_4593# a_13802_4589# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X440 VGND VDPWR a_11595_5833# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X441 VDPWR VDPWR a_11986_4593# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X442 a_7113_13395# a_6862_13645# VDPWR w_6756_13609# sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5830,267 d=13600,536
X443 a_11091_12911# a_9875_13765# a_11019_12911# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=1764,126
X444 a_8785_5039# a_7845_5295# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X445 a_11623_4593# a_10639_4597# VDPWR w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X446 a_7845_5295# a_6915_5043# a_8262_5039# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X447 a_14325_4589# a_13385_4845# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X448 a_9557_5471# VDPWR a_9461_5471# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X449 VDPWR VDPWR a_15309_4585# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X450 VDPWR VGND a_9753_4597# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X451 VDPWR a_8785_5039# a_17339_4938# w_16764_4814# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=6334,279
X452 VGND a_11230_4567# a_11178_4593# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X453 a_7731_5039# VDPWR a_7635_5039# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X454 a_24774_14701# ui_in[0] VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X455 VDPWR VGND a_12250_1773# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X456 a_23677_14701# sky130_fd_sc_hd__mux4_1_0.A0 VDPWR sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.36 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X457 VGND VGND a_4505_13107# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X458 VGND VDPWR a_2706_5417# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X459 a_5636_5017# a_5099_5047# a_5861_5409# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X460 a_4183_2153# a_4129_2043# a_3790_1761# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X461 a_3949_5413# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X462 a_6392_5409# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X463 ua[0] a_24962_14701# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X464 a_9801_12841# a_9467_13091# a_9717_13091# w_9394_13055# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X465 a_13732_2135# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X466 a_2145_1791# VDPWR a_2049_1791# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X467 a_6726_5043# VDPWR a_5975_5299# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X468 a_15936_1765# VDPWR a_15185_2021# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X469 a_5809_14763# a_4849_11293# VDPWR w_5712_14949# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X470 a_6029_5409# a_5099_5047# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X471 VGND VGND a_14108_5829# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X472 a_11916_1773# VGND VDPWR w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X473 VGND a_9801_12841# a_11091_12911# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5266,228
X474 VDPWR VDPWR a_11553_1773# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X475 VDPWR VGND a_8566_1779# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X476 a_15113_5459# VDPWR a_15017_5459# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X477 VGND a_11243_11891# a_12631_13987# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2772,150 d=2268,138
X478 VDPWR a_4837_16089# a_6635_15235# w_6570_15449# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X479 VGND VGND a_15239_2131# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X480 a_13018_5437# a_12481_5467# a_13243_5829# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X481 a_8755_1779# a_7815_2035# VDPWR w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X482 a_9753_4963# VDPWR VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X483 VDPWR VDPWR a_4546_1787# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X484 VGND VDPWR a_10088_5837# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X485 a_7476_1753# a_6885_1783# a_7701_1779# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X486 a_13802_4589# VGND VDPWR w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X487 a_12713_13987# a_9877_10533# a_12631_13987# w_12566_13951# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2772,150
X488 a_8232_1779# VGND VDPWR w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X489 a_10611_5471# a_9671_5727# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X490 a_11331_5833# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X491 a_2313_2157# a_2187_1765# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X492 a_11767_15219# a_9809_14509# a_11679_15219# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X493 a_11824_13629# a_11291_12911# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X494 a_5099_5047# a_4159_5303# VDPWR w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X495 a_11289_2139# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X496 VGND a_9332_5445# a_9280_5471# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X497 a_3820_5021# a_3229_5051# a_4045_5047# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X498 VGND VDPWR a_5999_2149# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X499 a_22274_16171# a_21506_16181# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X500 a_10813_13753# a_9811_11277# VDPWR w_10748_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X501 a_4505_13107# VDPWR VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X502 VGND VGND a_11595_5833# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X503 a_13439_4589# a_12509_4593# VDPWR w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X504 a_15045_4585# a_14946_4905# VDPWR w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X505 a_6635_15235# a_6629_15387# VDPWR w_6570_15449# sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X506 VGND VDPWR a_4713_12141# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X507 a_15281_5825# a_14297_5463# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X508 VGND VGND a_4515_11543# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X509 a_10639_4597# a_9699_4853# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X510 VGND a_9801_12841# a_10857_14747# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X511 VDPWR a_14946_4905# a_15309_4585# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X512 a_14946_4905# a_14916_4559# a_14864_4585# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.11427 pd=1.24175 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X513 a_11049_14719# a_10771_14747# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X514 a_9597_13793# VGND VDPWR w_9500_13979# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X515 VGND VGND a_11553_2139# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X516 VDPWR VDPWR a_4213_5047# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X517 VDPWR VGND a_6726_5043# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X518 a_4880_2153# VDPWR a_4129_2043# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X519 a_11569_4849# a_10639_4597# a_11986_4959# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X520 a_9715_16073# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X521 a_2676_1791# VGND VDPWR w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X522 VDPWR a_11160_1747# a_11108_1773# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X523 a_7869_2145# a_7815_2035# a_7476_1753# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X524 a_5765_5409# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X525 VGND VGND a_14136_4955# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X526 a_4837_16089# VDPWR a_4753_16089# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X527 a_6915_5043# a_5975_5299# VDPWR w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X528 a_4913_13781# a_4635_13809# VDPWR w_4538_13995# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X529 VDPWR a_4839_12857# a_5975_12927# w_5910_13141# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0805 ps=0.94333 w=0.42 l=0.15
**devattr s=2646,147 d=5689,267
X530 a_6329_12927# a_5975_12927# VDPWR w_5910_13141# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5689,267 d=10400,504
X531 VGND a_1950_5025# a_1898_5051# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X532 a_13315_2025# a_12439_1773# a_13732_1769# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X533 VDPWR a_9811_11277# a_10937_12911# w_10872_13125# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0805 ps=0.94333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X534 VDPWR VDPWR a_11916_1773# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X535 a_11541_5723# a_10611_5471# a_11958_5467# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X536 a_15644_5459# VGND VDPWR w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X537 a_9675_12125# VGND a_9589_12125# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X538 a_15602_1765# VGND VDPWR w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X539 a_11597_15219# a_11049_14719# VDPWR w_11532_15433# sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X540 a_24234_14385# ui_in[1] a_24241_14651# sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1274 pd=1.16667 as=0.10855 ps=1.36 w=0.42 l=0.15
**devattr s=4316,272 d=2268,138
X541 VDPWR VDPWR a_9717_13091# w_9394_13055# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X542 a_6281_11907# a_6003_11935# VDPWR w_5906_12121# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X543 a_9811_11277# VDPWR a_9727_11277# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X544 VGND a_3790_1761# a_3738_1787# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X545 VDPWR a_4905_12113# a_6003_11935# w_5906_12121# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X546 a_9685_10561# VGND a_9599_10561# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X547 a_15239_1765# a_14255_1769# VDPWR w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X548 VDPWR a_7476_1753# a_7424_1779# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X549 a_4847_14525# a_4513_14775# a_4763_14775# w_4440_14739# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X550 a_5069_1787# a_4129_2043# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X551 a_15672_4951# a_14946_4905# a_14946_4905# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.07384 ps=0.80236 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X552 a_9809_14509# a_9475_14759# a_9725_14759# w_9402_14723# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X553 a_10895_13753# a_9811_11277# a_10813_13753# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
X554 a_4515_11543# VDPWR VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X555 VGND VDPWR a_13774_5829# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X556 a_10857_14747# a_9811_11277# a_10771_14747# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X557 a_7605_1779# VGND VDPWR w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X558 a_7847_14003# a_6281_11907# a_7751_14003# w_7604_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X559 a_15309_4951# a_14325_4589# a_14946_4905# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.07384 ps=0.80236 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X560 a_13357_5719# a_12481_5467# a_13774_5463# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X561 a_9683_1777# a_9629_2033# a_9290_1751# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X562 a_17125_5265# a_16871_4938# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=5796,222 d=2772,150
X563 a_24241_14651# sky130_fd_sc_hd__mux4_1_0.A2 VDPWR sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.36 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X564 a_4045_5413# VDPWR a_3949_5413# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X565 VGND VGND a_13411_5829# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X566 VGND VGND a_4880_2153# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X567 VGND a_9465_16323# a_9799_16073# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X568 VGND VGND a_5999_2149# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X569 a_4183_1787# a_3199_1791# VDPWR w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X570 VDPWR VDPWR a_4576_5047# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X571 a_6021_13769# a_4903_15345# a_5933_13769# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X572 VDPWR a_1920_1765# a_1868_1791# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X573 VGND sky130_fd_sc_hd__mux4_1_0.A3 a_24152_14385# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.10855 ps=1.36 w=0.42 l=0.15
**devattr s=4316,272 d=2268,138
X574 a_6127_13769# a_4837_16089# a_6021_13769# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X575 a_4627_12141# VGND VDPWR w_4530_12327# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X576 a_6885_1783# a_5945_2039# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X577 a_9753_4963# a_9699_4853# a_9360_4571# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X578 VDPWR VGND a_4213_5047# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X579 a_12292_5833# VDPWR a_11541_5723# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X580 a_4546_2153# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X581 VGND VDPWR a_11986_4959# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X582 a_4637_10577# VGND VDPWR w_4540_10763# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X583 VDPWR sky130_fd_sc_hd__mux4_1_0.A3 a_2217_5025# w_6074_6018# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X584 a_10569_1777# a_9629_2033# VDPWR w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X585 a_11623_4959# a_10639_4597# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X586 VDPWR VGND a_15978_5459# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X587 a_9717_13091# VGND VDPWR w_9394_13055# sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X588 a_9727_11277# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X589 a_7815_2035# a_6885_1783# a_8232_2145# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X590 a_7899_5039# a_6915_5043# VDPWR w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X591 VGND ui_in[1] a_23731_14309# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X592 VDPWR a_14846_1739# a_14794_1765# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X593 a_6003_11935# a_4849_11293# VDPWR w_5906_12121# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X594 a_9557_5837# VDPWR a_9461_5837# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X595 VDPWR VDPWR a_6362_1783# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X596 a_12250_2139# VDPWR a_11499_2029# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X597 VDPWR VDPWR a_13732_1769# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X598 a_16486_16197# sky130_fd_sc_hd__mux4_1_0.A0 VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X599 VGND VDPWR a_4721_13809# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X600 a_9725_5471# a_9671_5727# a_9332_5445# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X601 VDPWR VDPWR a_9753_4597# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X602 a_11455_4593# VDPWR a_11359_4593# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X603 a_16167_5459# a_15227_5715# VDPWR w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X604 a_9877_10533# a_9599_10561# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X605 VGND a_11202_5441# a_11150_5467# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X606 a_14975_1765# VGND VDPWR w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X607 a_14888_5433# a_14297_5463# a_15113_5459# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X608 VGND a_12075_13379# a_12631_13987# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2268,138 d=4075,198
X609 VDPWR a_9801_12841# a_10937_12911# w_10872_13125# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0805 ps=0.94333 w=0.42 l=0.15
**devattr s=2646,147 d=5689,267
X610 VDPWR VDPWR a_11958_5467# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X611 a_2343_5051# a_2217_5025# VDPWR w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X612 VGND VGND a_13369_2135# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X613 VGND VDPWR a_13802_4955# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X614 a_7173_15235# a_6635_15235# VDPWR w_6570_15449# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X615 a_24234_14385# a_24774_14701# a_24962_14701# sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1274 pd=1.16667 as=0.09209 ps=0.99 w=0.42 l=0.15
**devattr s=3683,198 d=10752,424
X616 a_6726_5409# VDPWR a_5975_5299# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X617 VDPWR VDPWR a_6029_5043# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X618 a_2313_1791# a_2259_2047# a_1920_1765# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X619 a_12881_13987# a_12135_15219# a_12809_13987# w_12566_13951# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X620 a_4576_5413# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X621 a_4755_12857# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X622 VGND a_4515_11543# a_4849_11293# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X623 VDPWR a_7506_5013# a_7454_5039# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X624 a_9515_1777# VDPWR a_9419_1777# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X625 VGND a_12976_1743# a_12924_1769# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X626 a_13201_2135# VDPWR a_13105_2135# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X627 a_15185_2021# a_14255_1769# a_15602_2131# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X628 VGND VGND a_12292_5833# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X629 a_10088_5471# VGND VDPWR w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X630 a_4585_16339# VDPWR a_4503_16339# w_4430_16303# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X631 VGND a_9477_11527# a_9811_11277# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X632 VDPWR a_14946_4905# a_16006_4585# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X633 VDPWR a_4839_12857# a_5809_14763# w_5712_14949# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X634 a_7635_5039# VGND VDPWR w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X635 VGND VGND a_9465_16323# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X636 a_4595_14775# VDPWR a_4513_14775# w_4440_14739# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X637 VGND VGND a_12250_2139# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X638 VDPWR a_9360_4571# a_9308_4597# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X639 a_15309_4951# a_15255_4841# a_14916_4559# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X640 a_9585_4963# VDPWR a_9489_4963# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X641 VDPWR VGND a_7899_5039# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X642 a_15978_5825# VDPWR a_15227_5715# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X643 a_3790_1761# a_3199_1791# a_4015_2153# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X644 a_11958_5833# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X645 a_4015_1787# VDPWR a_3919_1787# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X646 a_16195_4585# a_15255_4841# VDPWR w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X647 VGND VDPWR a_8232_2145# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X648 a_2049_1791# VGND VDPWR w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X649 a_2145_2157# VDPWR a_2049_2157# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X650 a_14916_4559# a_14325_4589# a_15141_4585# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X651 sky130_fd_sc_hd__mux4_1_0.A1 a_12631_13987# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4075,198 d=7020,368
X652 a_11351_13753# a_10813_13753# VDPWR w_10748_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X653 a_11916_2139# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X654 a_13271_4589# VDPWR a_13175_4589# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X655 a_6389_13769# a_5851_13769# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X656 a_4839_12857# a_4505_13107# a_4755_13107# w_4432_13071# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X657 VGND VGND a_6726_5409# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X658 VGND VDPWR a_4183_2153# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X659 VGND VDPWR a_11553_2139# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X660 a_19510_16177# a_18742_16187# VDPWR w_19322_16391# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X661 VGND a_4839_12857# a_6127_13769# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X662 VGND a_11351_13753# a_11824_13629# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4010,197
X663 a_3010_1791# VDPWR a_2259_2047# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X664 a_13369_1769# a_12439_1773# VDPWR w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X665 a_23511_14335# ui_in[1] ui_in[0] sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.09322 ps=1.07 w=0.42 l=0.15
**devattr s=3409,185 d=4368,272
X666 a_9725_14759# VGND VDPWR w_9402_14723# sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X667 a_4765_11293# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X668 VDPWR VGND a_6029_5043# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X669 a_5999_1783# a_5945_2039# a_5606_1757# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X670 VDPWR VGND a_15281_5459# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X671 a_21506_16181# a_20384_16179# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X672 VDPWR VDPWR a_9597_13793# w_9500_13979# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X673 a_4903_15345# a_4625_15373# VDPWR w_4528_15559# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X674 a_9629_2033# a_8755_1779# a_10046_2143# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X675 VGND a_9799_16073# a_11873_15219# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X676 a_9465_16323# VDPWR VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X677 a_14066_2135# VDPWR a_13315_2025# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X678 a_9799_16073# VDPWR a_9715_16073# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X679 VGND VDPWR a_8262_5405# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X680 a_11595_5467# a_11541_5723# a_11202_5441# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X681 VGND a_13018_5437# a_12966_5463# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X682 VGND VDPWR a_15602_2131# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X683 a_2343_5051# a_2289_5307# a_1950_5025# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X684 a_7669_14003# a_4915_10549# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4368,272 d=2772,150
X685 a_15071_1765# VDPWR a_14975_1765# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X686 a_9683_2143# a_8755_1779# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X687 a_16006_4951# VDPWR a_15255_4841# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X688 VDPWR a_6389_13769# a_6944_13645# w_6756_13609# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5830,267
X689 VDPWR a_8785_5039# a_16871_4938# w_16764_4814# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2772,150
X690 a_13411_5463# a_12481_5467# VDPWR w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X691 a_13357_5719# a_12481_5467# a_13774_5829# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X692 VDPWR VGND a_9549_13091# w_9394_13055# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X693 VGND VDPWR a_9675_12125# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X694 VGND VGND a_9477_11527# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X695 a_24407_14651# a_23731_14309# a_24234_14385# sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09013 pd=0.995 as=0.1274 ps=1.16667 w=0.42 l=0.15
**devattr s=2268,138 d=3605,199
X696 VGND a_4839_12857# a_6129_12927# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5266,228
X697 a_2676_2157# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X698 a_11679_15219# a_8113_13753# a_11597_15219# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
X699 VGND VDPWR a_9685_10561# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X700 a_4213_5413# a_4159_5303# a_3820_5021# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X701 a_9699_4853# VDPWR a_10116_4597# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X702 a_15141_4951# VDPWR a_15045_4951# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X703 a_9587_15357# VGND VDPWR w_9490_15543# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X704 a_11019_12911# a_9811_11277# a_10937_12911# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X705 a_11243_11891# a_10965_11919# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X706 VGND VDPWR a_11916_2139# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X707 a_14136_4589# VDPWR a_13385_4845# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X708 a_4159_5303# a_3229_5051# a_4576_5047# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X709 VDPWR VDPWR a_15672_4585# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X710 VGND a_8785_5039# a_17346_5265# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=4514,209
X711 VGND VGND a_4183_2153# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X712 a_8596_5039# VDPWR a_7845_5295# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X713 VGND a_9290_1751# a_9238_1777# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X714 a_9875_13765# a_9597_13793# VDPWR w_9500_13979# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X715 a_18742_16187# a_18128_16189# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X716 a_7869_2145# a_6885_1783# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X717 a_8113_13753# a_7669_14003# VDPWR w_7604_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5930,268 d=10800,508
X718 a_6329_12927# a_5975_12927# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=5266,228 d=6760,364
X719 sky130_fd_sc_hd__mux4_1_0.A2 a_15185_2021# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X720 VDPWR VGND a_15936_1765# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X721 VGND VGND a_14066_2135# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X722 a_9725_5837# a_9671_5727# a_9332_5445# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X723 a_5945_2039# a_5069_1787# a_6362_1783# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X724 a_11455_4959# VDPWR a_11359_4959# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X725 sky130_fd_sc_hd__mux4_1_0.A0 a_22274_16171# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X726 a_10965_11919# a_9811_11277# VDPWR w_10868_12105# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X727 a_24318_14385# sky130_fd_sc_hd__mux4_1_0.A2 VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.10858 pd=1.36 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X728 a_11623_4593# a_11569_4849# a_11230_4567# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X729 a_9801_12841# VDPWR a_9717_12841# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X730 VDPWR VDPWR a_4627_12141# w_4530_12327# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X731 a_6281_11907# a_6003_11935# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X732 a_10380_1777# VDPWR a_9629_2033# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X733 VGND VDPWR a_10046_2143# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X734 a_4915_10549# a_4637_10577# VDPWR w_4540_10763# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X735 a_2343_5417# a_2217_5025# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X736 a_9290_1751# a_8755_1779# a_9515_1777# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X737 a_12976_1743# a_12439_1773# a_13201_2135# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X738 a_5831_1783# VDPWR a_5735_1783# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X739 a_24318_14385# a_23731_14309# a_24234_14385# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.10858 pd=1.36 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=4318,272
X740 a_9549_13091# VDPWR a_9467_13091# w_9394_13055# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X741 a_9477_11527# VDPWR VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X742 a_3229_5051# a_2289_5307# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X743 a_6087_14735# a_5809_14763# VDPWR w_5712_14949# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X744 VDPWR VDPWR a_4637_10577# w_4540_10763# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X745 VGND VDPWR a_6029_5409# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X746 a_12481_5467# a_11541_5723# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X747 a_11499_2029# a_10569_1777# a_11916_1773# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X748 a_13369_1769# a_13315_2025# a_12976_1743# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X749 a_11427_5467# VDPWR a_11331_5467# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X750 VGND VDPWR a_13369_2135# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X751 a_4753_16339# VGND VDPWR w_4430_16303# sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X752 a_2175_5051# VDPWR a_2079_5051# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X753 a_10450_4963# VDPWR a_9699_4853# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X754 VDPWR VDPWR a_9683_1777# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X755 a_4763_14775# VGND VDPWR w_4440_14739# sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X756 a_9360_4571# VDPWR a_9585_4963# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X757 a_18128_16189# a_17254_16187# VDPWR w_17940_16403# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X758 a_4910_5413# VDPWR a_4159_5303# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X759 a_13439_4955# a_13385_4845# a_13046_4563# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X760 VDPWR VGND a_8596_5039# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X761 a_10088_5837# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X762 a_15017_5825# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X763 a_7899_5405# a_7845_5295# a_7506_5013# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X764 a_10422_5471# VDPWR a_9671_5727# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X765 VGND VDPWR a_6362_2149# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X766 VDPWR VDPWR a_10116_4597# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X767 a_13046_4563# a_12509_4593# a_13271_4589# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X768 a_9332_5445# VGND a_9557_5471# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X769 a_9599_10561# VGND VDPWR w_9502_10747# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X770 a_11359_4593# VGND VDPWR w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X771 a_8785_5039# a_7845_5295# VDPWR w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X772 VGND a_3820_5021# a_3768_5047# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X773 a_11595_5833# a_10611_5471# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X774 VDPWR VDPWR a_7869_1779# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X775 VDPWR VDPWR a_13439_4589# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X776 a_7506_5013# a_6915_5043# a_7731_5039# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X777 VGND VDPWR a_15281_5825# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X778 VGND VGND a_7869_2145# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X779 a_9717_12841# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X780 a_8262_5039# VGND VDPWR w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X781 VDPWR VGND a_9557_14759# w_9402_14723# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X782 a_9867_12097# a_9589_12125# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X783 VDPWR VDPWR a_9725_5471# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X784 VDPWR VGND a_10380_1777# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X785 a_4839_12857# VDPWR a_4755_12857# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X786 a_3199_1791# a_2259_2047# VDPWR w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X787 a_12439_1773# a_11499_2029# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X788 a_9799_16073# a_9465_16323# a_9715_16323# w_9392_16287# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X789 a_12809_13987# a_11243_11891# a_12713_13987# w_12566_13951# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X790 a_2313_2157# a_2259_2047# a_1920_1765# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X791 VDPWR ui_in[1] a_23731_14309# sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.1083 ps=1.36 w=0.42 l=0.15
**devattr s=4332,272 d=4316,272
X792 a_1920_1765# a_2187_1765# a_2145_1791# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X793 VDPWR VGND a_4585_16339# w_4430_16303# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X794 a_17053_4938# a_16871_4938# VDPWR w_16764_4814# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X795 a_12075_13379# a_11824_13629# VDPWR w_11718_13593# sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5830,267 d=13600,536
X796 VDPWR VGND a_4595_14775# w_4440_14739# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X797 a_7701_2145# VDPWR a_7605_2145# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X798 VGND VGND a_10450_4963# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X799 a_15281_5825# a_15227_5715# a_14888_5433# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X800 a_10046_1777# VGND VDPWR w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X801 a_9419_1777# VGND VDPWR w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X802 VDPWR VDPWR a_2313_1791# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X803 a_13105_2135# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X804 VGND VGND a_4910_5413# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X805 a_2706_5051# VGND VDPWR w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X806 a_15227_5715# a_14297_5463# a_15644_5459# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X807 a_17254_16187# a_16486_16197# VDPWR w_17066_16401# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X808 VGND VGND a_6029_5409# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X809 a_14846_1739# a_14255_1769# a_15071_1765# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X810 a_6635_15235# a_6087_14735# VDPWR w_6570_15449# sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X811 a_5975_5299# a_5099_5047# a_6392_5043# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X812 a_11553_1773# a_10569_1777# VDPWR w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X813 ui_in[0] a_23731_14309# a_23511_14701# sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X814 VDPWR VGND a_10422_5471# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X815 VDPWR VGND a_9683_1777# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X816 VDPWR VDPWR a_15239_1765# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X817 a_10116_4963# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X818 a_9489_4963# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X819 a_13385_4845# a_12509_4593# a_13802_4955# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X820 a_24962_14701# ui_in[0] ui_in[0] sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09209 pd=0.99 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=3683,198
X821 a_3919_1787# VGND VDPWR w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X822 VDPWR a_13046_4563# a_12994_4589# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X823 VGND a_7113_13395# a_7669_14003# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2268,138 d=4075,198
X824 VGND a_9467_13091# a_9801_12841# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X825 a_10611_5471# a_9671_5727# VDPWR w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X826 a_2049_2157# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X827 a_9557_14759# VDPWR a_9475_14759# w_9402_14723# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X828 a_2343_5417# a_2289_5307# a_1950_5025# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X829 a_7845_5295# a_6915_5043# a_8262_5405# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X830 VDPWR a_9332_5445# a_9280_5471# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X831 VGND sky130_fd_sc_hd__mux4_1_0.A2 a_2187_1765# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X832 a_14946_4905# VDPWR a_15309_4951# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.07384 pd=0.80236 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X833 VGND VGND a_9753_4963# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X834 VDPWR VDPWR a_9725_14759# w_9402_14723# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X835 a_13175_4589# VGND VDPWR w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X836 a_4849_11293# VDPWR a_4765_11293# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X837 a_13411_5829# a_12481_5467# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X838 a_7731_5405# VDPWR a_7635_5405# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X839 a_14297_5463# a_13357_5719# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X840 VDPWR VGND a_13439_4589# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X841 a_9461_5471# VGND VDPWR w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X842 a_15239_2131# a_15185_2021# a_14846_1739# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X843 a_3010_2157# VDPWR a_2259_2047# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X844 a_7173_15235# a_6635_15235# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X845 a_13243_5463# VDPWR a_13147_5463# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X846 a_5851_13769# a_4837_16089# VDPWR w_5786_13983# sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X847 a_4849_11293# a_4515_11543# a_4765_11543# w_4442_11507# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X848 VDPWR VGND a_9725_5471# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X849 a_14255_1769# a_13315_2025# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X850 VGND a_4905_12113# a_6089_11935# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X851 a_4213_5047# a_3229_5051# VDPWR w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X852 a_5999_2149# a_5945_2039# a_5606_1757# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X853 a_4129_2043# a_3199_1791# a_4546_2153# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X854 a_9811_11277# a_9477_11527# a_9727_11527# w_9404_11491# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X855 a_20384_16179# a_19510_16177# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X856 a_6911_15235# a_6087_14735# a_6805_15235# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X857 VDPWR a_4839_12857# a_5851_13769# w_5786_13983# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X858 VDPWR a_1950_5025# a_1898_5051# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X859 a_8566_2145# VDPWR a_7815_2035# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X860 VDPWR VDPWR a_2676_1791# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X861 VDPWR VDPWR a_7899_5039# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
.ends

