magic
tech sky130A
magscale 1 2
timestamp 1754603109
<< nwell >>
rect 9392 16287 10112 16608
rect 9490 15543 10026 15864
rect 11532 15433 12252 15754
rect 9402 14723 10122 15044
rect 10674 14933 11210 15254
rect 9500 13979 10036 14300
rect 10748 13967 11468 14288
rect 12566 13951 13194 14272
rect 11718 13593 12254 13914
rect 9394 13055 10114 13376
rect 10872 13125 11408 13446
rect 9492 12311 10028 12632
rect 10868 12105 11404 12426
rect 9404 11491 10124 11812
rect 9502 10747 10038 11068
rect 6074 6018 6426 6339
rect 9180 5386 10728 5707
rect 11050 5382 12598 5703
rect 12866 5378 14414 5699
rect 14736 5374 16284 5695
rect 1798 4966 3346 5287
rect 3668 4962 5216 5283
rect 5484 4958 7032 5279
rect 7354 4954 8902 5275
rect 9208 4512 10756 4833
rect 11078 4508 12626 4829
rect 12894 4504 14442 4825
rect 14764 4500 16312 4821
rect 1768 1706 3316 2027
rect 3638 1702 5186 2023
rect 5454 1698 7002 2019
rect 7324 1694 8872 2015
rect 9138 1692 10686 2013
rect 11008 1688 12556 2009
rect 12824 1684 14372 2005
rect 14694 1680 16242 2001
<< pwell >>
rect 9439 16047 10073 16229
rect 9459 16009 9493 16047
rect 9757 15467 9947 15485
rect 9561 15303 9947 15467
rect 11986 15329 12213 15375
rect 9561 15299 9591 15303
rect 9557 15265 9591 15299
rect 11571 15193 12213 15329
rect 11599 15155 11633 15193
rect 10941 14857 11131 14875
rect 10745 14693 11131 14857
rect 10745 14689 10775 14693
rect 9449 14483 10083 14665
rect 10741 14655 10775 14689
rect 9469 14445 9503 14483
rect 9767 13903 9957 13921
rect 9571 13739 9957 13903
rect 11202 13863 11429 13909
rect 9571 13735 9601 13739
rect 9567 13701 9601 13735
rect 10787 13727 11429 13863
rect 10815 13689 10849 13727
rect 12966 13853 13155 13893
rect 12605 13717 13155 13853
rect 12634 13673 12668 13717
rect 12966 13711 13155 13717
rect 11967 13489 12153 13535
rect 11786 13353 12153 13489
rect 11786 13349 11819 13353
rect 11785 13315 11819 13349
rect 11185 13021 11369 13067
rect 9441 12815 10075 12997
rect 10911 12885 11369 13021
rect 10939 12847 10973 12885
rect 9461 12777 9495 12815
rect 9759 12235 9949 12253
rect 9563 12071 9949 12235
rect 9563 12067 9593 12071
rect 9559 12033 9593 12067
rect 11135 12029 11325 12047
rect 10939 11865 11325 12029
rect 10939 11861 10969 11865
rect 10935 11827 10969 11861
rect 9451 11251 10085 11433
rect 9471 11213 9505 11251
rect 9769 10671 9959 10689
rect 9573 10507 9959 10671
rect 9573 10503 9603 10507
rect 9569 10469 9603 10503
rect 6325 6583 6359 6617
rect 6325 6579 6346 6583
rect 6160 6397 6346 6579
rect 10626 5947 10660 5985
rect 9254 5811 10689 5947
rect 12496 5943 12530 5981
rect 9254 5765 9440 5811
rect 10503 5765 10689 5811
rect 11124 5807 12559 5943
rect 14312 5939 14346 5977
rect 11124 5761 11310 5807
rect 12373 5761 12559 5807
rect 12940 5803 14375 5939
rect 16182 5935 16216 5973
rect 12940 5757 13126 5803
rect 14189 5757 14375 5803
rect 14810 5799 16245 5935
rect 14810 5753 14996 5799
rect 16059 5753 16245 5799
rect 3244 5527 3278 5565
rect 1872 5391 3307 5527
rect 5114 5523 5148 5561
rect 1872 5345 2058 5391
rect 3121 5345 3307 5391
rect 3742 5387 5177 5523
rect 6930 5519 6964 5557
rect 3742 5341 3928 5387
rect 4991 5341 5177 5387
rect 5558 5383 6993 5519
rect 8800 5515 8834 5553
rect 5558 5337 5744 5383
rect 6807 5337 6993 5383
rect 7428 5379 8863 5515
rect 7428 5333 7614 5379
rect 8677 5333 8863 5379
rect 10654 5073 10688 5111
rect 9282 4937 10717 5073
rect 12524 5069 12558 5107
rect 9282 4891 9468 4937
rect 10531 4891 10717 4937
rect 11152 4933 12587 5069
rect 14340 5065 14374 5103
rect 11152 4887 11338 4933
rect 12401 4887 12587 4933
rect 12968 4929 14403 5065
rect 16210 5061 16244 5099
rect 12968 4883 13154 4929
rect 14217 4883 14403 4929
rect 14838 4925 16273 5061
rect 14838 4879 15024 4925
rect 16087 4879 16273 4925
rect 3214 2267 3248 2305
rect 1842 2131 3277 2267
rect 5084 2263 5118 2301
rect 1842 2085 2028 2131
rect 3091 2085 3277 2131
rect 3712 2127 5147 2263
rect 6900 2259 6934 2297
rect 3712 2081 3898 2127
rect 4961 2081 5147 2127
rect 5528 2123 6963 2259
rect 8770 2255 8804 2293
rect 5528 2077 5714 2123
rect 6777 2077 6963 2123
rect 7398 2119 8833 2255
rect 10584 2253 10618 2291
rect 7398 2073 7584 2119
rect 8647 2073 8833 2119
rect 9212 2117 10647 2253
rect 12454 2249 12488 2287
rect 9212 2071 9398 2117
rect 10461 2071 10647 2117
rect 11082 2113 12517 2249
rect 14270 2245 14304 2283
rect 11082 2067 11268 2113
rect 12331 2067 12517 2113
rect 12898 2109 14333 2245
rect 16140 2241 16174 2279
rect 12898 2063 13084 2109
rect 14147 2063 14333 2109
rect 14768 2105 16203 2241
rect 14768 2059 14954 2105
rect 16017 2059 16203 2105
<< ndiff >>
rect 9465 16121 9517 16203
rect 9465 16087 9473 16121
rect 9507 16087 9517 16121
rect 9465 16073 9517 16087
rect 9547 16143 9601 16203
rect 9547 16109 9557 16143
rect 9591 16109 9601 16143
rect 9547 16073 9601 16109
rect 9631 16121 9685 16203
rect 9631 16087 9641 16121
rect 9675 16087 9685 16121
rect 9631 16073 9685 16087
rect 9715 16073 9769 16203
rect 9799 16123 9953 16203
rect 9799 16089 9809 16123
rect 9843 16089 9909 16123
rect 9943 16089 9953 16123
rect 9799 16073 9953 16089
rect 9983 16194 10047 16203
rect 9983 16160 9999 16194
rect 10033 16160 10047 16194
rect 9983 16126 10047 16160
rect 9983 16092 9999 16126
rect 10033 16092 10047 16126
rect 9983 16073 10047 16092
rect 9783 15441 9835 15459
rect 9587 15403 9643 15441
rect 9587 15369 9599 15403
rect 9633 15369 9643 15403
rect 9587 15357 9643 15369
rect 9673 15357 9727 15441
rect 9757 15375 9835 15441
rect 9757 15357 9791 15375
rect 9783 15341 9791 15357
rect 9825 15341 9835 15375
rect 9783 15329 9835 15341
rect 9865 15375 9921 15459
rect 9865 15341 9875 15375
rect 9909 15341 9921 15375
rect 9865 15329 9921 15341
rect 12012 15333 12105 15349
rect 12012 15303 12046 15333
rect 11597 15273 11649 15303
rect 11597 15239 11605 15273
rect 11639 15239 11649 15273
rect 11597 15219 11649 15239
rect 11679 15219 11737 15303
rect 11767 15219 11843 15303
rect 11873 15219 11939 15303
rect 11969 15299 12046 15303
rect 12080 15299 12105 15333
rect 11969 15265 12105 15299
rect 11969 15231 12046 15265
rect 12080 15231 12105 15265
rect 11969 15219 12105 15231
rect 12135 15333 12187 15349
rect 12135 15299 12145 15333
rect 12179 15299 12187 15333
rect 12135 15265 12187 15299
rect 12135 15231 12145 15265
rect 12179 15231 12187 15265
rect 12135 15219 12187 15231
rect 10967 14831 11019 14849
rect 10771 14793 10827 14831
rect 10771 14759 10783 14793
rect 10817 14759 10827 14793
rect 10771 14747 10827 14759
rect 10857 14747 10911 14831
rect 10941 14765 11019 14831
rect 10941 14747 10975 14765
rect 10967 14731 10975 14747
rect 11009 14731 11019 14765
rect 10967 14719 11019 14731
rect 11049 14765 11105 14849
rect 11049 14731 11059 14765
rect 11093 14731 11105 14765
rect 11049 14719 11105 14731
rect 9475 14557 9527 14639
rect 9475 14523 9483 14557
rect 9517 14523 9527 14557
rect 9475 14509 9527 14523
rect 9557 14579 9611 14639
rect 9557 14545 9567 14579
rect 9601 14545 9611 14579
rect 9557 14509 9611 14545
rect 9641 14557 9695 14639
rect 9641 14523 9651 14557
rect 9685 14523 9695 14557
rect 9641 14509 9695 14523
rect 9725 14509 9779 14639
rect 9809 14559 9963 14639
rect 9809 14525 9819 14559
rect 9853 14525 9919 14559
rect 9953 14525 9963 14559
rect 9809 14509 9963 14525
rect 9993 14630 10057 14639
rect 9993 14596 10009 14630
rect 10043 14596 10057 14630
rect 9993 14562 10057 14596
rect 9993 14528 10009 14562
rect 10043 14528 10057 14562
rect 9993 14509 10057 14528
rect 9793 13877 9845 13895
rect 9597 13839 9653 13877
rect 9597 13805 9609 13839
rect 9643 13805 9653 13839
rect 9597 13793 9653 13805
rect 9683 13793 9737 13877
rect 9767 13811 9845 13877
rect 9767 13793 9801 13811
rect 9793 13777 9801 13793
rect 9835 13777 9845 13811
rect 9793 13765 9845 13777
rect 9875 13811 9931 13895
rect 11228 13867 11321 13883
rect 11228 13837 11262 13867
rect 9875 13777 9885 13811
rect 9919 13777 9931 13811
rect 9875 13765 9931 13777
rect 10813 13807 10865 13837
rect 10813 13773 10821 13807
rect 10855 13773 10865 13807
rect 10813 13753 10865 13773
rect 10895 13753 10953 13837
rect 10983 13753 11059 13837
rect 11089 13753 11155 13837
rect 11185 13833 11262 13837
rect 11296 13833 11321 13867
rect 11185 13799 11321 13833
rect 11185 13765 11262 13799
rect 11296 13765 11321 13799
rect 11185 13753 11321 13765
rect 11351 13867 11403 13883
rect 11351 13833 11361 13867
rect 11395 13833 11403 13867
rect 11351 13799 11403 13833
rect 11351 13765 11361 13799
rect 11395 13765 11403 13799
rect 11351 13753 11403 13765
rect 12992 13827 13045 13867
rect 12631 13807 12683 13827
rect 12631 13773 12639 13807
rect 12673 13773 12683 13807
rect 12631 13743 12683 13773
rect 12713 13801 12779 13827
rect 12713 13767 12729 13801
rect 12763 13767 12779 13801
rect 12713 13743 12779 13767
rect 12809 13787 12863 13827
rect 12809 13753 12819 13787
rect 12853 13753 12863 13787
rect 12809 13743 12863 13753
rect 12893 13801 12947 13827
rect 12893 13767 12903 13801
rect 12937 13767 12947 13801
rect 12893 13743 12947 13767
rect 12977 13787 13045 13827
rect 12977 13753 12997 13787
rect 13031 13753 13045 13787
rect 12977 13743 13045 13753
rect 12992 13737 13045 13743
rect 13075 13825 13129 13867
rect 13075 13791 13085 13825
rect 13119 13791 13129 13825
rect 13075 13737 13129 13791
rect 11993 13463 12045 13509
rect 11812 13435 11864 13463
rect 11812 13401 11820 13435
rect 11854 13401 11864 13435
rect 11812 13379 11864 13401
rect 11894 13435 11948 13463
rect 11894 13401 11904 13435
rect 11938 13401 11948 13435
rect 11894 13379 11948 13401
rect 11978 13435 12045 13463
rect 11978 13401 12000 13435
rect 12034 13401 12045 13435
rect 11978 13379 12045 13401
rect 12075 13495 12127 13509
rect 12075 13461 12085 13495
rect 12119 13461 12127 13495
rect 12075 13427 12127 13461
rect 12075 13393 12085 13427
rect 12119 13393 12127 13427
rect 12075 13379 12127 13393
rect 11211 12995 11261 13041
rect 9467 12889 9519 12971
rect 9467 12855 9475 12889
rect 9509 12855 9519 12889
rect 9467 12841 9519 12855
rect 9549 12911 9603 12971
rect 9549 12877 9559 12911
rect 9593 12877 9603 12911
rect 9549 12841 9603 12877
rect 9633 12889 9687 12971
rect 9633 12855 9643 12889
rect 9677 12855 9687 12889
rect 9633 12841 9687 12855
rect 9717 12841 9771 12971
rect 9801 12891 9955 12971
rect 9801 12857 9811 12891
rect 9845 12857 9911 12891
rect 9945 12857 9955 12891
rect 9801 12841 9955 12857
rect 9985 12962 10049 12971
rect 9985 12928 10001 12962
rect 10035 12928 10049 12962
rect 9985 12894 10049 12928
rect 10937 12957 10989 12995
rect 10937 12923 10945 12957
rect 10979 12923 10989 12957
rect 10937 12911 10989 12923
rect 11019 12911 11061 12995
rect 11091 12911 11133 12995
rect 11163 12973 11261 12995
rect 11163 12939 11217 12973
rect 11251 12939 11261 12973
rect 11163 12911 11261 12939
rect 11291 12983 11343 13041
rect 11291 12949 11301 12983
rect 11335 12949 11343 12983
rect 11291 12911 11343 12949
rect 9985 12860 10001 12894
rect 10035 12860 10049 12894
rect 9985 12841 10049 12860
rect 9785 12209 9837 12227
rect 9589 12171 9645 12209
rect 9589 12137 9601 12171
rect 9635 12137 9645 12171
rect 9589 12125 9645 12137
rect 9675 12125 9729 12209
rect 9759 12143 9837 12209
rect 9759 12125 9793 12143
rect 9785 12109 9793 12125
rect 9827 12109 9837 12143
rect 9785 12097 9837 12109
rect 9867 12143 9923 12227
rect 9867 12109 9877 12143
rect 9911 12109 9923 12143
rect 9867 12097 9923 12109
rect 11161 12003 11213 12021
rect 10965 11965 11021 12003
rect 10965 11931 10977 11965
rect 11011 11931 11021 11965
rect 10965 11919 11021 11931
rect 11051 11919 11105 12003
rect 11135 11937 11213 12003
rect 11135 11919 11169 11937
rect 11161 11903 11169 11919
rect 11203 11903 11213 11937
rect 11161 11891 11213 11903
rect 11243 11937 11299 12021
rect 11243 11903 11253 11937
rect 11287 11903 11299 11937
rect 11243 11891 11299 11903
rect 9477 11325 9529 11407
rect 9477 11291 9485 11325
rect 9519 11291 9529 11325
rect 9477 11277 9529 11291
rect 9559 11347 9613 11407
rect 9559 11313 9569 11347
rect 9603 11313 9613 11347
rect 9559 11277 9613 11313
rect 9643 11325 9697 11407
rect 9643 11291 9653 11325
rect 9687 11291 9697 11325
rect 9643 11277 9697 11291
rect 9727 11277 9781 11407
rect 9811 11327 9965 11407
rect 9811 11293 9821 11327
rect 9855 11293 9921 11327
rect 9955 11293 9965 11327
rect 9811 11277 9965 11293
rect 9995 11398 10059 11407
rect 9995 11364 10011 11398
rect 10045 11364 10059 11398
rect 9995 11330 10059 11364
rect 9995 11296 10011 11330
rect 10045 11296 10059 11330
rect 9995 11277 10059 11296
rect 9795 10645 9847 10663
rect 9599 10607 9655 10645
rect 9599 10573 9611 10607
rect 9645 10573 9655 10607
rect 9599 10561 9655 10573
rect 9685 10561 9739 10645
rect 9769 10579 9847 10645
rect 9769 10561 9803 10579
rect 9795 10545 9803 10561
rect 9837 10545 9847 10579
rect 9795 10533 9847 10545
rect 9877 10579 9933 10663
rect 9877 10545 9887 10579
rect 9921 10545 9933 10579
rect 9877 10533 9933 10545
rect 6186 6537 6238 6553
rect 6186 6503 6194 6537
rect 6228 6503 6238 6537
rect 6186 6469 6238 6503
rect 6186 6435 6194 6469
rect 6228 6435 6238 6469
rect 6186 6423 6238 6435
rect 6268 6537 6320 6553
rect 6268 6503 6278 6537
rect 6312 6503 6320 6537
rect 6268 6469 6320 6503
rect 6268 6435 6278 6469
rect 6312 6435 6320 6469
rect 6268 6423 6320 6435
rect 9280 5873 9332 5921
rect 9280 5839 9288 5873
rect 9322 5839 9332 5873
rect 9280 5791 9332 5839
rect 9362 5913 9431 5921
rect 9362 5879 9387 5913
rect 9421 5879 9431 5913
rect 9362 5837 9431 5879
rect 9461 5837 9527 5921
rect 9557 5837 9599 5921
rect 9629 5901 9695 5921
rect 9629 5867 9639 5901
rect 9673 5867 9695 5901
rect 9629 5837 9695 5867
rect 9725 5896 9784 5921
rect 9725 5862 9740 5896
rect 9774 5862 9784 5896
rect 9725 5837 9784 5862
rect 9814 5913 9868 5921
rect 9814 5879 9824 5913
rect 9858 5879 9868 5913
rect 9814 5837 9868 5879
rect 9898 5896 9952 5921
rect 9898 5862 9908 5896
rect 9942 5862 9952 5896
rect 9898 5837 9952 5862
rect 9982 5904 10034 5921
rect 9982 5870 9992 5904
rect 10026 5870 10034 5904
rect 9982 5837 10034 5870
rect 10088 5896 10140 5921
rect 10088 5862 10096 5896
rect 10130 5862 10140 5896
rect 10088 5837 10140 5862
rect 10170 5913 10224 5921
rect 10170 5879 10180 5913
rect 10214 5879 10224 5913
rect 10170 5837 10224 5879
rect 10254 5896 10308 5921
rect 10254 5862 10264 5896
rect 10298 5862 10308 5896
rect 10254 5837 10308 5862
rect 10338 5896 10392 5921
rect 10338 5862 10348 5896
rect 10382 5862 10392 5896
rect 10338 5837 10392 5862
rect 10422 5837 10482 5921
rect 10512 5909 10581 5921
rect 10512 5875 10537 5909
rect 10571 5875 10581 5909
rect 10512 5837 10581 5875
rect 9362 5791 9414 5837
rect 1898 5453 1950 5501
rect 1898 5419 1906 5453
rect 1940 5419 1950 5453
rect 1898 5371 1950 5419
rect 1980 5493 2049 5501
rect 1980 5459 2005 5493
rect 2039 5459 2049 5493
rect 1980 5417 2049 5459
rect 2079 5417 2145 5501
rect 2175 5417 2217 5501
rect 2247 5481 2313 5501
rect 2247 5447 2257 5481
rect 2291 5447 2313 5481
rect 2247 5417 2313 5447
rect 2343 5476 2402 5501
rect 2343 5442 2358 5476
rect 2392 5442 2402 5476
rect 2343 5417 2402 5442
rect 2432 5493 2486 5501
rect 2432 5459 2442 5493
rect 2476 5459 2486 5493
rect 2432 5417 2486 5459
rect 2516 5476 2570 5501
rect 2516 5442 2526 5476
rect 2560 5442 2570 5476
rect 2516 5417 2570 5442
rect 2600 5484 2652 5501
rect 2600 5450 2610 5484
rect 2644 5450 2652 5484
rect 2600 5417 2652 5450
rect 2706 5476 2758 5501
rect 2706 5442 2714 5476
rect 2748 5442 2758 5476
rect 2706 5417 2758 5442
rect 2788 5493 2842 5501
rect 2788 5459 2798 5493
rect 2832 5459 2842 5493
rect 2788 5417 2842 5459
rect 2872 5476 2926 5501
rect 2872 5442 2882 5476
rect 2916 5442 2926 5476
rect 2872 5417 2926 5442
rect 2956 5476 3010 5501
rect 2956 5442 2966 5476
rect 3000 5442 3010 5476
rect 2956 5417 3010 5442
rect 3040 5417 3100 5501
rect 3130 5489 3199 5501
rect 3130 5455 3155 5489
rect 3189 5455 3199 5489
rect 3130 5417 3199 5455
rect 1980 5371 2032 5417
rect 3147 5371 3199 5417
rect 3229 5453 3281 5501
rect 3229 5419 3239 5453
rect 3273 5419 3281 5453
rect 3229 5371 3281 5419
rect 3768 5449 3820 5497
rect 3768 5415 3776 5449
rect 3810 5415 3820 5449
rect 3768 5367 3820 5415
rect 3850 5489 3919 5497
rect 3850 5455 3875 5489
rect 3909 5455 3919 5489
rect 3850 5413 3919 5455
rect 3949 5413 4015 5497
rect 4045 5413 4087 5497
rect 4117 5477 4183 5497
rect 4117 5443 4127 5477
rect 4161 5443 4183 5477
rect 4117 5413 4183 5443
rect 4213 5472 4272 5497
rect 4213 5438 4228 5472
rect 4262 5438 4272 5472
rect 4213 5413 4272 5438
rect 4302 5489 4356 5497
rect 4302 5455 4312 5489
rect 4346 5455 4356 5489
rect 4302 5413 4356 5455
rect 4386 5472 4440 5497
rect 4386 5438 4396 5472
rect 4430 5438 4440 5472
rect 4386 5413 4440 5438
rect 4470 5480 4522 5497
rect 4470 5446 4480 5480
rect 4514 5446 4522 5480
rect 4470 5413 4522 5446
rect 4576 5472 4628 5497
rect 4576 5438 4584 5472
rect 4618 5438 4628 5472
rect 4576 5413 4628 5438
rect 4658 5489 4712 5497
rect 4658 5455 4668 5489
rect 4702 5455 4712 5489
rect 4658 5413 4712 5455
rect 4742 5472 4796 5497
rect 4742 5438 4752 5472
rect 4786 5438 4796 5472
rect 4742 5413 4796 5438
rect 4826 5472 4880 5497
rect 4826 5438 4836 5472
rect 4870 5438 4880 5472
rect 4826 5413 4880 5438
rect 4910 5413 4970 5497
rect 5000 5485 5069 5497
rect 5000 5451 5025 5485
rect 5059 5451 5069 5485
rect 5000 5413 5069 5451
rect 3850 5367 3902 5413
rect 5017 5367 5069 5413
rect 5099 5449 5151 5497
rect 5099 5415 5109 5449
rect 5143 5415 5151 5449
rect 5099 5367 5151 5415
rect 5584 5445 5636 5493
rect 5584 5411 5592 5445
rect 5626 5411 5636 5445
rect 5584 5363 5636 5411
rect 5666 5485 5735 5493
rect 5666 5451 5691 5485
rect 5725 5451 5735 5485
rect 5666 5409 5735 5451
rect 5765 5409 5831 5493
rect 5861 5409 5903 5493
rect 5933 5473 5999 5493
rect 5933 5439 5943 5473
rect 5977 5439 5999 5473
rect 5933 5409 5999 5439
rect 6029 5468 6088 5493
rect 6029 5434 6044 5468
rect 6078 5434 6088 5468
rect 6029 5409 6088 5434
rect 6118 5485 6172 5493
rect 6118 5451 6128 5485
rect 6162 5451 6172 5485
rect 6118 5409 6172 5451
rect 6202 5468 6256 5493
rect 6202 5434 6212 5468
rect 6246 5434 6256 5468
rect 6202 5409 6256 5434
rect 6286 5476 6338 5493
rect 6286 5442 6296 5476
rect 6330 5442 6338 5476
rect 6286 5409 6338 5442
rect 6392 5468 6444 5493
rect 6392 5434 6400 5468
rect 6434 5434 6444 5468
rect 6392 5409 6444 5434
rect 6474 5485 6528 5493
rect 6474 5451 6484 5485
rect 6518 5451 6528 5485
rect 6474 5409 6528 5451
rect 6558 5468 6612 5493
rect 6558 5434 6568 5468
rect 6602 5434 6612 5468
rect 6558 5409 6612 5434
rect 6642 5468 6696 5493
rect 6642 5434 6652 5468
rect 6686 5434 6696 5468
rect 6642 5409 6696 5434
rect 6726 5409 6786 5493
rect 6816 5481 6885 5493
rect 6816 5447 6841 5481
rect 6875 5447 6885 5481
rect 6816 5409 6885 5447
rect 5666 5363 5718 5409
rect 6833 5363 6885 5409
rect 6915 5445 6967 5493
rect 6915 5411 6925 5445
rect 6959 5411 6967 5445
rect 6915 5363 6967 5411
rect 7454 5441 7506 5489
rect 7454 5407 7462 5441
rect 7496 5407 7506 5441
rect 7454 5359 7506 5407
rect 7536 5481 7605 5489
rect 7536 5447 7561 5481
rect 7595 5447 7605 5481
rect 7536 5405 7605 5447
rect 7635 5405 7701 5489
rect 7731 5405 7773 5489
rect 7803 5469 7869 5489
rect 7803 5435 7813 5469
rect 7847 5435 7869 5469
rect 7803 5405 7869 5435
rect 7899 5464 7958 5489
rect 7899 5430 7914 5464
rect 7948 5430 7958 5464
rect 7899 5405 7958 5430
rect 7988 5481 8042 5489
rect 7988 5447 7998 5481
rect 8032 5447 8042 5481
rect 7988 5405 8042 5447
rect 8072 5464 8126 5489
rect 8072 5430 8082 5464
rect 8116 5430 8126 5464
rect 8072 5405 8126 5430
rect 8156 5472 8208 5489
rect 8156 5438 8166 5472
rect 8200 5438 8208 5472
rect 8156 5405 8208 5438
rect 8262 5464 8314 5489
rect 8262 5430 8270 5464
rect 8304 5430 8314 5464
rect 8262 5405 8314 5430
rect 8344 5481 8398 5489
rect 8344 5447 8354 5481
rect 8388 5447 8398 5481
rect 8344 5405 8398 5447
rect 8428 5464 8482 5489
rect 8428 5430 8438 5464
rect 8472 5430 8482 5464
rect 8428 5405 8482 5430
rect 8512 5464 8566 5489
rect 8512 5430 8522 5464
rect 8556 5430 8566 5464
rect 8512 5405 8566 5430
rect 8596 5405 8656 5489
rect 8686 5477 8755 5489
rect 8686 5443 8711 5477
rect 8745 5443 8755 5477
rect 8686 5405 8755 5443
rect 7536 5359 7588 5405
rect 8703 5359 8755 5405
rect 8785 5441 8837 5489
rect 10529 5791 10581 5837
rect 10611 5873 10663 5921
rect 10611 5839 10621 5873
rect 10655 5839 10663 5873
rect 10611 5791 10663 5839
rect 11150 5869 11202 5917
rect 11150 5835 11158 5869
rect 11192 5835 11202 5869
rect 11150 5787 11202 5835
rect 11232 5909 11301 5917
rect 11232 5875 11257 5909
rect 11291 5875 11301 5909
rect 11232 5833 11301 5875
rect 11331 5833 11397 5917
rect 11427 5833 11469 5917
rect 11499 5897 11565 5917
rect 11499 5863 11509 5897
rect 11543 5863 11565 5897
rect 11499 5833 11565 5863
rect 11595 5892 11654 5917
rect 11595 5858 11610 5892
rect 11644 5858 11654 5892
rect 11595 5833 11654 5858
rect 11684 5909 11738 5917
rect 11684 5875 11694 5909
rect 11728 5875 11738 5909
rect 11684 5833 11738 5875
rect 11768 5892 11822 5917
rect 11768 5858 11778 5892
rect 11812 5858 11822 5892
rect 11768 5833 11822 5858
rect 11852 5900 11904 5917
rect 11852 5866 11862 5900
rect 11896 5866 11904 5900
rect 11852 5833 11904 5866
rect 11958 5892 12010 5917
rect 11958 5858 11966 5892
rect 12000 5858 12010 5892
rect 11958 5833 12010 5858
rect 12040 5909 12094 5917
rect 12040 5875 12050 5909
rect 12084 5875 12094 5909
rect 12040 5833 12094 5875
rect 12124 5892 12178 5917
rect 12124 5858 12134 5892
rect 12168 5858 12178 5892
rect 12124 5833 12178 5858
rect 12208 5892 12262 5917
rect 12208 5858 12218 5892
rect 12252 5858 12262 5892
rect 12208 5833 12262 5858
rect 12292 5833 12352 5917
rect 12382 5905 12451 5917
rect 12382 5871 12407 5905
rect 12441 5871 12451 5905
rect 12382 5833 12451 5871
rect 11232 5787 11284 5833
rect 12399 5787 12451 5833
rect 12481 5869 12533 5917
rect 12481 5835 12491 5869
rect 12525 5835 12533 5869
rect 12481 5787 12533 5835
rect 12966 5865 13018 5913
rect 12966 5831 12974 5865
rect 13008 5831 13018 5865
rect 12966 5783 13018 5831
rect 13048 5905 13117 5913
rect 13048 5871 13073 5905
rect 13107 5871 13117 5905
rect 13048 5829 13117 5871
rect 13147 5829 13213 5913
rect 13243 5829 13285 5913
rect 13315 5893 13381 5913
rect 13315 5859 13325 5893
rect 13359 5859 13381 5893
rect 13315 5829 13381 5859
rect 13411 5888 13470 5913
rect 13411 5854 13426 5888
rect 13460 5854 13470 5888
rect 13411 5829 13470 5854
rect 13500 5905 13554 5913
rect 13500 5871 13510 5905
rect 13544 5871 13554 5905
rect 13500 5829 13554 5871
rect 13584 5888 13638 5913
rect 13584 5854 13594 5888
rect 13628 5854 13638 5888
rect 13584 5829 13638 5854
rect 13668 5896 13720 5913
rect 13668 5862 13678 5896
rect 13712 5862 13720 5896
rect 13668 5829 13720 5862
rect 13774 5888 13826 5913
rect 13774 5854 13782 5888
rect 13816 5854 13826 5888
rect 13774 5829 13826 5854
rect 13856 5905 13910 5913
rect 13856 5871 13866 5905
rect 13900 5871 13910 5905
rect 13856 5829 13910 5871
rect 13940 5888 13994 5913
rect 13940 5854 13950 5888
rect 13984 5854 13994 5888
rect 13940 5829 13994 5854
rect 14024 5888 14078 5913
rect 14024 5854 14034 5888
rect 14068 5854 14078 5888
rect 14024 5829 14078 5854
rect 14108 5829 14168 5913
rect 14198 5901 14267 5913
rect 14198 5867 14223 5901
rect 14257 5867 14267 5901
rect 14198 5829 14267 5867
rect 13048 5783 13100 5829
rect 14215 5783 14267 5829
rect 14297 5865 14349 5913
rect 14297 5831 14307 5865
rect 14341 5831 14349 5865
rect 14297 5783 14349 5831
rect 14836 5861 14888 5909
rect 14836 5827 14844 5861
rect 14878 5827 14888 5861
rect 14836 5779 14888 5827
rect 14918 5901 14987 5909
rect 14918 5867 14943 5901
rect 14977 5867 14987 5901
rect 14918 5825 14987 5867
rect 15017 5825 15083 5909
rect 15113 5825 15155 5909
rect 15185 5889 15251 5909
rect 15185 5855 15195 5889
rect 15229 5855 15251 5889
rect 15185 5825 15251 5855
rect 15281 5884 15340 5909
rect 15281 5850 15296 5884
rect 15330 5850 15340 5884
rect 15281 5825 15340 5850
rect 15370 5901 15424 5909
rect 15370 5867 15380 5901
rect 15414 5867 15424 5901
rect 15370 5825 15424 5867
rect 15454 5884 15508 5909
rect 15454 5850 15464 5884
rect 15498 5850 15508 5884
rect 15454 5825 15508 5850
rect 15538 5892 15590 5909
rect 15538 5858 15548 5892
rect 15582 5858 15590 5892
rect 15538 5825 15590 5858
rect 15644 5884 15696 5909
rect 15644 5850 15652 5884
rect 15686 5850 15696 5884
rect 15644 5825 15696 5850
rect 15726 5901 15780 5909
rect 15726 5867 15736 5901
rect 15770 5867 15780 5901
rect 15726 5825 15780 5867
rect 15810 5884 15864 5909
rect 15810 5850 15820 5884
rect 15854 5850 15864 5884
rect 15810 5825 15864 5850
rect 15894 5884 15948 5909
rect 15894 5850 15904 5884
rect 15938 5850 15948 5884
rect 15894 5825 15948 5850
rect 15978 5825 16038 5909
rect 16068 5897 16137 5909
rect 16068 5863 16093 5897
rect 16127 5863 16137 5897
rect 16068 5825 16137 5863
rect 14918 5779 14970 5825
rect 8785 5407 8795 5441
rect 8829 5407 8837 5441
rect 16085 5779 16137 5825
rect 16167 5861 16219 5909
rect 16167 5827 16177 5861
rect 16211 5827 16219 5861
rect 16167 5779 16219 5827
rect 8785 5359 8837 5407
rect 9308 4999 9360 5047
rect 9308 4965 9316 4999
rect 9350 4965 9360 4999
rect 9308 4917 9360 4965
rect 9390 5039 9459 5047
rect 9390 5005 9415 5039
rect 9449 5005 9459 5039
rect 9390 4963 9459 5005
rect 9489 4963 9555 5047
rect 9585 4963 9627 5047
rect 9657 5027 9723 5047
rect 9657 4993 9667 5027
rect 9701 4993 9723 5027
rect 9657 4963 9723 4993
rect 9753 5022 9812 5047
rect 9753 4988 9768 5022
rect 9802 4988 9812 5022
rect 9753 4963 9812 4988
rect 9842 5039 9896 5047
rect 9842 5005 9852 5039
rect 9886 5005 9896 5039
rect 9842 4963 9896 5005
rect 9926 5022 9980 5047
rect 9926 4988 9936 5022
rect 9970 4988 9980 5022
rect 9926 4963 9980 4988
rect 10010 5030 10062 5047
rect 10010 4996 10020 5030
rect 10054 4996 10062 5030
rect 10010 4963 10062 4996
rect 10116 5022 10168 5047
rect 10116 4988 10124 5022
rect 10158 4988 10168 5022
rect 10116 4963 10168 4988
rect 10198 5039 10252 5047
rect 10198 5005 10208 5039
rect 10242 5005 10252 5039
rect 10198 4963 10252 5005
rect 10282 5022 10336 5047
rect 10282 4988 10292 5022
rect 10326 4988 10336 5022
rect 10282 4963 10336 4988
rect 10366 5022 10420 5047
rect 10366 4988 10376 5022
rect 10410 4988 10420 5022
rect 10366 4963 10420 4988
rect 10450 4963 10510 5047
rect 10540 5035 10609 5047
rect 10540 5001 10565 5035
rect 10599 5001 10609 5035
rect 10540 4963 10609 5001
rect 9390 4917 9442 4963
rect 10557 4917 10609 4963
rect 10639 4999 10691 5047
rect 10639 4965 10649 4999
rect 10683 4965 10691 4999
rect 10639 4917 10691 4965
rect 11178 4995 11230 5043
rect 11178 4961 11186 4995
rect 11220 4961 11230 4995
rect 11178 4913 11230 4961
rect 11260 5035 11329 5043
rect 11260 5001 11285 5035
rect 11319 5001 11329 5035
rect 11260 4959 11329 5001
rect 11359 4959 11425 5043
rect 11455 4959 11497 5043
rect 11527 5023 11593 5043
rect 11527 4989 11537 5023
rect 11571 4989 11593 5023
rect 11527 4959 11593 4989
rect 11623 5018 11682 5043
rect 11623 4984 11638 5018
rect 11672 4984 11682 5018
rect 11623 4959 11682 4984
rect 11712 5035 11766 5043
rect 11712 5001 11722 5035
rect 11756 5001 11766 5035
rect 11712 4959 11766 5001
rect 11796 5018 11850 5043
rect 11796 4984 11806 5018
rect 11840 4984 11850 5018
rect 11796 4959 11850 4984
rect 11880 5026 11932 5043
rect 11880 4992 11890 5026
rect 11924 4992 11932 5026
rect 11880 4959 11932 4992
rect 11986 5018 12038 5043
rect 11986 4984 11994 5018
rect 12028 4984 12038 5018
rect 11986 4959 12038 4984
rect 12068 5035 12122 5043
rect 12068 5001 12078 5035
rect 12112 5001 12122 5035
rect 12068 4959 12122 5001
rect 12152 5018 12206 5043
rect 12152 4984 12162 5018
rect 12196 4984 12206 5018
rect 12152 4959 12206 4984
rect 12236 5018 12290 5043
rect 12236 4984 12246 5018
rect 12280 4984 12290 5018
rect 12236 4959 12290 4984
rect 12320 4959 12380 5043
rect 12410 5031 12479 5043
rect 12410 4997 12435 5031
rect 12469 4997 12479 5031
rect 12410 4959 12479 4997
rect 11260 4913 11312 4959
rect 12427 4913 12479 4959
rect 12509 4995 12561 5043
rect 12509 4961 12519 4995
rect 12553 4961 12561 4995
rect 12509 4913 12561 4961
rect 12994 4991 13046 5039
rect 12994 4957 13002 4991
rect 13036 4957 13046 4991
rect 12994 4909 13046 4957
rect 13076 5031 13145 5039
rect 13076 4997 13101 5031
rect 13135 4997 13145 5031
rect 13076 4955 13145 4997
rect 13175 4955 13241 5039
rect 13271 4955 13313 5039
rect 13343 5019 13409 5039
rect 13343 4985 13353 5019
rect 13387 4985 13409 5019
rect 13343 4955 13409 4985
rect 13439 5014 13498 5039
rect 13439 4980 13454 5014
rect 13488 4980 13498 5014
rect 13439 4955 13498 4980
rect 13528 5031 13582 5039
rect 13528 4997 13538 5031
rect 13572 4997 13582 5031
rect 13528 4955 13582 4997
rect 13612 5014 13666 5039
rect 13612 4980 13622 5014
rect 13656 4980 13666 5014
rect 13612 4955 13666 4980
rect 13696 5022 13748 5039
rect 13696 4988 13706 5022
rect 13740 4988 13748 5022
rect 13696 4955 13748 4988
rect 13802 5014 13854 5039
rect 13802 4980 13810 5014
rect 13844 4980 13854 5014
rect 13802 4955 13854 4980
rect 13884 5031 13938 5039
rect 13884 4997 13894 5031
rect 13928 4997 13938 5031
rect 13884 4955 13938 4997
rect 13968 5014 14022 5039
rect 13968 4980 13978 5014
rect 14012 4980 14022 5014
rect 13968 4955 14022 4980
rect 14052 5014 14106 5039
rect 14052 4980 14062 5014
rect 14096 4980 14106 5014
rect 14052 4955 14106 4980
rect 14136 4955 14196 5039
rect 14226 5027 14295 5039
rect 14226 4993 14251 5027
rect 14285 4993 14295 5027
rect 14226 4955 14295 4993
rect 13076 4909 13128 4955
rect 14243 4909 14295 4955
rect 14325 4991 14377 5039
rect 14325 4957 14335 4991
rect 14369 4957 14377 4991
rect 14325 4909 14377 4957
rect 14864 4987 14916 5035
rect 14864 4953 14872 4987
rect 14906 4953 14916 4987
rect 14864 4905 14916 4953
rect 14946 5027 15015 5035
rect 14946 4993 14971 5027
rect 15005 4993 15015 5027
rect 14946 4951 15015 4993
rect 15045 4951 15111 5035
rect 15141 4951 15183 5035
rect 15213 5015 15279 5035
rect 15213 4981 15223 5015
rect 15257 4981 15279 5015
rect 15213 4951 15279 4981
rect 15309 5010 15368 5035
rect 15309 4976 15324 5010
rect 15358 4976 15368 5010
rect 15309 4951 15368 4976
rect 15398 5027 15452 5035
rect 15398 4993 15408 5027
rect 15442 4993 15452 5027
rect 15398 4951 15452 4993
rect 15482 5010 15536 5035
rect 15482 4976 15492 5010
rect 15526 4976 15536 5010
rect 15482 4951 15536 4976
rect 15566 5018 15618 5035
rect 15566 4984 15576 5018
rect 15610 4984 15618 5018
rect 15566 4951 15618 4984
rect 15672 5010 15724 5035
rect 15672 4976 15680 5010
rect 15714 4976 15724 5010
rect 15672 4951 15724 4976
rect 15754 5027 15808 5035
rect 15754 4993 15764 5027
rect 15798 4993 15808 5027
rect 15754 4951 15808 4993
rect 15838 5010 15892 5035
rect 15838 4976 15848 5010
rect 15882 4976 15892 5010
rect 15838 4951 15892 4976
rect 15922 5010 15976 5035
rect 15922 4976 15932 5010
rect 15966 4976 15976 5010
rect 15922 4951 15976 4976
rect 16006 4951 16066 5035
rect 16096 5023 16165 5035
rect 16096 4989 16121 5023
rect 16155 4989 16165 5023
rect 16096 4951 16165 4989
rect 14946 4905 14998 4951
rect 16113 4905 16165 4951
rect 16195 4987 16247 5035
rect 16195 4953 16205 4987
rect 16239 4953 16247 4987
rect 16195 4905 16247 4953
rect 1868 2193 1920 2241
rect 1868 2159 1876 2193
rect 1910 2159 1920 2193
rect 1868 2111 1920 2159
rect 1950 2233 2019 2241
rect 1950 2199 1975 2233
rect 2009 2199 2019 2233
rect 1950 2157 2019 2199
rect 2049 2157 2115 2241
rect 2145 2157 2187 2241
rect 2217 2221 2283 2241
rect 2217 2187 2227 2221
rect 2261 2187 2283 2221
rect 2217 2157 2283 2187
rect 2313 2216 2372 2241
rect 2313 2182 2328 2216
rect 2362 2182 2372 2216
rect 2313 2157 2372 2182
rect 2402 2233 2456 2241
rect 2402 2199 2412 2233
rect 2446 2199 2456 2233
rect 2402 2157 2456 2199
rect 2486 2216 2540 2241
rect 2486 2182 2496 2216
rect 2530 2182 2540 2216
rect 2486 2157 2540 2182
rect 2570 2224 2622 2241
rect 2570 2190 2580 2224
rect 2614 2190 2622 2224
rect 2570 2157 2622 2190
rect 2676 2216 2728 2241
rect 2676 2182 2684 2216
rect 2718 2182 2728 2216
rect 2676 2157 2728 2182
rect 2758 2233 2812 2241
rect 2758 2199 2768 2233
rect 2802 2199 2812 2233
rect 2758 2157 2812 2199
rect 2842 2216 2896 2241
rect 2842 2182 2852 2216
rect 2886 2182 2896 2216
rect 2842 2157 2896 2182
rect 2926 2216 2980 2241
rect 2926 2182 2936 2216
rect 2970 2182 2980 2216
rect 2926 2157 2980 2182
rect 3010 2157 3070 2241
rect 3100 2229 3169 2241
rect 3100 2195 3125 2229
rect 3159 2195 3169 2229
rect 3100 2157 3169 2195
rect 1950 2111 2002 2157
rect 3117 2111 3169 2157
rect 3199 2193 3251 2241
rect 3199 2159 3209 2193
rect 3243 2159 3251 2193
rect 3199 2111 3251 2159
rect 3738 2189 3790 2237
rect 3738 2155 3746 2189
rect 3780 2155 3790 2189
rect 3738 2107 3790 2155
rect 3820 2229 3889 2237
rect 3820 2195 3845 2229
rect 3879 2195 3889 2229
rect 3820 2153 3889 2195
rect 3919 2153 3985 2237
rect 4015 2153 4057 2237
rect 4087 2217 4153 2237
rect 4087 2183 4097 2217
rect 4131 2183 4153 2217
rect 4087 2153 4153 2183
rect 4183 2212 4242 2237
rect 4183 2178 4198 2212
rect 4232 2178 4242 2212
rect 4183 2153 4242 2178
rect 4272 2229 4326 2237
rect 4272 2195 4282 2229
rect 4316 2195 4326 2229
rect 4272 2153 4326 2195
rect 4356 2212 4410 2237
rect 4356 2178 4366 2212
rect 4400 2178 4410 2212
rect 4356 2153 4410 2178
rect 4440 2220 4492 2237
rect 4440 2186 4450 2220
rect 4484 2186 4492 2220
rect 4440 2153 4492 2186
rect 4546 2212 4598 2237
rect 4546 2178 4554 2212
rect 4588 2178 4598 2212
rect 4546 2153 4598 2178
rect 4628 2229 4682 2237
rect 4628 2195 4638 2229
rect 4672 2195 4682 2229
rect 4628 2153 4682 2195
rect 4712 2212 4766 2237
rect 4712 2178 4722 2212
rect 4756 2178 4766 2212
rect 4712 2153 4766 2178
rect 4796 2212 4850 2237
rect 4796 2178 4806 2212
rect 4840 2178 4850 2212
rect 4796 2153 4850 2178
rect 4880 2153 4940 2237
rect 4970 2225 5039 2237
rect 4970 2191 4995 2225
rect 5029 2191 5039 2225
rect 4970 2153 5039 2191
rect 3820 2107 3872 2153
rect 4987 2107 5039 2153
rect 5069 2189 5121 2237
rect 5069 2155 5079 2189
rect 5113 2155 5121 2189
rect 5069 2107 5121 2155
rect 5554 2185 5606 2233
rect 5554 2151 5562 2185
rect 5596 2151 5606 2185
rect 5554 2103 5606 2151
rect 5636 2225 5705 2233
rect 5636 2191 5661 2225
rect 5695 2191 5705 2225
rect 5636 2149 5705 2191
rect 5735 2149 5801 2233
rect 5831 2149 5873 2233
rect 5903 2213 5969 2233
rect 5903 2179 5913 2213
rect 5947 2179 5969 2213
rect 5903 2149 5969 2179
rect 5999 2208 6058 2233
rect 5999 2174 6014 2208
rect 6048 2174 6058 2208
rect 5999 2149 6058 2174
rect 6088 2225 6142 2233
rect 6088 2191 6098 2225
rect 6132 2191 6142 2225
rect 6088 2149 6142 2191
rect 6172 2208 6226 2233
rect 6172 2174 6182 2208
rect 6216 2174 6226 2208
rect 6172 2149 6226 2174
rect 6256 2216 6308 2233
rect 6256 2182 6266 2216
rect 6300 2182 6308 2216
rect 6256 2149 6308 2182
rect 6362 2208 6414 2233
rect 6362 2174 6370 2208
rect 6404 2174 6414 2208
rect 6362 2149 6414 2174
rect 6444 2225 6498 2233
rect 6444 2191 6454 2225
rect 6488 2191 6498 2225
rect 6444 2149 6498 2191
rect 6528 2208 6582 2233
rect 6528 2174 6538 2208
rect 6572 2174 6582 2208
rect 6528 2149 6582 2174
rect 6612 2208 6666 2233
rect 6612 2174 6622 2208
rect 6656 2174 6666 2208
rect 6612 2149 6666 2174
rect 6696 2149 6756 2233
rect 6786 2221 6855 2233
rect 6786 2187 6811 2221
rect 6845 2187 6855 2221
rect 6786 2149 6855 2187
rect 5636 2103 5688 2149
rect 6803 2103 6855 2149
rect 6885 2185 6937 2233
rect 6885 2151 6895 2185
rect 6929 2151 6937 2185
rect 6885 2103 6937 2151
rect 7424 2181 7476 2229
rect 7424 2147 7432 2181
rect 7466 2147 7476 2181
rect 7424 2099 7476 2147
rect 7506 2221 7575 2229
rect 7506 2187 7531 2221
rect 7565 2187 7575 2221
rect 7506 2145 7575 2187
rect 7605 2145 7671 2229
rect 7701 2145 7743 2229
rect 7773 2209 7839 2229
rect 7773 2175 7783 2209
rect 7817 2175 7839 2209
rect 7773 2145 7839 2175
rect 7869 2204 7928 2229
rect 7869 2170 7884 2204
rect 7918 2170 7928 2204
rect 7869 2145 7928 2170
rect 7958 2221 8012 2229
rect 7958 2187 7968 2221
rect 8002 2187 8012 2221
rect 7958 2145 8012 2187
rect 8042 2204 8096 2229
rect 8042 2170 8052 2204
rect 8086 2170 8096 2204
rect 8042 2145 8096 2170
rect 8126 2212 8178 2229
rect 8126 2178 8136 2212
rect 8170 2178 8178 2212
rect 8126 2145 8178 2178
rect 8232 2204 8284 2229
rect 8232 2170 8240 2204
rect 8274 2170 8284 2204
rect 8232 2145 8284 2170
rect 8314 2221 8368 2229
rect 8314 2187 8324 2221
rect 8358 2187 8368 2221
rect 8314 2145 8368 2187
rect 8398 2204 8452 2229
rect 8398 2170 8408 2204
rect 8442 2170 8452 2204
rect 8398 2145 8452 2170
rect 8482 2204 8536 2229
rect 8482 2170 8492 2204
rect 8526 2170 8536 2204
rect 8482 2145 8536 2170
rect 8566 2145 8626 2229
rect 8656 2217 8725 2229
rect 8656 2183 8681 2217
rect 8715 2183 8725 2217
rect 8656 2145 8725 2183
rect 7506 2099 7558 2145
rect 8673 2099 8725 2145
rect 8755 2181 8807 2229
rect 8755 2147 8765 2181
rect 8799 2147 8807 2181
rect 8755 2099 8807 2147
rect 9238 2179 9290 2227
rect 9238 2145 9246 2179
rect 9280 2145 9290 2179
rect 9238 2097 9290 2145
rect 9320 2219 9389 2227
rect 9320 2185 9345 2219
rect 9379 2185 9389 2219
rect 9320 2143 9389 2185
rect 9419 2143 9485 2227
rect 9515 2143 9557 2227
rect 9587 2207 9653 2227
rect 9587 2173 9597 2207
rect 9631 2173 9653 2207
rect 9587 2143 9653 2173
rect 9683 2202 9742 2227
rect 9683 2168 9698 2202
rect 9732 2168 9742 2202
rect 9683 2143 9742 2168
rect 9772 2219 9826 2227
rect 9772 2185 9782 2219
rect 9816 2185 9826 2219
rect 9772 2143 9826 2185
rect 9856 2202 9910 2227
rect 9856 2168 9866 2202
rect 9900 2168 9910 2202
rect 9856 2143 9910 2168
rect 9940 2210 9992 2227
rect 9940 2176 9950 2210
rect 9984 2176 9992 2210
rect 9940 2143 9992 2176
rect 10046 2202 10098 2227
rect 10046 2168 10054 2202
rect 10088 2168 10098 2202
rect 10046 2143 10098 2168
rect 10128 2219 10182 2227
rect 10128 2185 10138 2219
rect 10172 2185 10182 2219
rect 10128 2143 10182 2185
rect 10212 2202 10266 2227
rect 10212 2168 10222 2202
rect 10256 2168 10266 2202
rect 10212 2143 10266 2168
rect 10296 2202 10350 2227
rect 10296 2168 10306 2202
rect 10340 2168 10350 2202
rect 10296 2143 10350 2168
rect 10380 2143 10440 2227
rect 10470 2215 10539 2227
rect 10470 2181 10495 2215
rect 10529 2181 10539 2215
rect 10470 2143 10539 2181
rect 9320 2097 9372 2143
rect 10487 2097 10539 2143
rect 10569 2179 10621 2227
rect 10569 2145 10579 2179
rect 10613 2145 10621 2179
rect 10569 2097 10621 2145
rect 11108 2175 11160 2223
rect 11108 2141 11116 2175
rect 11150 2141 11160 2175
rect 11108 2093 11160 2141
rect 11190 2215 11259 2223
rect 11190 2181 11215 2215
rect 11249 2181 11259 2215
rect 11190 2139 11259 2181
rect 11289 2139 11355 2223
rect 11385 2139 11427 2223
rect 11457 2203 11523 2223
rect 11457 2169 11467 2203
rect 11501 2169 11523 2203
rect 11457 2139 11523 2169
rect 11553 2198 11612 2223
rect 11553 2164 11568 2198
rect 11602 2164 11612 2198
rect 11553 2139 11612 2164
rect 11642 2215 11696 2223
rect 11642 2181 11652 2215
rect 11686 2181 11696 2215
rect 11642 2139 11696 2181
rect 11726 2198 11780 2223
rect 11726 2164 11736 2198
rect 11770 2164 11780 2198
rect 11726 2139 11780 2164
rect 11810 2206 11862 2223
rect 11810 2172 11820 2206
rect 11854 2172 11862 2206
rect 11810 2139 11862 2172
rect 11916 2198 11968 2223
rect 11916 2164 11924 2198
rect 11958 2164 11968 2198
rect 11916 2139 11968 2164
rect 11998 2215 12052 2223
rect 11998 2181 12008 2215
rect 12042 2181 12052 2215
rect 11998 2139 12052 2181
rect 12082 2198 12136 2223
rect 12082 2164 12092 2198
rect 12126 2164 12136 2198
rect 12082 2139 12136 2164
rect 12166 2198 12220 2223
rect 12166 2164 12176 2198
rect 12210 2164 12220 2198
rect 12166 2139 12220 2164
rect 12250 2139 12310 2223
rect 12340 2211 12409 2223
rect 12340 2177 12365 2211
rect 12399 2177 12409 2211
rect 12340 2139 12409 2177
rect 11190 2093 11242 2139
rect 12357 2093 12409 2139
rect 12439 2175 12491 2223
rect 12439 2141 12449 2175
rect 12483 2141 12491 2175
rect 12439 2093 12491 2141
rect 12924 2171 12976 2219
rect 12924 2137 12932 2171
rect 12966 2137 12976 2171
rect 12924 2089 12976 2137
rect 13006 2211 13075 2219
rect 13006 2177 13031 2211
rect 13065 2177 13075 2211
rect 13006 2135 13075 2177
rect 13105 2135 13171 2219
rect 13201 2135 13243 2219
rect 13273 2199 13339 2219
rect 13273 2165 13283 2199
rect 13317 2165 13339 2199
rect 13273 2135 13339 2165
rect 13369 2194 13428 2219
rect 13369 2160 13384 2194
rect 13418 2160 13428 2194
rect 13369 2135 13428 2160
rect 13458 2211 13512 2219
rect 13458 2177 13468 2211
rect 13502 2177 13512 2211
rect 13458 2135 13512 2177
rect 13542 2194 13596 2219
rect 13542 2160 13552 2194
rect 13586 2160 13596 2194
rect 13542 2135 13596 2160
rect 13626 2202 13678 2219
rect 13626 2168 13636 2202
rect 13670 2168 13678 2202
rect 13626 2135 13678 2168
rect 13732 2194 13784 2219
rect 13732 2160 13740 2194
rect 13774 2160 13784 2194
rect 13732 2135 13784 2160
rect 13814 2211 13868 2219
rect 13814 2177 13824 2211
rect 13858 2177 13868 2211
rect 13814 2135 13868 2177
rect 13898 2194 13952 2219
rect 13898 2160 13908 2194
rect 13942 2160 13952 2194
rect 13898 2135 13952 2160
rect 13982 2194 14036 2219
rect 13982 2160 13992 2194
rect 14026 2160 14036 2194
rect 13982 2135 14036 2160
rect 14066 2135 14126 2219
rect 14156 2207 14225 2219
rect 14156 2173 14181 2207
rect 14215 2173 14225 2207
rect 14156 2135 14225 2173
rect 13006 2089 13058 2135
rect 14173 2089 14225 2135
rect 14255 2171 14307 2219
rect 14255 2137 14265 2171
rect 14299 2137 14307 2171
rect 14255 2089 14307 2137
rect 14794 2167 14846 2215
rect 14794 2133 14802 2167
rect 14836 2133 14846 2167
rect 14794 2085 14846 2133
rect 14876 2207 14945 2215
rect 14876 2173 14901 2207
rect 14935 2173 14945 2207
rect 14876 2131 14945 2173
rect 14975 2131 15041 2215
rect 15071 2131 15113 2215
rect 15143 2195 15209 2215
rect 15143 2161 15153 2195
rect 15187 2161 15209 2195
rect 15143 2131 15209 2161
rect 15239 2190 15298 2215
rect 15239 2156 15254 2190
rect 15288 2156 15298 2190
rect 15239 2131 15298 2156
rect 15328 2207 15382 2215
rect 15328 2173 15338 2207
rect 15372 2173 15382 2207
rect 15328 2131 15382 2173
rect 15412 2190 15466 2215
rect 15412 2156 15422 2190
rect 15456 2156 15466 2190
rect 15412 2131 15466 2156
rect 15496 2198 15548 2215
rect 15496 2164 15506 2198
rect 15540 2164 15548 2198
rect 15496 2131 15548 2164
rect 15602 2190 15654 2215
rect 15602 2156 15610 2190
rect 15644 2156 15654 2190
rect 15602 2131 15654 2156
rect 15684 2207 15738 2215
rect 15684 2173 15694 2207
rect 15728 2173 15738 2207
rect 15684 2131 15738 2173
rect 15768 2190 15822 2215
rect 15768 2156 15778 2190
rect 15812 2156 15822 2190
rect 15768 2131 15822 2156
rect 15852 2190 15906 2215
rect 15852 2156 15862 2190
rect 15896 2156 15906 2190
rect 15852 2131 15906 2156
rect 15936 2131 15996 2215
rect 16026 2203 16095 2215
rect 16026 2169 16051 2203
rect 16085 2169 16095 2203
rect 16026 2131 16095 2169
rect 14876 2085 14928 2131
rect 16043 2085 16095 2131
rect 16125 2167 16177 2215
rect 16125 2133 16135 2167
rect 16169 2133 16177 2167
rect 16125 2085 16177 2133
<< pdiff >>
rect 9465 16511 9517 16523
rect 9465 16477 9473 16511
rect 9507 16477 9517 16511
rect 9465 16443 9517 16477
rect 9465 16409 9473 16443
rect 9507 16409 9517 16443
rect 9465 16323 9517 16409
rect 9547 16323 9601 16523
rect 9631 16501 9685 16523
rect 9631 16467 9641 16501
rect 9675 16467 9685 16501
rect 9631 16433 9685 16467
rect 9631 16399 9641 16433
rect 9675 16399 9685 16433
rect 9631 16323 9685 16399
rect 9715 16501 9769 16523
rect 9715 16467 9725 16501
rect 9759 16467 9769 16501
rect 9715 16433 9769 16467
rect 9715 16399 9725 16433
rect 9759 16399 9769 16433
rect 9715 16323 9769 16399
rect 9799 16501 9851 16523
rect 9799 16467 9809 16501
rect 9843 16467 9851 16501
rect 9799 16323 9851 16467
rect 9905 16501 9957 16523
rect 9905 16467 9913 16501
rect 9947 16467 9957 16501
rect 9905 16433 9957 16467
rect 9905 16399 9913 16433
rect 9947 16399 9957 16433
rect 9905 16323 9957 16399
rect 9987 16503 10047 16523
rect 9987 16469 9997 16503
rect 10031 16469 10047 16503
rect 9987 16435 10047 16469
rect 9987 16401 9997 16435
rect 10031 16401 10047 16435
rect 9987 16367 10047 16401
rect 9987 16333 9997 16367
rect 10031 16333 10047 16367
rect 9987 16323 10047 16333
rect 9783 15767 9835 15779
rect 9783 15737 9791 15767
rect 9587 15725 9643 15737
rect 9587 15691 9599 15725
rect 9633 15691 9643 15725
rect 9587 15653 9643 15691
rect 9673 15725 9727 15737
rect 9673 15691 9683 15725
rect 9717 15691 9727 15725
rect 9673 15653 9727 15691
rect 9757 15733 9791 15737
rect 9825 15733 9835 15767
rect 9757 15699 9835 15733
rect 9757 15665 9791 15699
rect 9825 15665 9835 15699
rect 9757 15653 9835 15665
rect 9773 15579 9835 15653
rect 9865 15767 9960 15779
rect 9865 15733 9895 15767
rect 9929 15733 9960 15767
rect 9865 15699 9960 15733
rect 9865 15665 9895 15699
rect 9929 15665 9960 15699
rect 9865 15579 9960 15665
rect 11597 15657 11649 15669
rect 11597 15623 11605 15657
rect 11639 15623 11649 15657
rect 11597 15585 11649 15623
rect 11679 15649 11749 15669
rect 11679 15615 11697 15649
rect 11731 15615 11749 15649
rect 11679 15585 11749 15615
rect 11779 15657 11853 15669
rect 11779 15623 11799 15657
rect 11833 15623 11853 15657
rect 11779 15585 11853 15623
rect 11883 15649 11939 15669
rect 11883 15615 11894 15649
rect 11928 15615 11939 15649
rect 11883 15585 11939 15615
rect 11969 15657 12105 15669
rect 11969 15623 12045 15657
rect 12079 15623 12105 15657
rect 11969 15589 12105 15623
rect 11969 15585 12045 15589
rect 11988 15555 12045 15585
rect 12079 15555 12105 15589
rect 11988 15469 12105 15555
rect 12135 15657 12187 15669
rect 12135 15623 12145 15657
rect 12179 15623 12187 15657
rect 12135 15589 12187 15623
rect 12135 15555 12145 15589
rect 12179 15555 12187 15589
rect 12135 15521 12187 15555
rect 12135 15487 12145 15521
rect 12179 15487 12187 15521
rect 12135 15469 12187 15487
rect 10967 15157 11019 15169
rect 10967 15127 10975 15157
rect 10771 15115 10827 15127
rect 10771 15081 10783 15115
rect 10817 15081 10827 15115
rect 10771 15043 10827 15081
rect 10857 15115 10911 15127
rect 10857 15081 10867 15115
rect 10901 15081 10911 15115
rect 10857 15043 10911 15081
rect 10941 15123 10975 15127
rect 11009 15123 11019 15157
rect 10941 15089 11019 15123
rect 10941 15055 10975 15089
rect 11009 15055 11019 15089
rect 10941 15043 11019 15055
rect 9475 14947 9527 14959
rect 9475 14913 9483 14947
rect 9517 14913 9527 14947
rect 9475 14879 9527 14913
rect 9475 14845 9483 14879
rect 9517 14845 9527 14879
rect 9475 14759 9527 14845
rect 9557 14759 9611 14959
rect 9641 14937 9695 14959
rect 9641 14903 9651 14937
rect 9685 14903 9695 14937
rect 9641 14869 9695 14903
rect 9641 14835 9651 14869
rect 9685 14835 9695 14869
rect 9641 14759 9695 14835
rect 9725 14937 9779 14959
rect 9725 14903 9735 14937
rect 9769 14903 9779 14937
rect 9725 14869 9779 14903
rect 9725 14835 9735 14869
rect 9769 14835 9779 14869
rect 9725 14759 9779 14835
rect 9809 14937 9861 14959
rect 9809 14903 9819 14937
rect 9853 14903 9861 14937
rect 9809 14759 9861 14903
rect 9915 14937 9967 14959
rect 9915 14903 9923 14937
rect 9957 14903 9967 14937
rect 9915 14869 9967 14903
rect 9915 14835 9923 14869
rect 9957 14835 9967 14869
rect 9915 14759 9967 14835
rect 9997 14939 10057 14959
rect 9997 14905 10007 14939
rect 10041 14905 10057 14939
rect 9997 14871 10057 14905
rect 9997 14837 10007 14871
rect 10041 14837 10057 14871
rect 9997 14803 10057 14837
rect 10957 14969 11019 15043
rect 11049 15157 11144 15169
rect 11049 15123 11079 15157
rect 11113 15123 11144 15157
rect 11049 15089 11144 15123
rect 11049 15055 11079 15089
rect 11113 15055 11144 15089
rect 11049 14969 11144 15055
rect 9997 14769 10007 14803
rect 10041 14769 10057 14803
rect 9997 14759 10057 14769
rect 9793 14203 9845 14215
rect 9793 14173 9801 14203
rect 9597 14161 9653 14173
rect 9597 14127 9609 14161
rect 9643 14127 9653 14161
rect 9597 14089 9653 14127
rect 9683 14161 9737 14173
rect 9683 14127 9693 14161
rect 9727 14127 9737 14161
rect 9683 14089 9737 14127
rect 9767 14169 9801 14173
rect 9835 14169 9845 14203
rect 9767 14135 9845 14169
rect 9767 14101 9801 14135
rect 9835 14101 9845 14135
rect 9767 14089 9845 14101
rect 9783 14015 9845 14089
rect 9875 14203 9970 14215
rect 9875 14169 9905 14203
rect 9939 14169 9970 14203
rect 9875 14135 9970 14169
rect 9875 14101 9905 14135
rect 9939 14101 9970 14135
rect 10813 14191 10865 14203
rect 10813 14157 10821 14191
rect 10855 14157 10865 14191
rect 10813 14119 10865 14157
rect 10895 14183 10965 14203
rect 10895 14149 10913 14183
rect 10947 14149 10965 14183
rect 10895 14119 10965 14149
rect 10995 14191 11069 14203
rect 10995 14157 11015 14191
rect 11049 14157 11069 14191
rect 10995 14119 11069 14157
rect 11099 14183 11155 14203
rect 11099 14149 11110 14183
rect 11144 14149 11155 14183
rect 11099 14119 11155 14149
rect 11185 14191 11321 14203
rect 11185 14157 11261 14191
rect 11295 14157 11321 14191
rect 11185 14123 11321 14157
rect 11185 14119 11261 14123
rect 9875 14015 9970 14101
rect 11204 14089 11261 14119
rect 11295 14089 11321 14123
rect 11204 14003 11321 14089
rect 11351 14191 11403 14203
rect 11351 14157 11361 14191
rect 11395 14157 11403 14191
rect 12992 14175 13045 14187
rect 11351 14123 11403 14157
rect 11351 14089 11361 14123
rect 11395 14089 11403 14123
rect 12992 14141 13000 14175
rect 13034 14141 13045 14175
rect 11351 14055 11403 14089
rect 12992 14107 13045 14141
rect 12992 14073 13000 14107
rect 13034 14073 13045 14107
rect 12992 14071 13045 14073
rect 11351 14021 11361 14055
rect 11395 14021 11403 14055
rect 11351 14003 11403 14021
rect 12631 14044 12683 14071
rect 12631 14010 12639 14044
rect 12673 14010 12683 14044
rect 12631 13987 12683 14010
rect 12713 13987 12779 14071
rect 12809 13987 12851 14071
rect 12881 13987 12947 14071
rect 12977 13987 13045 14071
rect 13075 14144 13129 14187
rect 13075 14110 13085 14144
rect 13119 14110 13129 14144
rect 13075 14076 13129 14110
rect 13075 14042 13085 14076
rect 13119 14042 13129 14076
rect 13075 13987 13129 14042
rect 11993 13801 12045 13829
rect 11993 13767 12001 13801
rect 12035 13767 12045 13801
rect 11993 13733 12045 13767
rect 11993 13713 12001 13733
rect 11824 13681 11876 13713
rect 11824 13647 11832 13681
rect 11866 13647 11876 13681
rect 11824 13629 11876 13647
rect 11906 13629 11948 13713
rect 11978 13699 12001 13713
rect 12035 13699 12045 13733
rect 11978 13629 12045 13699
rect 12075 13817 12143 13829
rect 12075 13783 12101 13817
rect 12135 13783 12143 13817
rect 12075 13749 12143 13783
rect 12075 13715 12101 13749
rect 12135 13715 12143 13749
rect 12075 13629 12143 13715
rect 9467 13279 9519 13291
rect 9467 13245 9475 13279
rect 9509 13245 9519 13279
rect 9467 13211 9519 13245
rect 9467 13177 9475 13211
rect 9509 13177 9519 13211
rect 9467 13091 9519 13177
rect 9549 13091 9603 13291
rect 9633 13269 9687 13291
rect 9633 13235 9643 13269
rect 9677 13235 9687 13269
rect 9633 13201 9687 13235
rect 9633 13167 9643 13201
rect 9677 13167 9687 13201
rect 9633 13091 9687 13167
rect 9717 13269 9771 13291
rect 9717 13235 9727 13269
rect 9761 13235 9771 13269
rect 9717 13201 9771 13235
rect 9717 13167 9727 13201
rect 9761 13167 9771 13201
rect 9717 13091 9771 13167
rect 9801 13269 9853 13291
rect 9801 13235 9811 13269
rect 9845 13235 9853 13269
rect 9801 13091 9853 13235
rect 9907 13269 9959 13291
rect 9907 13235 9915 13269
rect 9949 13235 9959 13269
rect 9907 13201 9959 13235
rect 9907 13167 9915 13201
rect 9949 13167 9959 13201
rect 9907 13091 9959 13167
rect 9989 13271 10049 13291
rect 11209 13349 11261 13361
rect 11209 13315 11217 13349
rect 11251 13315 11261 13349
rect 11209 13302 11261 13315
rect 9989 13237 9999 13271
rect 10033 13237 10049 13271
rect 11211 13248 11261 13302
rect 9989 13203 10049 13237
rect 9989 13169 9999 13203
rect 10033 13169 10049 13203
rect 9989 13135 10049 13169
rect 10937 13210 10989 13248
rect 10937 13176 10945 13210
rect 10979 13176 10989 13210
rect 10937 13164 10989 13176
rect 11019 13240 11073 13248
rect 11019 13206 11029 13240
rect 11063 13206 11073 13240
rect 11019 13164 11073 13206
rect 11103 13221 11166 13248
rect 11103 13187 11122 13221
rect 11156 13187 11166 13221
rect 11103 13164 11166 13187
rect 11196 13164 11261 13248
rect 9989 13101 9999 13135
rect 10033 13101 10049 13135
rect 9989 13091 10049 13101
rect 11211 13161 11261 13164
rect 11291 13335 11343 13361
rect 11291 13301 11301 13335
rect 11335 13301 11343 13335
rect 11291 13267 11343 13301
rect 11291 13233 11301 13267
rect 11335 13233 11343 13267
rect 11291 13161 11343 13233
rect 9785 12535 9837 12547
rect 9785 12505 9793 12535
rect 9589 12493 9645 12505
rect 9589 12459 9601 12493
rect 9635 12459 9645 12493
rect 9589 12421 9645 12459
rect 9675 12493 9729 12505
rect 9675 12459 9685 12493
rect 9719 12459 9729 12493
rect 9675 12421 9729 12459
rect 9759 12501 9793 12505
rect 9827 12501 9837 12535
rect 9759 12467 9837 12501
rect 9759 12433 9793 12467
rect 9827 12433 9837 12467
rect 9759 12421 9837 12433
rect 9775 12347 9837 12421
rect 9867 12535 9962 12547
rect 9867 12501 9897 12535
rect 9931 12501 9962 12535
rect 9867 12467 9962 12501
rect 9867 12433 9897 12467
rect 9931 12433 9962 12467
rect 9867 12347 9962 12433
rect 11161 12329 11213 12341
rect 11161 12299 11169 12329
rect 10965 12287 11021 12299
rect 10965 12253 10977 12287
rect 11011 12253 11021 12287
rect 10965 12215 11021 12253
rect 11051 12287 11105 12299
rect 11051 12253 11061 12287
rect 11095 12253 11105 12287
rect 11051 12215 11105 12253
rect 11135 12295 11169 12299
rect 11203 12295 11213 12329
rect 11135 12261 11213 12295
rect 11135 12227 11169 12261
rect 11203 12227 11213 12261
rect 11135 12215 11213 12227
rect 11151 12141 11213 12215
rect 11243 12329 11338 12341
rect 11243 12295 11273 12329
rect 11307 12295 11338 12329
rect 11243 12261 11338 12295
rect 11243 12227 11273 12261
rect 11307 12227 11338 12261
rect 11243 12141 11338 12227
rect 9477 11715 9529 11727
rect 9477 11681 9485 11715
rect 9519 11681 9529 11715
rect 9477 11647 9529 11681
rect 9477 11613 9485 11647
rect 9519 11613 9529 11647
rect 9477 11527 9529 11613
rect 9559 11527 9613 11727
rect 9643 11705 9697 11727
rect 9643 11671 9653 11705
rect 9687 11671 9697 11705
rect 9643 11637 9697 11671
rect 9643 11603 9653 11637
rect 9687 11603 9697 11637
rect 9643 11527 9697 11603
rect 9727 11705 9781 11727
rect 9727 11671 9737 11705
rect 9771 11671 9781 11705
rect 9727 11637 9781 11671
rect 9727 11603 9737 11637
rect 9771 11603 9781 11637
rect 9727 11527 9781 11603
rect 9811 11705 9863 11727
rect 9811 11671 9821 11705
rect 9855 11671 9863 11705
rect 9811 11527 9863 11671
rect 9917 11705 9969 11727
rect 9917 11671 9925 11705
rect 9959 11671 9969 11705
rect 9917 11637 9969 11671
rect 9917 11603 9925 11637
rect 9959 11603 9969 11637
rect 9917 11527 9969 11603
rect 9999 11707 10059 11727
rect 9999 11673 10009 11707
rect 10043 11673 10059 11707
rect 9999 11639 10059 11673
rect 9999 11605 10009 11639
rect 10043 11605 10059 11639
rect 9999 11571 10059 11605
rect 9999 11537 10009 11571
rect 10043 11537 10059 11571
rect 9999 11527 10059 11537
rect 9795 10971 9847 10983
rect 9795 10941 9803 10971
rect 9599 10929 9655 10941
rect 9599 10895 9611 10929
rect 9645 10895 9655 10929
rect 9599 10857 9655 10895
rect 9685 10929 9739 10941
rect 9685 10895 9695 10929
rect 9729 10895 9739 10929
rect 9685 10857 9739 10895
rect 9769 10937 9803 10941
rect 9837 10937 9847 10971
rect 9769 10903 9847 10937
rect 9769 10869 9803 10903
rect 9837 10869 9847 10903
rect 9769 10857 9847 10869
rect 9785 10783 9847 10857
rect 9877 10971 9972 10983
rect 9877 10937 9907 10971
rect 9941 10937 9972 10971
rect 9877 10903 9972 10937
rect 9877 10869 9907 10903
rect 9941 10869 9972 10903
rect 9877 10783 9972 10869
rect 6186 6285 6238 6303
rect 6186 6251 6194 6285
rect 6228 6251 6238 6285
rect 6186 6217 6238 6251
rect 6186 6183 6194 6217
rect 6228 6183 6238 6217
rect 6186 6149 6238 6183
rect 6186 6115 6194 6149
rect 6228 6115 6238 6149
rect 6186 6103 6238 6115
rect 6268 6285 6320 6303
rect 6268 6251 6278 6285
rect 6312 6251 6320 6285
rect 6268 6217 6320 6251
rect 6268 6183 6278 6217
rect 6312 6183 6320 6217
rect 6268 6149 6320 6183
rect 6268 6115 6278 6149
rect 6312 6115 6320 6149
rect 6268 6103 6320 6115
rect 9280 5633 9332 5671
rect 9280 5599 9288 5633
rect 9322 5599 9332 5633
rect 9280 5543 9332 5599
rect 1898 5213 1950 5251
rect 1898 5179 1906 5213
rect 1940 5179 1950 5213
rect 1898 5123 1950 5179
rect 1898 5089 1906 5123
rect 1940 5089 1950 5123
rect 1898 5051 1950 5089
rect 1980 5135 2032 5251
rect 3147 5135 3199 5251
rect 1980 5093 2049 5135
rect 1980 5059 1990 5093
rect 2024 5059 2049 5093
rect 1980 5051 2049 5059
rect 2079 5051 2145 5135
rect 2175 5051 2217 5135
rect 2247 5105 2313 5135
rect 2247 5071 2257 5105
rect 2291 5071 2313 5105
rect 2247 5051 2313 5071
rect 2343 5110 2402 5135
rect 2343 5076 2358 5110
rect 2392 5076 2402 5110
rect 2343 5051 2402 5076
rect 2432 5093 2486 5135
rect 2432 5059 2442 5093
rect 2476 5059 2486 5093
rect 2432 5051 2486 5059
rect 2516 5110 2570 5135
rect 2516 5076 2526 5110
rect 2560 5076 2570 5110
rect 2516 5051 2570 5076
rect 2600 5097 2652 5135
rect 2600 5063 2610 5097
rect 2644 5063 2652 5097
rect 2600 5051 2652 5063
rect 2706 5110 2758 5135
rect 2706 5076 2714 5110
rect 2748 5076 2758 5110
rect 2706 5051 2758 5076
rect 2788 5093 2842 5135
rect 2788 5059 2798 5093
rect 2832 5059 2842 5093
rect 2788 5051 2842 5059
rect 2872 5110 2926 5135
rect 2872 5076 2882 5110
rect 2916 5076 2926 5110
rect 2872 5051 2926 5076
rect 2956 5110 3010 5135
rect 2956 5076 2966 5110
rect 3000 5076 3010 5110
rect 2956 5051 3010 5076
rect 3040 5051 3100 5135
rect 3130 5101 3199 5135
rect 3130 5067 3155 5101
rect 3189 5067 3199 5101
rect 3130 5051 3199 5067
rect 3229 5210 3281 5251
rect 3229 5176 3239 5210
rect 3273 5176 3281 5210
rect 3229 5116 3281 5176
rect 3229 5082 3239 5116
rect 3273 5082 3281 5116
rect 3229 5051 3281 5082
rect 3768 5209 3820 5247
rect 3768 5175 3776 5209
rect 3810 5175 3820 5209
rect 3768 5119 3820 5175
rect 3768 5085 3776 5119
rect 3810 5085 3820 5119
rect 3768 5047 3820 5085
rect 3850 5131 3902 5247
rect 5017 5131 5069 5247
rect 3850 5089 3919 5131
rect 3850 5055 3860 5089
rect 3894 5055 3919 5089
rect 3850 5047 3919 5055
rect 3949 5047 4015 5131
rect 4045 5047 4087 5131
rect 4117 5101 4183 5131
rect 4117 5067 4127 5101
rect 4161 5067 4183 5101
rect 4117 5047 4183 5067
rect 4213 5106 4272 5131
rect 4213 5072 4228 5106
rect 4262 5072 4272 5106
rect 4213 5047 4272 5072
rect 4302 5089 4356 5131
rect 4302 5055 4312 5089
rect 4346 5055 4356 5089
rect 4302 5047 4356 5055
rect 4386 5106 4440 5131
rect 4386 5072 4396 5106
rect 4430 5072 4440 5106
rect 4386 5047 4440 5072
rect 4470 5093 4522 5131
rect 4470 5059 4480 5093
rect 4514 5059 4522 5093
rect 4470 5047 4522 5059
rect 4576 5106 4628 5131
rect 4576 5072 4584 5106
rect 4618 5072 4628 5106
rect 4576 5047 4628 5072
rect 4658 5089 4712 5131
rect 4658 5055 4668 5089
rect 4702 5055 4712 5089
rect 4658 5047 4712 5055
rect 4742 5106 4796 5131
rect 4742 5072 4752 5106
rect 4786 5072 4796 5106
rect 4742 5047 4796 5072
rect 4826 5106 4880 5131
rect 4826 5072 4836 5106
rect 4870 5072 4880 5106
rect 4826 5047 4880 5072
rect 4910 5047 4970 5131
rect 5000 5097 5069 5131
rect 5000 5063 5025 5097
rect 5059 5063 5069 5097
rect 5000 5047 5069 5063
rect 5099 5206 5151 5247
rect 5099 5172 5109 5206
rect 5143 5172 5151 5206
rect 5099 5112 5151 5172
rect 5099 5078 5109 5112
rect 5143 5078 5151 5112
rect 5099 5047 5151 5078
rect 5584 5205 5636 5243
rect 5584 5171 5592 5205
rect 5626 5171 5636 5205
rect 5584 5115 5636 5171
rect 5584 5081 5592 5115
rect 5626 5081 5636 5115
rect 5584 5043 5636 5081
rect 5666 5127 5718 5243
rect 9280 5509 9288 5543
rect 9322 5509 9332 5543
rect 6833 5127 6885 5243
rect 5666 5085 5735 5127
rect 5666 5051 5676 5085
rect 5710 5051 5735 5085
rect 5666 5043 5735 5051
rect 5765 5043 5831 5127
rect 5861 5043 5903 5127
rect 5933 5097 5999 5127
rect 5933 5063 5943 5097
rect 5977 5063 5999 5097
rect 5933 5043 5999 5063
rect 6029 5102 6088 5127
rect 6029 5068 6044 5102
rect 6078 5068 6088 5102
rect 6029 5043 6088 5068
rect 6118 5085 6172 5127
rect 6118 5051 6128 5085
rect 6162 5051 6172 5085
rect 6118 5043 6172 5051
rect 6202 5102 6256 5127
rect 6202 5068 6212 5102
rect 6246 5068 6256 5102
rect 6202 5043 6256 5068
rect 6286 5089 6338 5127
rect 6286 5055 6296 5089
rect 6330 5055 6338 5089
rect 6286 5043 6338 5055
rect 6392 5102 6444 5127
rect 6392 5068 6400 5102
rect 6434 5068 6444 5102
rect 6392 5043 6444 5068
rect 6474 5085 6528 5127
rect 6474 5051 6484 5085
rect 6518 5051 6528 5085
rect 6474 5043 6528 5051
rect 6558 5102 6612 5127
rect 6558 5068 6568 5102
rect 6602 5068 6612 5102
rect 6558 5043 6612 5068
rect 6642 5102 6696 5127
rect 6642 5068 6652 5102
rect 6686 5068 6696 5102
rect 6642 5043 6696 5068
rect 6726 5043 6786 5127
rect 6816 5093 6885 5127
rect 6816 5059 6841 5093
rect 6875 5059 6885 5093
rect 6816 5043 6885 5059
rect 6915 5202 6967 5243
rect 6915 5168 6925 5202
rect 6959 5168 6967 5202
rect 6915 5108 6967 5168
rect 6915 5074 6925 5108
rect 6959 5074 6967 5108
rect 6915 5043 6967 5074
rect 7454 5201 7506 5239
rect 7454 5167 7462 5201
rect 7496 5167 7506 5201
rect 7454 5111 7506 5167
rect 7454 5077 7462 5111
rect 7496 5077 7506 5111
rect 7454 5039 7506 5077
rect 7536 5123 7588 5239
rect 9280 5471 9332 5509
rect 9362 5555 9414 5671
rect 10529 5555 10581 5671
rect 9362 5513 9431 5555
rect 9362 5479 9372 5513
rect 9406 5479 9431 5513
rect 9362 5471 9431 5479
rect 9461 5471 9527 5555
rect 9557 5471 9599 5555
rect 9629 5525 9695 5555
rect 9629 5491 9639 5525
rect 9673 5491 9695 5525
rect 9629 5471 9695 5491
rect 9725 5530 9784 5555
rect 9725 5496 9740 5530
rect 9774 5496 9784 5530
rect 9725 5471 9784 5496
rect 9814 5513 9868 5555
rect 9814 5479 9824 5513
rect 9858 5479 9868 5513
rect 9814 5471 9868 5479
rect 9898 5530 9952 5555
rect 9898 5496 9908 5530
rect 9942 5496 9952 5530
rect 9898 5471 9952 5496
rect 9982 5517 10034 5555
rect 9982 5483 9992 5517
rect 10026 5483 10034 5517
rect 9982 5471 10034 5483
rect 10088 5530 10140 5555
rect 10088 5496 10096 5530
rect 10130 5496 10140 5530
rect 10088 5471 10140 5496
rect 10170 5513 10224 5555
rect 10170 5479 10180 5513
rect 10214 5479 10224 5513
rect 10170 5471 10224 5479
rect 10254 5530 10308 5555
rect 10254 5496 10264 5530
rect 10298 5496 10308 5530
rect 10254 5471 10308 5496
rect 10338 5530 10392 5555
rect 10338 5496 10348 5530
rect 10382 5496 10392 5530
rect 10338 5471 10392 5496
rect 10422 5471 10482 5555
rect 10512 5521 10581 5555
rect 10512 5487 10537 5521
rect 10571 5487 10581 5521
rect 10512 5471 10581 5487
rect 10611 5630 10663 5671
rect 10611 5596 10621 5630
rect 10655 5596 10663 5630
rect 10611 5536 10663 5596
rect 10611 5502 10621 5536
rect 10655 5502 10663 5536
rect 10611 5471 10663 5502
rect 11150 5629 11202 5667
rect 11150 5595 11158 5629
rect 11192 5595 11202 5629
rect 11150 5539 11202 5595
rect 11150 5505 11158 5539
rect 11192 5505 11202 5539
rect 11150 5467 11202 5505
rect 11232 5551 11284 5667
rect 12399 5551 12451 5667
rect 11232 5509 11301 5551
rect 11232 5475 11242 5509
rect 11276 5475 11301 5509
rect 11232 5467 11301 5475
rect 11331 5467 11397 5551
rect 11427 5467 11469 5551
rect 11499 5521 11565 5551
rect 11499 5487 11509 5521
rect 11543 5487 11565 5521
rect 11499 5467 11565 5487
rect 11595 5526 11654 5551
rect 11595 5492 11610 5526
rect 11644 5492 11654 5526
rect 11595 5467 11654 5492
rect 11684 5509 11738 5551
rect 11684 5475 11694 5509
rect 11728 5475 11738 5509
rect 11684 5467 11738 5475
rect 11768 5526 11822 5551
rect 11768 5492 11778 5526
rect 11812 5492 11822 5526
rect 11768 5467 11822 5492
rect 11852 5513 11904 5551
rect 11852 5479 11862 5513
rect 11896 5479 11904 5513
rect 11852 5467 11904 5479
rect 11958 5526 12010 5551
rect 11958 5492 11966 5526
rect 12000 5492 12010 5526
rect 11958 5467 12010 5492
rect 12040 5509 12094 5551
rect 12040 5475 12050 5509
rect 12084 5475 12094 5509
rect 12040 5467 12094 5475
rect 12124 5526 12178 5551
rect 12124 5492 12134 5526
rect 12168 5492 12178 5526
rect 12124 5467 12178 5492
rect 12208 5526 12262 5551
rect 12208 5492 12218 5526
rect 12252 5492 12262 5526
rect 12208 5467 12262 5492
rect 12292 5467 12352 5551
rect 12382 5517 12451 5551
rect 12382 5483 12407 5517
rect 12441 5483 12451 5517
rect 12382 5467 12451 5483
rect 12481 5626 12533 5667
rect 12481 5592 12491 5626
rect 12525 5592 12533 5626
rect 12481 5532 12533 5592
rect 12481 5498 12491 5532
rect 12525 5498 12533 5532
rect 12481 5467 12533 5498
rect 12966 5625 13018 5663
rect 12966 5591 12974 5625
rect 13008 5591 13018 5625
rect 12966 5535 13018 5591
rect 12966 5501 12974 5535
rect 13008 5501 13018 5535
rect 12966 5463 13018 5501
rect 13048 5547 13100 5663
rect 14215 5547 14267 5663
rect 13048 5505 13117 5547
rect 13048 5471 13058 5505
rect 13092 5471 13117 5505
rect 13048 5463 13117 5471
rect 13147 5463 13213 5547
rect 13243 5463 13285 5547
rect 13315 5517 13381 5547
rect 13315 5483 13325 5517
rect 13359 5483 13381 5517
rect 13315 5463 13381 5483
rect 13411 5522 13470 5547
rect 13411 5488 13426 5522
rect 13460 5488 13470 5522
rect 13411 5463 13470 5488
rect 13500 5505 13554 5547
rect 13500 5471 13510 5505
rect 13544 5471 13554 5505
rect 13500 5463 13554 5471
rect 13584 5522 13638 5547
rect 13584 5488 13594 5522
rect 13628 5488 13638 5522
rect 13584 5463 13638 5488
rect 13668 5509 13720 5547
rect 13668 5475 13678 5509
rect 13712 5475 13720 5509
rect 13668 5463 13720 5475
rect 13774 5522 13826 5547
rect 13774 5488 13782 5522
rect 13816 5488 13826 5522
rect 13774 5463 13826 5488
rect 13856 5505 13910 5547
rect 13856 5471 13866 5505
rect 13900 5471 13910 5505
rect 13856 5463 13910 5471
rect 13940 5522 13994 5547
rect 13940 5488 13950 5522
rect 13984 5488 13994 5522
rect 13940 5463 13994 5488
rect 14024 5522 14078 5547
rect 14024 5488 14034 5522
rect 14068 5488 14078 5522
rect 14024 5463 14078 5488
rect 14108 5463 14168 5547
rect 14198 5513 14267 5547
rect 14198 5479 14223 5513
rect 14257 5479 14267 5513
rect 14198 5463 14267 5479
rect 14297 5622 14349 5663
rect 14297 5588 14307 5622
rect 14341 5588 14349 5622
rect 14297 5528 14349 5588
rect 14297 5494 14307 5528
rect 14341 5494 14349 5528
rect 14297 5463 14349 5494
rect 14836 5621 14888 5659
rect 14836 5587 14844 5621
rect 14878 5587 14888 5621
rect 14836 5531 14888 5587
rect 14836 5497 14844 5531
rect 14878 5497 14888 5531
rect 14836 5459 14888 5497
rect 14918 5543 14970 5659
rect 16085 5543 16137 5659
rect 14918 5501 14987 5543
rect 14918 5467 14928 5501
rect 14962 5467 14987 5501
rect 14918 5459 14987 5467
rect 15017 5459 15083 5543
rect 15113 5459 15155 5543
rect 15185 5513 15251 5543
rect 15185 5479 15195 5513
rect 15229 5479 15251 5513
rect 15185 5459 15251 5479
rect 15281 5518 15340 5543
rect 15281 5484 15296 5518
rect 15330 5484 15340 5518
rect 15281 5459 15340 5484
rect 15370 5501 15424 5543
rect 15370 5467 15380 5501
rect 15414 5467 15424 5501
rect 15370 5459 15424 5467
rect 15454 5518 15508 5543
rect 15454 5484 15464 5518
rect 15498 5484 15508 5518
rect 15454 5459 15508 5484
rect 15538 5505 15590 5543
rect 15538 5471 15548 5505
rect 15582 5471 15590 5505
rect 15538 5459 15590 5471
rect 15644 5518 15696 5543
rect 15644 5484 15652 5518
rect 15686 5484 15696 5518
rect 15644 5459 15696 5484
rect 15726 5501 15780 5543
rect 15726 5467 15736 5501
rect 15770 5467 15780 5501
rect 15726 5459 15780 5467
rect 15810 5518 15864 5543
rect 15810 5484 15820 5518
rect 15854 5484 15864 5518
rect 15810 5459 15864 5484
rect 15894 5518 15948 5543
rect 15894 5484 15904 5518
rect 15938 5484 15948 5518
rect 15894 5459 15948 5484
rect 15978 5459 16038 5543
rect 16068 5509 16137 5543
rect 16068 5475 16093 5509
rect 16127 5475 16137 5509
rect 16068 5459 16137 5475
rect 16167 5618 16219 5659
rect 16167 5584 16177 5618
rect 16211 5584 16219 5618
rect 16167 5524 16219 5584
rect 16167 5490 16177 5524
rect 16211 5490 16219 5524
rect 16167 5459 16219 5490
rect 8703 5123 8755 5239
rect 7536 5081 7605 5123
rect 7536 5047 7546 5081
rect 7580 5047 7605 5081
rect 7536 5039 7605 5047
rect 7635 5039 7701 5123
rect 7731 5039 7773 5123
rect 7803 5093 7869 5123
rect 7803 5059 7813 5093
rect 7847 5059 7869 5093
rect 7803 5039 7869 5059
rect 7899 5098 7958 5123
rect 7899 5064 7914 5098
rect 7948 5064 7958 5098
rect 7899 5039 7958 5064
rect 7988 5081 8042 5123
rect 7988 5047 7998 5081
rect 8032 5047 8042 5081
rect 7988 5039 8042 5047
rect 8072 5098 8126 5123
rect 8072 5064 8082 5098
rect 8116 5064 8126 5098
rect 8072 5039 8126 5064
rect 8156 5085 8208 5123
rect 8156 5051 8166 5085
rect 8200 5051 8208 5085
rect 8156 5039 8208 5051
rect 8262 5098 8314 5123
rect 8262 5064 8270 5098
rect 8304 5064 8314 5098
rect 8262 5039 8314 5064
rect 8344 5081 8398 5123
rect 8344 5047 8354 5081
rect 8388 5047 8398 5081
rect 8344 5039 8398 5047
rect 8428 5098 8482 5123
rect 8428 5064 8438 5098
rect 8472 5064 8482 5098
rect 8428 5039 8482 5064
rect 8512 5098 8566 5123
rect 8512 5064 8522 5098
rect 8556 5064 8566 5098
rect 8512 5039 8566 5064
rect 8596 5039 8656 5123
rect 8686 5089 8755 5123
rect 8686 5055 8711 5089
rect 8745 5055 8755 5089
rect 8686 5039 8755 5055
rect 8785 5198 8837 5239
rect 8785 5164 8795 5198
rect 8829 5164 8837 5198
rect 8785 5104 8837 5164
rect 8785 5070 8795 5104
rect 8829 5070 8837 5104
rect 8785 5039 8837 5070
rect 9308 4759 9360 4797
rect 9308 4725 9316 4759
rect 9350 4725 9360 4759
rect 9308 4669 9360 4725
rect 9308 4635 9316 4669
rect 9350 4635 9360 4669
rect 9308 4597 9360 4635
rect 9390 4681 9442 4797
rect 10557 4681 10609 4797
rect 9390 4639 9459 4681
rect 9390 4605 9400 4639
rect 9434 4605 9459 4639
rect 9390 4597 9459 4605
rect 9489 4597 9555 4681
rect 9585 4597 9627 4681
rect 9657 4651 9723 4681
rect 9657 4617 9667 4651
rect 9701 4617 9723 4651
rect 9657 4597 9723 4617
rect 9753 4656 9812 4681
rect 9753 4622 9768 4656
rect 9802 4622 9812 4656
rect 9753 4597 9812 4622
rect 9842 4639 9896 4681
rect 9842 4605 9852 4639
rect 9886 4605 9896 4639
rect 9842 4597 9896 4605
rect 9926 4656 9980 4681
rect 9926 4622 9936 4656
rect 9970 4622 9980 4656
rect 9926 4597 9980 4622
rect 10010 4643 10062 4681
rect 10010 4609 10020 4643
rect 10054 4609 10062 4643
rect 10010 4597 10062 4609
rect 10116 4656 10168 4681
rect 10116 4622 10124 4656
rect 10158 4622 10168 4656
rect 10116 4597 10168 4622
rect 10198 4639 10252 4681
rect 10198 4605 10208 4639
rect 10242 4605 10252 4639
rect 10198 4597 10252 4605
rect 10282 4656 10336 4681
rect 10282 4622 10292 4656
rect 10326 4622 10336 4656
rect 10282 4597 10336 4622
rect 10366 4656 10420 4681
rect 10366 4622 10376 4656
rect 10410 4622 10420 4656
rect 10366 4597 10420 4622
rect 10450 4597 10510 4681
rect 10540 4647 10609 4681
rect 10540 4613 10565 4647
rect 10599 4613 10609 4647
rect 10540 4597 10609 4613
rect 10639 4756 10691 4797
rect 10639 4722 10649 4756
rect 10683 4722 10691 4756
rect 10639 4662 10691 4722
rect 10639 4628 10649 4662
rect 10683 4628 10691 4662
rect 10639 4597 10691 4628
rect 11178 4755 11230 4793
rect 11178 4721 11186 4755
rect 11220 4721 11230 4755
rect 11178 4665 11230 4721
rect 11178 4631 11186 4665
rect 11220 4631 11230 4665
rect 11178 4593 11230 4631
rect 11260 4677 11312 4793
rect 12427 4677 12479 4793
rect 11260 4635 11329 4677
rect 11260 4601 11270 4635
rect 11304 4601 11329 4635
rect 11260 4593 11329 4601
rect 11359 4593 11425 4677
rect 11455 4593 11497 4677
rect 11527 4647 11593 4677
rect 11527 4613 11537 4647
rect 11571 4613 11593 4647
rect 11527 4593 11593 4613
rect 11623 4652 11682 4677
rect 11623 4618 11638 4652
rect 11672 4618 11682 4652
rect 11623 4593 11682 4618
rect 11712 4635 11766 4677
rect 11712 4601 11722 4635
rect 11756 4601 11766 4635
rect 11712 4593 11766 4601
rect 11796 4652 11850 4677
rect 11796 4618 11806 4652
rect 11840 4618 11850 4652
rect 11796 4593 11850 4618
rect 11880 4639 11932 4677
rect 11880 4605 11890 4639
rect 11924 4605 11932 4639
rect 11880 4593 11932 4605
rect 11986 4652 12038 4677
rect 11986 4618 11994 4652
rect 12028 4618 12038 4652
rect 11986 4593 12038 4618
rect 12068 4635 12122 4677
rect 12068 4601 12078 4635
rect 12112 4601 12122 4635
rect 12068 4593 12122 4601
rect 12152 4652 12206 4677
rect 12152 4618 12162 4652
rect 12196 4618 12206 4652
rect 12152 4593 12206 4618
rect 12236 4652 12290 4677
rect 12236 4618 12246 4652
rect 12280 4618 12290 4652
rect 12236 4593 12290 4618
rect 12320 4593 12380 4677
rect 12410 4643 12479 4677
rect 12410 4609 12435 4643
rect 12469 4609 12479 4643
rect 12410 4593 12479 4609
rect 12509 4752 12561 4793
rect 12509 4718 12519 4752
rect 12553 4718 12561 4752
rect 12509 4658 12561 4718
rect 12509 4624 12519 4658
rect 12553 4624 12561 4658
rect 12509 4593 12561 4624
rect 12994 4751 13046 4789
rect 12994 4717 13002 4751
rect 13036 4717 13046 4751
rect 12994 4661 13046 4717
rect 12994 4627 13002 4661
rect 13036 4627 13046 4661
rect 12994 4589 13046 4627
rect 13076 4673 13128 4789
rect 14243 4673 14295 4789
rect 13076 4631 13145 4673
rect 13076 4597 13086 4631
rect 13120 4597 13145 4631
rect 13076 4589 13145 4597
rect 13175 4589 13241 4673
rect 13271 4589 13313 4673
rect 13343 4643 13409 4673
rect 13343 4609 13353 4643
rect 13387 4609 13409 4643
rect 13343 4589 13409 4609
rect 13439 4648 13498 4673
rect 13439 4614 13454 4648
rect 13488 4614 13498 4648
rect 13439 4589 13498 4614
rect 13528 4631 13582 4673
rect 13528 4597 13538 4631
rect 13572 4597 13582 4631
rect 13528 4589 13582 4597
rect 13612 4648 13666 4673
rect 13612 4614 13622 4648
rect 13656 4614 13666 4648
rect 13612 4589 13666 4614
rect 13696 4635 13748 4673
rect 13696 4601 13706 4635
rect 13740 4601 13748 4635
rect 13696 4589 13748 4601
rect 13802 4648 13854 4673
rect 13802 4614 13810 4648
rect 13844 4614 13854 4648
rect 13802 4589 13854 4614
rect 13884 4631 13938 4673
rect 13884 4597 13894 4631
rect 13928 4597 13938 4631
rect 13884 4589 13938 4597
rect 13968 4648 14022 4673
rect 13968 4614 13978 4648
rect 14012 4614 14022 4648
rect 13968 4589 14022 4614
rect 14052 4648 14106 4673
rect 14052 4614 14062 4648
rect 14096 4614 14106 4648
rect 14052 4589 14106 4614
rect 14136 4589 14196 4673
rect 14226 4639 14295 4673
rect 14226 4605 14251 4639
rect 14285 4605 14295 4639
rect 14226 4589 14295 4605
rect 14325 4748 14377 4789
rect 14325 4714 14335 4748
rect 14369 4714 14377 4748
rect 14325 4654 14377 4714
rect 14325 4620 14335 4654
rect 14369 4620 14377 4654
rect 14325 4589 14377 4620
rect 14864 4747 14916 4785
rect 14864 4713 14872 4747
rect 14906 4713 14916 4747
rect 14864 4657 14916 4713
rect 14864 4623 14872 4657
rect 14906 4623 14916 4657
rect 14864 4585 14916 4623
rect 14946 4669 14998 4785
rect 16113 4669 16165 4785
rect 14946 4627 15015 4669
rect 14946 4593 14956 4627
rect 14990 4593 15015 4627
rect 14946 4585 15015 4593
rect 15045 4585 15111 4669
rect 15141 4585 15183 4669
rect 15213 4639 15279 4669
rect 15213 4605 15223 4639
rect 15257 4605 15279 4639
rect 15213 4585 15279 4605
rect 15309 4644 15368 4669
rect 15309 4610 15324 4644
rect 15358 4610 15368 4644
rect 15309 4585 15368 4610
rect 15398 4627 15452 4669
rect 15398 4593 15408 4627
rect 15442 4593 15452 4627
rect 15398 4585 15452 4593
rect 15482 4644 15536 4669
rect 15482 4610 15492 4644
rect 15526 4610 15536 4644
rect 15482 4585 15536 4610
rect 15566 4631 15618 4669
rect 15566 4597 15576 4631
rect 15610 4597 15618 4631
rect 15566 4585 15618 4597
rect 15672 4644 15724 4669
rect 15672 4610 15680 4644
rect 15714 4610 15724 4644
rect 15672 4585 15724 4610
rect 15754 4627 15808 4669
rect 15754 4593 15764 4627
rect 15798 4593 15808 4627
rect 15754 4585 15808 4593
rect 15838 4644 15892 4669
rect 15838 4610 15848 4644
rect 15882 4610 15892 4644
rect 15838 4585 15892 4610
rect 15922 4644 15976 4669
rect 15922 4610 15932 4644
rect 15966 4610 15976 4644
rect 15922 4585 15976 4610
rect 16006 4585 16066 4669
rect 16096 4635 16165 4669
rect 16096 4601 16121 4635
rect 16155 4601 16165 4635
rect 16096 4585 16165 4601
rect 16195 4744 16247 4785
rect 16195 4710 16205 4744
rect 16239 4710 16247 4744
rect 16195 4650 16247 4710
rect 16195 4616 16205 4650
rect 16239 4616 16247 4650
rect 16195 4585 16247 4616
rect 1868 1953 1920 1991
rect 1868 1919 1876 1953
rect 1910 1919 1920 1953
rect 1868 1863 1920 1919
rect 1868 1829 1876 1863
rect 1910 1829 1920 1863
rect 1868 1791 1920 1829
rect 1950 1875 2002 1991
rect 3117 1875 3169 1991
rect 1950 1833 2019 1875
rect 1950 1799 1960 1833
rect 1994 1799 2019 1833
rect 1950 1791 2019 1799
rect 2049 1791 2115 1875
rect 2145 1791 2187 1875
rect 2217 1845 2283 1875
rect 2217 1811 2227 1845
rect 2261 1811 2283 1845
rect 2217 1791 2283 1811
rect 2313 1850 2372 1875
rect 2313 1816 2328 1850
rect 2362 1816 2372 1850
rect 2313 1791 2372 1816
rect 2402 1833 2456 1875
rect 2402 1799 2412 1833
rect 2446 1799 2456 1833
rect 2402 1791 2456 1799
rect 2486 1850 2540 1875
rect 2486 1816 2496 1850
rect 2530 1816 2540 1850
rect 2486 1791 2540 1816
rect 2570 1837 2622 1875
rect 2570 1803 2580 1837
rect 2614 1803 2622 1837
rect 2570 1791 2622 1803
rect 2676 1850 2728 1875
rect 2676 1816 2684 1850
rect 2718 1816 2728 1850
rect 2676 1791 2728 1816
rect 2758 1833 2812 1875
rect 2758 1799 2768 1833
rect 2802 1799 2812 1833
rect 2758 1791 2812 1799
rect 2842 1850 2896 1875
rect 2842 1816 2852 1850
rect 2886 1816 2896 1850
rect 2842 1791 2896 1816
rect 2926 1850 2980 1875
rect 2926 1816 2936 1850
rect 2970 1816 2980 1850
rect 2926 1791 2980 1816
rect 3010 1791 3070 1875
rect 3100 1841 3169 1875
rect 3100 1807 3125 1841
rect 3159 1807 3169 1841
rect 3100 1791 3169 1807
rect 3199 1950 3251 1991
rect 3199 1916 3209 1950
rect 3243 1916 3251 1950
rect 3199 1856 3251 1916
rect 3199 1822 3209 1856
rect 3243 1822 3251 1856
rect 3199 1791 3251 1822
rect 3738 1949 3790 1987
rect 3738 1915 3746 1949
rect 3780 1915 3790 1949
rect 3738 1859 3790 1915
rect 3738 1825 3746 1859
rect 3780 1825 3790 1859
rect 3738 1787 3790 1825
rect 3820 1871 3872 1987
rect 4987 1871 5039 1987
rect 3820 1829 3889 1871
rect 3820 1795 3830 1829
rect 3864 1795 3889 1829
rect 3820 1787 3889 1795
rect 3919 1787 3985 1871
rect 4015 1787 4057 1871
rect 4087 1841 4153 1871
rect 4087 1807 4097 1841
rect 4131 1807 4153 1841
rect 4087 1787 4153 1807
rect 4183 1846 4242 1871
rect 4183 1812 4198 1846
rect 4232 1812 4242 1846
rect 4183 1787 4242 1812
rect 4272 1829 4326 1871
rect 4272 1795 4282 1829
rect 4316 1795 4326 1829
rect 4272 1787 4326 1795
rect 4356 1846 4410 1871
rect 4356 1812 4366 1846
rect 4400 1812 4410 1846
rect 4356 1787 4410 1812
rect 4440 1833 4492 1871
rect 4440 1799 4450 1833
rect 4484 1799 4492 1833
rect 4440 1787 4492 1799
rect 4546 1846 4598 1871
rect 4546 1812 4554 1846
rect 4588 1812 4598 1846
rect 4546 1787 4598 1812
rect 4628 1829 4682 1871
rect 4628 1795 4638 1829
rect 4672 1795 4682 1829
rect 4628 1787 4682 1795
rect 4712 1846 4766 1871
rect 4712 1812 4722 1846
rect 4756 1812 4766 1846
rect 4712 1787 4766 1812
rect 4796 1846 4850 1871
rect 4796 1812 4806 1846
rect 4840 1812 4850 1846
rect 4796 1787 4850 1812
rect 4880 1787 4940 1871
rect 4970 1837 5039 1871
rect 4970 1803 4995 1837
rect 5029 1803 5039 1837
rect 4970 1787 5039 1803
rect 5069 1946 5121 1987
rect 5069 1912 5079 1946
rect 5113 1912 5121 1946
rect 5069 1852 5121 1912
rect 5069 1818 5079 1852
rect 5113 1818 5121 1852
rect 5069 1787 5121 1818
rect 5554 1945 5606 1983
rect 5554 1911 5562 1945
rect 5596 1911 5606 1945
rect 5554 1855 5606 1911
rect 5554 1821 5562 1855
rect 5596 1821 5606 1855
rect 5554 1783 5606 1821
rect 5636 1867 5688 1983
rect 6803 1867 6855 1983
rect 5636 1825 5705 1867
rect 5636 1791 5646 1825
rect 5680 1791 5705 1825
rect 5636 1783 5705 1791
rect 5735 1783 5801 1867
rect 5831 1783 5873 1867
rect 5903 1837 5969 1867
rect 5903 1803 5913 1837
rect 5947 1803 5969 1837
rect 5903 1783 5969 1803
rect 5999 1842 6058 1867
rect 5999 1808 6014 1842
rect 6048 1808 6058 1842
rect 5999 1783 6058 1808
rect 6088 1825 6142 1867
rect 6088 1791 6098 1825
rect 6132 1791 6142 1825
rect 6088 1783 6142 1791
rect 6172 1842 6226 1867
rect 6172 1808 6182 1842
rect 6216 1808 6226 1842
rect 6172 1783 6226 1808
rect 6256 1829 6308 1867
rect 6256 1795 6266 1829
rect 6300 1795 6308 1829
rect 6256 1783 6308 1795
rect 6362 1842 6414 1867
rect 6362 1808 6370 1842
rect 6404 1808 6414 1842
rect 6362 1783 6414 1808
rect 6444 1825 6498 1867
rect 6444 1791 6454 1825
rect 6488 1791 6498 1825
rect 6444 1783 6498 1791
rect 6528 1842 6582 1867
rect 6528 1808 6538 1842
rect 6572 1808 6582 1842
rect 6528 1783 6582 1808
rect 6612 1842 6666 1867
rect 6612 1808 6622 1842
rect 6656 1808 6666 1842
rect 6612 1783 6666 1808
rect 6696 1783 6756 1867
rect 6786 1833 6855 1867
rect 6786 1799 6811 1833
rect 6845 1799 6855 1833
rect 6786 1783 6855 1799
rect 6885 1942 6937 1983
rect 6885 1908 6895 1942
rect 6929 1908 6937 1942
rect 6885 1848 6937 1908
rect 6885 1814 6895 1848
rect 6929 1814 6937 1848
rect 6885 1783 6937 1814
rect 7424 1941 7476 1979
rect 7424 1907 7432 1941
rect 7466 1907 7476 1941
rect 7424 1851 7476 1907
rect 7424 1817 7432 1851
rect 7466 1817 7476 1851
rect 7424 1779 7476 1817
rect 7506 1863 7558 1979
rect 8673 1863 8725 1979
rect 7506 1821 7575 1863
rect 7506 1787 7516 1821
rect 7550 1787 7575 1821
rect 7506 1779 7575 1787
rect 7605 1779 7671 1863
rect 7701 1779 7743 1863
rect 7773 1833 7839 1863
rect 7773 1799 7783 1833
rect 7817 1799 7839 1833
rect 7773 1779 7839 1799
rect 7869 1838 7928 1863
rect 7869 1804 7884 1838
rect 7918 1804 7928 1838
rect 7869 1779 7928 1804
rect 7958 1821 8012 1863
rect 7958 1787 7968 1821
rect 8002 1787 8012 1821
rect 7958 1779 8012 1787
rect 8042 1838 8096 1863
rect 8042 1804 8052 1838
rect 8086 1804 8096 1838
rect 8042 1779 8096 1804
rect 8126 1825 8178 1863
rect 8126 1791 8136 1825
rect 8170 1791 8178 1825
rect 8126 1779 8178 1791
rect 8232 1838 8284 1863
rect 8232 1804 8240 1838
rect 8274 1804 8284 1838
rect 8232 1779 8284 1804
rect 8314 1821 8368 1863
rect 8314 1787 8324 1821
rect 8358 1787 8368 1821
rect 8314 1779 8368 1787
rect 8398 1838 8452 1863
rect 8398 1804 8408 1838
rect 8442 1804 8452 1838
rect 8398 1779 8452 1804
rect 8482 1838 8536 1863
rect 8482 1804 8492 1838
rect 8526 1804 8536 1838
rect 8482 1779 8536 1804
rect 8566 1779 8626 1863
rect 8656 1829 8725 1863
rect 8656 1795 8681 1829
rect 8715 1795 8725 1829
rect 8656 1779 8725 1795
rect 8755 1938 8807 1979
rect 8755 1904 8765 1938
rect 8799 1904 8807 1938
rect 8755 1844 8807 1904
rect 8755 1810 8765 1844
rect 8799 1810 8807 1844
rect 8755 1779 8807 1810
rect 9238 1939 9290 1977
rect 9238 1905 9246 1939
rect 9280 1905 9290 1939
rect 9238 1849 9290 1905
rect 9238 1815 9246 1849
rect 9280 1815 9290 1849
rect 9238 1777 9290 1815
rect 9320 1861 9372 1977
rect 10487 1861 10539 1977
rect 9320 1819 9389 1861
rect 9320 1785 9330 1819
rect 9364 1785 9389 1819
rect 9320 1777 9389 1785
rect 9419 1777 9485 1861
rect 9515 1777 9557 1861
rect 9587 1831 9653 1861
rect 9587 1797 9597 1831
rect 9631 1797 9653 1831
rect 9587 1777 9653 1797
rect 9683 1836 9742 1861
rect 9683 1802 9698 1836
rect 9732 1802 9742 1836
rect 9683 1777 9742 1802
rect 9772 1819 9826 1861
rect 9772 1785 9782 1819
rect 9816 1785 9826 1819
rect 9772 1777 9826 1785
rect 9856 1836 9910 1861
rect 9856 1802 9866 1836
rect 9900 1802 9910 1836
rect 9856 1777 9910 1802
rect 9940 1823 9992 1861
rect 9940 1789 9950 1823
rect 9984 1789 9992 1823
rect 9940 1777 9992 1789
rect 10046 1836 10098 1861
rect 10046 1802 10054 1836
rect 10088 1802 10098 1836
rect 10046 1777 10098 1802
rect 10128 1819 10182 1861
rect 10128 1785 10138 1819
rect 10172 1785 10182 1819
rect 10128 1777 10182 1785
rect 10212 1836 10266 1861
rect 10212 1802 10222 1836
rect 10256 1802 10266 1836
rect 10212 1777 10266 1802
rect 10296 1836 10350 1861
rect 10296 1802 10306 1836
rect 10340 1802 10350 1836
rect 10296 1777 10350 1802
rect 10380 1777 10440 1861
rect 10470 1827 10539 1861
rect 10470 1793 10495 1827
rect 10529 1793 10539 1827
rect 10470 1777 10539 1793
rect 10569 1936 10621 1977
rect 10569 1902 10579 1936
rect 10613 1902 10621 1936
rect 10569 1842 10621 1902
rect 10569 1808 10579 1842
rect 10613 1808 10621 1842
rect 10569 1777 10621 1808
rect 11108 1935 11160 1973
rect 11108 1901 11116 1935
rect 11150 1901 11160 1935
rect 11108 1845 11160 1901
rect 11108 1811 11116 1845
rect 11150 1811 11160 1845
rect 11108 1773 11160 1811
rect 11190 1857 11242 1973
rect 12357 1857 12409 1973
rect 11190 1815 11259 1857
rect 11190 1781 11200 1815
rect 11234 1781 11259 1815
rect 11190 1773 11259 1781
rect 11289 1773 11355 1857
rect 11385 1773 11427 1857
rect 11457 1827 11523 1857
rect 11457 1793 11467 1827
rect 11501 1793 11523 1827
rect 11457 1773 11523 1793
rect 11553 1832 11612 1857
rect 11553 1798 11568 1832
rect 11602 1798 11612 1832
rect 11553 1773 11612 1798
rect 11642 1815 11696 1857
rect 11642 1781 11652 1815
rect 11686 1781 11696 1815
rect 11642 1773 11696 1781
rect 11726 1832 11780 1857
rect 11726 1798 11736 1832
rect 11770 1798 11780 1832
rect 11726 1773 11780 1798
rect 11810 1819 11862 1857
rect 11810 1785 11820 1819
rect 11854 1785 11862 1819
rect 11810 1773 11862 1785
rect 11916 1832 11968 1857
rect 11916 1798 11924 1832
rect 11958 1798 11968 1832
rect 11916 1773 11968 1798
rect 11998 1815 12052 1857
rect 11998 1781 12008 1815
rect 12042 1781 12052 1815
rect 11998 1773 12052 1781
rect 12082 1832 12136 1857
rect 12082 1798 12092 1832
rect 12126 1798 12136 1832
rect 12082 1773 12136 1798
rect 12166 1832 12220 1857
rect 12166 1798 12176 1832
rect 12210 1798 12220 1832
rect 12166 1773 12220 1798
rect 12250 1773 12310 1857
rect 12340 1823 12409 1857
rect 12340 1789 12365 1823
rect 12399 1789 12409 1823
rect 12340 1773 12409 1789
rect 12439 1932 12491 1973
rect 12439 1898 12449 1932
rect 12483 1898 12491 1932
rect 12439 1838 12491 1898
rect 12439 1804 12449 1838
rect 12483 1804 12491 1838
rect 12439 1773 12491 1804
rect 12924 1931 12976 1969
rect 12924 1897 12932 1931
rect 12966 1897 12976 1931
rect 12924 1841 12976 1897
rect 12924 1807 12932 1841
rect 12966 1807 12976 1841
rect 12924 1769 12976 1807
rect 13006 1853 13058 1969
rect 14173 1853 14225 1969
rect 13006 1811 13075 1853
rect 13006 1777 13016 1811
rect 13050 1777 13075 1811
rect 13006 1769 13075 1777
rect 13105 1769 13171 1853
rect 13201 1769 13243 1853
rect 13273 1823 13339 1853
rect 13273 1789 13283 1823
rect 13317 1789 13339 1823
rect 13273 1769 13339 1789
rect 13369 1828 13428 1853
rect 13369 1794 13384 1828
rect 13418 1794 13428 1828
rect 13369 1769 13428 1794
rect 13458 1811 13512 1853
rect 13458 1777 13468 1811
rect 13502 1777 13512 1811
rect 13458 1769 13512 1777
rect 13542 1828 13596 1853
rect 13542 1794 13552 1828
rect 13586 1794 13596 1828
rect 13542 1769 13596 1794
rect 13626 1815 13678 1853
rect 13626 1781 13636 1815
rect 13670 1781 13678 1815
rect 13626 1769 13678 1781
rect 13732 1828 13784 1853
rect 13732 1794 13740 1828
rect 13774 1794 13784 1828
rect 13732 1769 13784 1794
rect 13814 1811 13868 1853
rect 13814 1777 13824 1811
rect 13858 1777 13868 1811
rect 13814 1769 13868 1777
rect 13898 1828 13952 1853
rect 13898 1794 13908 1828
rect 13942 1794 13952 1828
rect 13898 1769 13952 1794
rect 13982 1828 14036 1853
rect 13982 1794 13992 1828
rect 14026 1794 14036 1828
rect 13982 1769 14036 1794
rect 14066 1769 14126 1853
rect 14156 1819 14225 1853
rect 14156 1785 14181 1819
rect 14215 1785 14225 1819
rect 14156 1769 14225 1785
rect 14255 1928 14307 1969
rect 14255 1894 14265 1928
rect 14299 1894 14307 1928
rect 14255 1834 14307 1894
rect 14255 1800 14265 1834
rect 14299 1800 14307 1834
rect 14255 1769 14307 1800
rect 14794 1927 14846 1965
rect 14794 1893 14802 1927
rect 14836 1893 14846 1927
rect 14794 1837 14846 1893
rect 14794 1803 14802 1837
rect 14836 1803 14846 1837
rect 14794 1765 14846 1803
rect 14876 1849 14928 1965
rect 16043 1849 16095 1965
rect 14876 1807 14945 1849
rect 14876 1773 14886 1807
rect 14920 1773 14945 1807
rect 14876 1765 14945 1773
rect 14975 1765 15041 1849
rect 15071 1765 15113 1849
rect 15143 1819 15209 1849
rect 15143 1785 15153 1819
rect 15187 1785 15209 1819
rect 15143 1765 15209 1785
rect 15239 1824 15298 1849
rect 15239 1790 15254 1824
rect 15288 1790 15298 1824
rect 15239 1765 15298 1790
rect 15328 1807 15382 1849
rect 15328 1773 15338 1807
rect 15372 1773 15382 1807
rect 15328 1765 15382 1773
rect 15412 1824 15466 1849
rect 15412 1790 15422 1824
rect 15456 1790 15466 1824
rect 15412 1765 15466 1790
rect 15496 1811 15548 1849
rect 15496 1777 15506 1811
rect 15540 1777 15548 1811
rect 15496 1765 15548 1777
rect 15602 1824 15654 1849
rect 15602 1790 15610 1824
rect 15644 1790 15654 1824
rect 15602 1765 15654 1790
rect 15684 1807 15738 1849
rect 15684 1773 15694 1807
rect 15728 1773 15738 1807
rect 15684 1765 15738 1773
rect 15768 1824 15822 1849
rect 15768 1790 15778 1824
rect 15812 1790 15822 1824
rect 15768 1765 15822 1790
rect 15852 1824 15906 1849
rect 15852 1790 15862 1824
rect 15896 1790 15906 1824
rect 15852 1765 15906 1790
rect 15936 1765 15996 1849
rect 16026 1815 16095 1849
rect 16026 1781 16051 1815
rect 16085 1781 16095 1815
rect 16026 1765 16095 1781
rect 16125 1924 16177 1965
rect 16125 1890 16135 1924
rect 16169 1890 16177 1924
rect 16125 1830 16177 1890
rect 16125 1796 16135 1830
rect 16169 1796 16177 1830
rect 16125 1765 16177 1796
<< ndiffc >>
rect 9473 16087 9507 16121
rect 9557 16109 9591 16143
rect 9641 16087 9675 16121
rect 9809 16089 9843 16123
rect 9909 16089 9943 16123
rect 9999 16160 10033 16194
rect 9999 16092 10033 16126
rect 9599 15369 9633 15403
rect 9791 15341 9825 15375
rect 9875 15341 9909 15375
rect 11605 15239 11639 15273
rect 12046 15299 12080 15333
rect 12046 15231 12080 15265
rect 12145 15299 12179 15333
rect 12145 15231 12179 15265
rect 10783 14759 10817 14793
rect 10975 14731 11009 14765
rect 11059 14731 11093 14765
rect 9483 14523 9517 14557
rect 9567 14545 9601 14579
rect 9651 14523 9685 14557
rect 9819 14525 9853 14559
rect 9919 14525 9953 14559
rect 10009 14596 10043 14630
rect 10009 14528 10043 14562
rect 9609 13805 9643 13839
rect 9801 13777 9835 13811
rect 9885 13777 9919 13811
rect 10821 13773 10855 13807
rect 11262 13833 11296 13867
rect 11262 13765 11296 13799
rect 11361 13833 11395 13867
rect 11361 13765 11395 13799
rect 12639 13773 12673 13807
rect 12729 13767 12763 13801
rect 12819 13753 12853 13787
rect 12903 13767 12937 13801
rect 12997 13753 13031 13787
rect 13085 13791 13119 13825
rect 11820 13401 11854 13435
rect 11904 13401 11938 13435
rect 12000 13401 12034 13435
rect 12085 13461 12119 13495
rect 12085 13393 12119 13427
rect 9475 12855 9509 12889
rect 9559 12877 9593 12911
rect 9643 12855 9677 12889
rect 9811 12857 9845 12891
rect 9911 12857 9945 12891
rect 10001 12928 10035 12962
rect 10945 12923 10979 12957
rect 11217 12939 11251 12973
rect 11301 12949 11335 12983
rect 10001 12860 10035 12894
rect 9601 12137 9635 12171
rect 9793 12109 9827 12143
rect 9877 12109 9911 12143
rect 10977 11931 11011 11965
rect 11169 11903 11203 11937
rect 11253 11903 11287 11937
rect 9485 11291 9519 11325
rect 9569 11313 9603 11347
rect 9653 11291 9687 11325
rect 9821 11293 9855 11327
rect 9921 11293 9955 11327
rect 10011 11364 10045 11398
rect 10011 11296 10045 11330
rect 9611 10573 9645 10607
rect 9803 10545 9837 10579
rect 9887 10545 9921 10579
rect 6194 6503 6228 6537
rect 6194 6435 6228 6469
rect 6278 6503 6312 6537
rect 6278 6435 6312 6469
rect 9288 5839 9322 5873
rect 9387 5879 9421 5913
rect 9639 5867 9673 5901
rect 9740 5862 9774 5896
rect 9824 5879 9858 5913
rect 9908 5862 9942 5896
rect 9992 5870 10026 5904
rect 10096 5862 10130 5896
rect 10180 5879 10214 5913
rect 10264 5862 10298 5896
rect 10348 5862 10382 5896
rect 10537 5875 10571 5909
rect 1906 5419 1940 5453
rect 2005 5459 2039 5493
rect 2257 5447 2291 5481
rect 2358 5442 2392 5476
rect 2442 5459 2476 5493
rect 2526 5442 2560 5476
rect 2610 5450 2644 5484
rect 2714 5442 2748 5476
rect 2798 5459 2832 5493
rect 2882 5442 2916 5476
rect 2966 5442 3000 5476
rect 3155 5455 3189 5489
rect 3239 5419 3273 5453
rect 3776 5415 3810 5449
rect 3875 5455 3909 5489
rect 4127 5443 4161 5477
rect 4228 5438 4262 5472
rect 4312 5455 4346 5489
rect 4396 5438 4430 5472
rect 4480 5446 4514 5480
rect 4584 5438 4618 5472
rect 4668 5455 4702 5489
rect 4752 5438 4786 5472
rect 4836 5438 4870 5472
rect 5025 5451 5059 5485
rect 5109 5415 5143 5449
rect 5592 5411 5626 5445
rect 5691 5451 5725 5485
rect 5943 5439 5977 5473
rect 6044 5434 6078 5468
rect 6128 5451 6162 5485
rect 6212 5434 6246 5468
rect 6296 5442 6330 5476
rect 6400 5434 6434 5468
rect 6484 5451 6518 5485
rect 6568 5434 6602 5468
rect 6652 5434 6686 5468
rect 6841 5447 6875 5481
rect 6925 5411 6959 5445
rect 7462 5407 7496 5441
rect 7561 5447 7595 5481
rect 7813 5435 7847 5469
rect 7914 5430 7948 5464
rect 7998 5447 8032 5481
rect 8082 5430 8116 5464
rect 8166 5438 8200 5472
rect 8270 5430 8304 5464
rect 8354 5447 8388 5481
rect 8438 5430 8472 5464
rect 8522 5430 8556 5464
rect 8711 5443 8745 5477
rect 10621 5839 10655 5873
rect 11158 5835 11192 5869
rect 11257 5875 11291 5909
rect 11509 5863 11543 5897
rect 11610 5858 11644 5892
rect 11694 5875 11728 5909
rect 11778 5858 11812 5892
rect 11862 5866 11896 5900
rect 11966 5858 12000 5892
rect 12050 5875 12084 5909
rect 12134 5858 12168 5892
rect 12218 5858 12252 5892
rect 12407 5871 12441 5905
rect 12491 5835 12525 5869
rect 12974 5831 13008 5865
rect 13073 5871 13107 5905
rect 13325 5859 13359 5893
rect 13426 5854 13460 5888
rect 13510 5871 13544 5905
rect 13594 5854 13628 5888
rect 13678 5862 13712 5896
rect 13782 5854 13816 5888
rect 13866 5871 13900 5905
rect 13950 5854 13984 5888
rect 14034 5854 14068 5888
rect 14223 5867 14257 5901
rect 14307 5831 14341 5865
rect 14844 5827 14878 5861
rect 14943 5867 14977 5901
rect 15195 5855 15229 5889
rect 15296 5850 15330 5884
rect 15380 5867 15414 5901
rect 15464 5850 15498 5884
rect 15548 5858 15582 5892
rect 15652 5850 15686 5884
rect 15736 5867 15770 5901
rect 15820 5850 15854 5884
rect 15904 5850 15938 5884
rect 16093 5863 16127 5897
rect 8795 5407 8829 5441
rect 16177 5827 16211 5861
rect 9316 4965 9350 4999
rect 9415 5005 9449 5039
rect 9667 4993 9701 5027
rect 9768 4988 9802 5022
rect 9852 5005 9886 5039
rect 9936 4988 9970 5022
rect 10020 4996 10054 5030
rect 10124 4988 10158 5022
rect 10208 5005 10242 5039
rect 10292 4988 10326 5022
rect 10376 4988 10410 5022
rect 10565 5001 10599 5035
rect 10649 4965 10683 4999
rect 11186 4961 11220 4995
rect 11285 5001 11319 5035
rect 11537 4989 11571 5023
rect 11638 4984 11672 5018
rect 11722 5001 11756 5035
rect 11806 4984 11840 5018
rect 11890 4992 11924 5026
rect 11994 4984 12028 5018
rect 12078 5001 12112 5035
rect 12162 4984 12196 5018
rect 12246 4984 12280 5018
rect 12435 4997 12469 5031
rect 12519 4961 12553 4995
rect 13002 4957 13036 4991
rect 13101 4997 13135 5031
rect 13353 4985 13387 5019
rect 13454 4980 13488 5014
rect 13538 4997 13572 5031
rect 13622 4980 13656 5014
rect 13706 4988 13740 5022
rect 13810 4980 13844 5014
rect 13894 4997 13928 5031
rect 13978 4980 14012 5014
rect 14062 4980 14096 5014
rect 14251 4993 14285 5027
rect 14335 4957 14369 4991
rect 14872 4953 14906 4987
rect 14971 4993 15005 5027
rect 15223 4981 15257 5015
rect 15324 4976 15358 5010
rect 15408 4993 15442 5027
rect 15492 4976 15526 5010
rect 15576 4984 15610 5018
rect 15680 4976 15714 5010
rect 15764 4993 15798 5027
rect 15848 4976 15882 5010
rect 15932 4976 15966 5010
rect 16121 4989 16155 5023
rect 16205 4953 16239 4987
rect 1876 2159 1910 2193
rect 1975 2199 2009 2233
rect 2227 2187 2261 2221
rect 2328 2182 2362 2216
rect 2412 2199 2446 2233
rect 2496 2182 2530 2216
rect 2580 2190 2614 2224
rect 2684 2182 2718 2216
rect 2768 2199 2802 2233
rect 2852 2182 2886 2216
rect 2936 2182 2970 2216
rect 3125 2195 3159 2229
rect 3209 2159 3243 2193
rect 3746 2155 3780 2189
rect 3845 2195 3879 2229
rect 4097 2183 4131 2217
rect 4198 2178 4232 2212
rect 4282 2195 4316 2229
rect 4366 2178 4400 2212
rect 4450 2186 4484 2220
rect 4554 2178 4588 2212
rect 4638 2195 4672 2229
rect 4722 2178 4756 2212
rect 4806 2178 4840 2212
rect 4995 2191 5029 2225
rect 5079 2155 5113 2189
rect 5562 2151 5596 2185
rect 5661 2191 5695 2225
rect 5913 2179 5947 2213
rect 6014 2174 6048 2208
rect 6098 2191 6132 2225
rect 6182 2174 6216 2208
rect 6266 2182 6300 2216
rect 6370 2174 6404 2208
rect 6454 2191 6488 2225
rect 6538 2174 6572 2208
rect 6622 2174 6656 2208
rect 6811 2187 6845 2221
rect 6895 2151 6929 2185
rect 7432 2147 7466 2181
rect 7531 2187 7565 2221
rect 7783 2175 7817 2209
rect 7884 2170 7918 2204
rect 7968 2187 8002 2221
rect 8052 2170 8086 2204
rect 8136 2178 8170 2212
rect 8240 2170 8274 2204
rect 8324 2187 8358 2221
rect 8408 2170 8442 2204
rect 8492 2170 8526 2204
rect 8681 2183 8715 2217
rect 8765 2147 8799 2181
rect 9246 2145 9280 2179
rect 9345 2185 9379 2219
rect 9597 2173 9631 2207
rect 9698 2168 9732 2202
rect 9782 2185 9816 2219
rect 9866 2168 9900 2202
rect 9950 2176 9984 2210
rect 10054 2168 10088 2202
rect 10138 2185 10172 2219
rect 10222 2168 10256 2202
rect 10306 2168 10340 2202
rect 10495 2181 10529 2215
rect 10579 2145 10613 2179
rect 11116 2141 11150 2175
rect 11215 2181 11249 2215
rect 11467 2169 11501 2203
rect 11568 2164 11602 2198
rect 11652 2181 11686 2215
rect 11736 2164 11770 2198
rect 11820 2172 11854 2206
rect 11924 2164 11958 2198
rect 12008 2181 12042 2215
rect 12092 2164 12126 2198
rect 12176 2164 12210 2198
rect 12365 2177 12399 2211
rect 12449 2141 12483 2175
rect 12932 2137 12966 2171
rect 13031 2177 13065 2211
rect 13283 2165 13317 2199
rect 13384 2160 13418 2194
rect 13468 2177 13502 2211
rect 13552 2160 13586 2194
rect 13636 2168 13670 2202
rect 13740 2160 13774 2194
rect 13824 2177 13858 2211
rect 13908 2160 13942 2194
rect 13992 2160 14026 2194
rect 14181 2173 14215 2207
rect 14265 2137 14299 2171
rect 14802 2133 14836 2167
rect 14901 2173 14935 2207
rect 15153 2161 15187 2195
rect 15254 2156 15288 2190
rect 15338 2173 15372 2207
rect 15422 2156 15456 2190
rect 15506 2164 15540 2198
rect 15610 2156 15644 2190
rect 15694 2173 15728 2207
rect 15778 2156 15812 2190
rect 15862 2156 15896 2190
rect 16051 2169 16085 2203
rect 16135 2133 16169 2167
<< pdiffc >>
rect 9473 16477 9507 16511
rect 9473 16409 9507 16443
rect 9641 16467 9675 16501
rect 9641 16399 9675 16433
rect 9725 16467 9759 16501
rect 9725 16399 9759 16433
rect 9809 16467 9843 16501
rect 9913 16467 9947 16501
rect 9913 16399 9947 16433
rect 9997 16469 10031 16503
rect 9997 16401 10031 16435
rect 9997 16333 10031 16367
rect 9599 15691 9633 15725
rect 9683 15691 9717 15725
rect 9791 15733 9825 15767
rect 9791 15665 9825 15699
rect 9895 15733 9929 15767
rect 9895 15665 9929 15699
rect 11605 15623 11639 15657
rect 11697 15615 11731 15649
rect 11799 15623 11833 15657
rect 11894 15615 11928 15649
rect 12045 15623 12079 15657
rect 12045 15555 12079 15589
rect 12145 15623 12179 15657
rect 12145 15555 12179 15589
rect 12145 15487 12179 15521
rect 10783 15081 10817 15115
rect 10867 15081 10901 15115
rect 10975 15123 11009 15157
rect 10975 15055 11009 15089
rect 9483 14913 9517 14947
rect 9483 14845 9517 14879
rect 9651 14903 9685 14937
rect 9651 14835 9685 14869
rect 9735 14903 9769 14937
rect 9735 14835 9769 14869
rect 9819 14903 9853 14937
rect 9923 14903 9957 14937
rect 9923 14835 9957 14869
rect 10007 14905 10041 14939
rect 10007 14837 10041 14871
rect 11079 15123 11113 15157
rect 11079 15055 11113 15089
rect 10007 14769 10041 14803
rect 9609 14127 9643 14161
rect 9693 14127 9727 14161
rect 9801 14169 9835 14203
rect 9801 14101 9835 14135
rect 9905 14169 9939 14203
rect 9905 14101 9939 14135
rect 10821 14157 10855 14191
rect 10913 14149 10947 14183
rect 11015 14157 11049 14191
rect 11110 14149 11144 14183
rect 11261 14157 11295 14191
rect 11261 14089 11295 14123
rect 11361 14157 11395 14191
rect 11361 14089 11395 14123
rect 13000 14141 13034 14175
rect 13000 14073 13034 14107
rect 11361 14021 11395 14055
rect 12639 14010 12673 14044
rect 13085 14110 13119 14144
rect 13085 14042 13119 14076
rect 12001 13767 12035 13801
rect 11832 13647 11866 13681
rect 12001 13699 12035 13733
rect 12101 13783 12135 13817
rect 12101 13715 12135 13749
rect 9475 13245 9509 13279
rect 9475 13177 9509 13211
rect 9643 13235 9677 13269
rect 9643 13167 9677 13201
rect 9727 13235 9761 13269
rect 9727 13167 9761 13201
rect 9811 13235 9845 13269
rect 9915 13235 9949 13269
rect 9915 13167 9949 13201
rect 11217 13315 11251 13349
rect 9999 13237 10033 13271
rect 9999 13169 10033 13203
rect 10945 13176 10979 13210
rect 11029 13206 11063 13240
rect 11122 13187 11156 13221
rect 9999 13101 10033 13135
rect 11301 13301 11335 13335
rect 11301 13233 11335 13267
rect 9601 12459 9635 12493
rect 9685 12459 9719 12493
rect 9793 12501 9827 12535
rect 9793 12433 9827 12467
rect 9897 12501 9931 12535
rect 9897 12433 9931 12467
rect 10977 12253 11011 12287
rect 11061 12253 11095 12287
rect 11169 12295 11203 12329
rect 11169 12227 11203 12261
rect 11273 12295 11307 12329
rect 11273 12227 11307 12261
rect 9485 11681 9519 11715
rect 9485 11613 9519 11647
rect 9653 11671 9687 11705
rect 9653 11603 9687 11637
rect 9737 11671 9771 11705
rect 9737 11603 9771 11637
rect 9821 11671 9855 11705
rect 9925 11671 9959 11705
rect 9925 11603 9959 11637
rect 10009 11673 10043 11707
rect 10009 11605 10043 11639
rect 10009 11537 10043 11571
rect 9611 10895 9645 10929
rect 9695 10895 9729 10929
rect 9803 10937 9837 10971
rect 9803 10869 9837 10903
rect 9907 10937 9941 10971
rect 9907 10869 9941 10903
rect 6194 6251 6228 6285
rect 6194 6183 6228 6217
rect 6194 6115 6228 6149
rect 6278 6251 6312 6285
rect 6278 6183 6312 6217
rect 6278 6115 6312 6149
rect 9288 5599 9322 5633
rect 1906 5179 1940 5213
rect 1906 5089 1940 5123
rect 1990 5059 2024 5093
rect 2257 5071 2291 5105
rect 2358 5076 2392 5110
rect 2442 5059 2476 5093
rect 2526 5076 2560 5110
rect 2610 5063 2644 5097
rect 2714 5076 2748 5110
rect 2798 5059 2832 5093
rect 2882 5076 2916 5110
rect 2966 5076 3000 5110
rect 3155 5067 3189 5101
rect 3239 5176 3273 5210
rect 3239 5082 3273 5116
rect 3776 5175 3810 5209
rect 3776 5085 3810 5119
rect 3860 5055 3894 5089
rect 4127 5067 4161 5101
rect 4228 5072 4262 5106
rect 4312 5055 4346 5089
rect 4396 5072 4430 5106
rect 4480 5059 4514 5093
rect 4584 5072 4618 5106
rect 4668 5055 4702 5089
rect 4752 5072 4786 5106
rect 4836 5072 4870 5106
rect 5025 5063 5059 5097
rect 5109 5172 5143 5206
rect 5109 5078 5143 5112
rect 5592 5171 5626 5205
rect 5592 5081 5626 5115
rect 9288 5509 9322 5543
rect 5676 5051 5710 5085
rect 5943 5063 5977 5097
rect 6044 5068 6078 5102
rect 6128 5051 6162 5085
rect 6212 5068 6246 5102
rect 6296 5055 6330 5089
rect 6400 5068 6434 5102
rect 6484 5051 6518 5085
rect 6568 5068 6602 5102
rect 6652 5068 6686 5102
rect 6841 5059 6875 5093
rect 6925 5168 6959 5202
rect 6925 5074 6959 5108
rect 7462 5167 7496 5201
rect 7462 5077 7496 5111
rect 9372 5479 9406 5513
rect 9639 5491 9673 5525
rect 9740 5496 9774 5530
rect 9824 5479 9858 5513
rect 9908 5496 9942 5530
rect 9992 5483 10026 5517
rect 10096 5496 10130 5530
rect 10180 5479 10214 5513
rect 10264 5496 10298 5530
rect 10348 5496 10382 5530
rect 10537 5487 10571 5521
rect 10621 5596 10655 5630
rect 10621 5502 10655 5536
rect 11158 5595 11192 5629
rect 11158 5505 11192 5539
rect 11242 5475 11276 5509
rect 11509 5487 11543 5521
rect 11610 5492 11644 5526
rect 11694 5475 11728 5509
rect 11778 5492 11812 5526
rect 11862 5479 11896 5513
rect 11966 5492 12000 5526
rect 12050 5475 12084 5509
rect 12134 5492 12168 5526
rect 12218 5492 12252 5526
rect 12407 5483 12441 5517
rect 12491 5592 12525 5626
rect 12491 5498 12525 5532
rect 12974 5591 13008 5625
rect 12974 5501 13008 5535
rect 13058 5471 13092 5505
rect 13325 5483 13359 5517
rect 13426 5488 13460 5522
rect 13510 5471 13544 5505
rect 13594 5488 13628 5522
rect 13678 5475 13712 5509
rect 13782 5488 13816 5522
rect 13866 5471 13900 5505
rect 13950 5488 13984 5522
rect 14034 5488 14068 5522
rect 14223 5479 14257 5513
rect 14307 5588 14341 5622
rect 14307 5494 14341 5528
rect 14844 5587 14878 5621
rect 14844 5497 14878 5531
rect 14928 5467 14962 5501
rect 15195 5479 15229 5513
rect 15296 5484 15330 5518
rect 15380 5467 15414 5501
rect 15464 5484 15498 5518
rect 15548 5471 15582 5505
rect 15652 5484 15686 5518
rect 15736 5467 15770 5501
rect 15820 5484 15854 5518
rect 15904 5484 15938 5518
rect 16093 5475 16127 5509
rect 16177 5584 16211 5618
rect 16177 5490 16211 5524
rect 7546 5047 7580 5081
rect 7813 5059 7847 5093
rect 7914 5064 7948 5098
rect 7998 5047 8032 5081
rect 8082 5064 8116 5098
rect 8166 5051 8200 5085
rect 8270 5064 8304 5098
rect 8354 5047 8388 5081
rect 8438 5064 8472 5098
rect 8522 5064 8556 5098
rect 8711 5055 8745 5089
rect 8795 5164 8829 5198
rect 8795 5070 8829 5104
rect 9316 4725 9350 4759
rect 9316 4635 9350 4669
rect 9400 4605 9434 4639
rect 9667 4617 9701 4651
rect 9768 4622 9802 4656
rect 9852 4605 9886 4639
rect 9936 4622 9970 4656
rect 10020 4609 10054 4643
rect 10124 4622 10158 4656
rect 10208 4605 10242 4639
rect 10292 4622 10326 4656
rect 10376 4622 10410 4656
rect 10565 4613 10599 4647
rect 10649 4722 10683 4756
rect 10649 4628 10683 4662
rect 11186 4721 11220 4755
rect 11186 4631 11220 4665
rect 11270 4601 11304 4635
rect 11537 4613 11571 4647
rect 11638 4618 11672 4652
rect 11722 4601 11756 4635
rect 11806 4618 11840 4652
rect 11890 4605 11924 4639
rect 11994 4618 12028 4652
rect 12078 4601 12112 4635
rect 12162 4618 12196 4652
rect 12246 4618 12280 4652
rect 12435 4609 12469 4643
rect 12519 4718 12553 4752
rect 12519 4624 12553 4658
rect 13002 4717 13036 4751
rect 13002 4627 13036 4661
rect 13086 4597 13120 4631
rect 13353 4609 13387 4643
rect 13454 4614 13488 4648
rect 13538 4597 13572 4631
rect 13622 4614 13656 4648
rect 13706 4601 13740 4635
rect 13810 4614 13844 4648
rect 13894 4597 13928 4631
rect 13978 4614 14012 4648
rect 14062 4614 14096 4648
rect 14251 4605 14285 4639
rect 14335 4714 14369 4748
rect 14335 4620 14369 4654
rect 14872 4713 14906 4747
rect 14872 4623 14906 4657
rect 14956 4593 14990 4627
rect 15223 4605 15257 4639
rect 15324 4610 15358 4644
rect 15408 4593 15442 4627
rect 15492 4610 15526 4644
rect 15576 4597 15610 4631
rect 15680 4610 15714 4644
rect 15764 4593 15798 4627
rect 15848 4610 15882 4644
rect 15932 4610 15966 4644
rect 16121 4601 16155 4635
rect 16205 4710 16239 4744
rect 16205 4616 16239 4650
rect 1876 1919 1910 1953
rect 1876 1829 1910 1863
rect 1960 1799 1994 1833
rect 2227 1811 2261 1845
rect 2328 1816 2362 1850
rect 2412 1799 2446 1833
rect 2496 1816 2530 1850
rect 2580 1803 2614 1837
rect 2684 1816 2718 1850
rect 2768 1799 2802 1833
rect 2852 1816 2886 1850
rect 2936 1816 2970 1850
rect 3125 1807 3159 1841
rect 3209 1916 3243 1950
rect 3209 1822 3243 1856
rect 3746 1915 3780 1949
rect 3746 1825 3780 1859
rect 3830 1795 3864 1829
rect 4097 1807 4131 1841
rect 4198 1812 4232 1846
rect 4282 1795 4316 1829
rect 4366 1812 4400 1846
rect 4450 1799 4484 1833
rect 4554 1812 4588 1846
rect 4638 1795 4672 1829
rect 4722 1812 4756 1846
rect 4806 1812 4840 1846
rect 4995 1803 5029 1837
rect 5079 1912 5113 1946
rect 5079 1818 5113 1852
rect 5562 1911 5596 1945
rect 5562 1821 5596 1855
rect 5646 1791 5680 1825
rect 5913 1803 5947 1837
rect 6014 1808 6048 1842
rect 6098 1791 6132 1825
rect 6182 1808 6216 1842
rect 6266 1795 6300 1829
rect 6370 1808 6404 1842
rect 6454 1791 6488 1825
rect 6538 1808 6572 1842
rect 6622 1808 6656 1842
rect 6811 1799 6845 1833
rect 6895 1908 6929 1942
rect 6895 1814 6929 1848
rect 7432 1907 7466 1941
rect 7432 1817 7466 1851
rect 7516 1787 7550 1821
rect 7783 1799 7817 1833
rect 7884 1804 7918 1838
rect 7968 1787 8002 1821
rect 8052 1804 8086 1838
rect 8136 1791 8170 1825
rect 8240 1804 8274 1838
rect 8324 1787 8358 1821
rect 8408 1804 8442 1838
rect 8492 1804 8526 1838
rect 8681 1795 8715 1829
rect 8765 1904 8799 1938
rect 8765 1810 8799 1844
rect 9246 1905 9280 1939
rect 9246 1815 9280 1849
rect 9330 1785 9364 1819
rect 9597 1797 9631 1831
rect 9698 1802 9732 1836
rect 9782 1785 9816 1819
rect 9866 1802 9900 1836
rect 9950 1789 9984 1823
rect 10054 1802 10088 1836
rect 10138 1785 10172 1819
rect 10222 1802 10256 1836
rect 10306 1802 10340 1836
rect 10495 1793 10529 1827
rect 10579 1902 10613 1936
rect 10579 1808 10613 1842
rect 11116 1901 11150 1935
rect 11116 1811 11150 1845
rect 11200 1781 11234 1815
rect 11467 1793 11501 1827
rect 11568 1798 11602 1832
rect 11652 1781 11686 1815
rect 11736 1798 11770 1832
rect 11820 1785 11854 1819
rect 11924 1798 11958 1832
rect 12008 1781 12042 1815
rect 12092 1798 12126 1832
rect 12176 1798 12210 1832
rect 12365 1789 12399 1823
rect 12449 1898 12483 1932
rect 12449 1804 12483 1838
rect 12932 1897 12966 1931
rect 12932 1807 12966 1841
rect 13016 1777 13050 1811
rect 13283 1789 13317 1823
rect 13384 1794 13418 1828
rect 13468 1777 13502 1811
rect 13552 1794 13586 1828
rect 13636 1781 13670 1815
rect 13740 1794 13774 1828
rect 13824 1777 13858 1811
rect 13908 1794 13942 1828
rect 13992 1794 14026 1828
rect 14181 1785 14215 1819
rect 14265 1894 14299 1928
rect 14265 1800 14299 1834
rect 14802 1893 14836 1927
rect 14802 1803 14836 1837
rect 14886 1773 14920 1807
rect 15153 1785 15187 1819
rect 15254 1790 15288 1824
rect 15338 1773 15372 1807
rect 15422 1790 15456 1824
rect 15506 1777 15540 1811
rect 15610 1790 15644 1824
rect 15694 1773 15728 1807
rect 15778 1790 15812 1824
rect 15862 1790 15896 1824
rect 16051 1781 16085 1815
rect 16135 1890 16169 1924
rect 16135 1796 16169 1830
<< poly >>
rect 9517 16523 9547 16549
rect 9601 16523 9631 16549
rect 9685 16523 9715 16549
rect 9769 16523 9799 16549
rect 9957 16523 9987 16549
rect 9517 16291 9547 16323
rect 9601 16291 9631 16323
rect 9685 16291 9715 16323
rect 9769 16291 9799 16323
rect 9957 16291 9987 16323
rect 9505 16275 9559 16291
rect 9505 16241 9515 16275
rect 9549 16241 9559 16275
rect 9505 16225 9559 16241
rect 9601 16275 9715 16291
rect 9601 16241 9632 16275
rect 9666 16241 9715 16275
rect 9601 16225 9715 16241
rect 9757 16275 9811 16291
rect 9757 16241 9767 16275
rect 9801 16241 9811 16275
rect 9757 16225 9811 16241
rect 9853 16275 9987 16291
rect 9853 16241 9863 16275
rect 9897 16258 9987 16275
rect 9897 16241 9983 16258
rect 9853 16225 9983 16241
rect 9517 16203 9547 16225
rect 9601 16203 9631 16225
rect 9685 16203 9715 16225
rect 9769 16203 9799 16225
rect 9953 16203 9983 16225
rect 9517 16047 9547 16073
rect 9601 16047 9631 16073
rect 9685 16047 9715 16073
rect 9769 16047 9799 16073
rect 9953 16047 9983 16073
rect 9835 15779 9865 15805
rect 9643 15737 9673 15763
rect 9727 15737 9757 15763
rect 9643 15547 9673 15653
rect 9586 15531 9673 15547
rect 9586 15497 9602 15531
rect 9636 15497 9673 15531
rect 9586 15481 9673 15497
rect 9643 15441 9673 15481
rect 9727 15547 9757 15653
rect 11649 15669 11679 15695
rect 11749 15669 11779 15695
rect 11853 15669 11883 15695
rect 11939 15669 11969 15695
rect 12105 15669 12135 15695
rect 9835 15547 9865 15579
rect 9727 15531 9793 15547
rect 9727 15497 9743 15531
rect 9777 15497 9793 15531
rect 9727 15481 9793 15497
rect 9835 15531 9901 15547
rect 9835 15497 9851 15531
rect 9885 15497 9901 15531
rect 9835 15481 9901 15497
rect 9727 15441 9757 15481
rect 9835 15459 9865 15481
rect 9643 15331 9673 15357
rect 9727 15331 9757 15357
rect 11649 15437 11679 15585
rect 11749 15437 11779 15585
rect 11853 15437 11883 15585
rect 11939 15437 11969 15585
rect 12105 15437 12135 15469
rect 11591 15421 11679 15437
rect 11591 15387 11601 15421
rect 11635 15387 11679 15421
rect 11591 15371 11679 15387
rect 9835 15303 9865 15329
rect 11649 15303 11679 15371
rect 11737 15421 11791 15437
rect 11737 15387 11747 15421
rect 11781 15387 11791 15421
rect 11737 15371 11791 15387
rect 11843 15421 11897 15437
rect 11843 15387 11853 15421
rect 11887 15387 11897 15421
rect 11843 15371 11897 15387
rect 11939 15421 12003 15437
rect 11939 15387 11949 15421
rect 11983 15387 12003 15421
rect 11939 15371 12003 15387
rect 12050 15421 12135 15437
rect 12050 15387 12060 15421
rect 12094 15387 12135 15421
rect 12050 15371 12135 15387
rect 11737 15303 11767 15371
rect 11843 15303 11873 15371
rect 11939 15303 11969 15371
rect 12105 15349 12135 15371
rect 11019 15169 11049 15195
rect 11649 15193 11679 15219
rect 11737 15193 11767 15219
rect 11843 15193 11873 15219
rect 11939 15193 11969 15219
rect 12105 15193 12135 15219
rect 10827 15127 10857 15153
rect 10911 15127 10941 15153
rect 9527 14959 9557 14985
rect 9611 14959 9641 14985
rect 9695 14959 9725 14985
rect 9779 14959 9809 14985
rect 9967 14959 9997 14985
rect 10827 14937 10857 15043
rect 10770 14921 10857 14937
rect 10770 14887 10786 14921
rect 10820 14887 10857 14921
rect 10770 14871 10857 14887
rect 10827 14831 10857 14871
rect 10911 14937 10941 15043
rect 11019 14937 11049 14969
rect 10911 14921 10977 14937
rect 10911 14887 10927 14921
rect 10961 14887 10977 14921
rect 10911 14871 10977 14887
rect 11019 14921 11085 14937
rect 11019 14887 11035 14921
rect 11069 14887 11085 14921
rect 11019 14871 11085 14887
rect 10911 14831 10941 14871
rect 11019 14849 11049 14871
rect 9527 14727 9557 14759
rect 9611 14727 9641 14759
rect 9695 14727 9725 14759
rect 9779 14727 9809 14759
rect 9967 14727 9997 14759
rect 9515 14711 9569 14727
rect 9515 14677 9525 14711
rect 9559 14677 9569 14711
rect 9515 14661 9569 14677
rect 9611 14711 9725 14727
rect 9611 14677 9642 14711
rect 9676 14677 9725 14711
rect 9611 14661 9725 14677
rect 9767 14711 9821 14727
rect 9767 14677 9777 14711
rect 9811 14677 9821 14711
rect 9767 14661 9821 14677
rect 9863 14711 9997 14727
rect 10827 14721 10857 14747
rect 10911 14721 10941 14747
rect 9863 14677 9873 14711
rect 9907 14694 9997 14711
rect 9907 14677 9993 14694
rect 11019 14693 11049 14719
rect 9863 14661 9993 14677
rect 9527 14639 9557 14661
rect 9611 14639 9641 14661
rect 9695 14639 9725 14661
rect 9779 14639 9809 14661
rect 9963 14639 9993 14661
rect 9527 14483 9557 14509
rect 9611 14483 9641 14509
rect 9695 14483 9725 14509
rect 9779 14483 9809 14509
rect 9963 14483 9993 14509
rect 9845 14215 9875 14241
rect 9653 14173 9683 14199
rect 9737 14173 9767 14199
rect 9653 13983 9683 14089
rect 9596 13967 9683 13983
rect 9596 13933 9612 13967
rect 9646 13933 9683 13967
rect 9596 13917 9683 13933
rect 9653 13877 9683 13917
rect 9737 13983 9767 14089
rect 10865 14203 10895 14229
rect 10965 14203 10995 14229
rect 11069 14203 11099 14229
rect 11155 14203 11185 14229
rect 11321 14203 11351 14229
rect 9845 13983 9875 14015
rect 9737 13967 9803 13983
rect 9737 13933 9753 13967
rect 9787 13933 9803 13967
rect 9737 13917 9803 13933
rect 9845 13967 9911 13983
rect 10865 13971 10895 14119
rect 10965 13971 10995 14119
rect 11069 13971 11099 14119
rect 11155 13971 11185 14119
rect 13045 14187 13075 14213
rect 12845 14163 12911 14173
rect 12845 14129 12861 14163
rect 12895 14129 12911 14163
rect 12845 14119 12911 14129
rect 12683 14071 12713 14097
rect 12779 14071 12809 14097
rect 12851 14071 12881 14119
rect 12947 14071 12977 14097
rect 11321 13971 11351 14003
rect 9845 13933 9861 13967
rect 9895 13933 9911 13967
rect 9845 13917 9911 13933
rect 10807 13955 10895 13971
rect 10807 13921 10817 13955
rect 10851 13921 10895 13955
rect 9737 13877 9767 13917
rect 9845 13895 9875 13917
rect 10807 13905 10895 13921
rect 9653 13767 9683 13793
rect 9737 13767 9767 13793
rect 10865 13837 10895 13905
rect 10953 13955 11007 13971
rect 10953 13921 10963 13955
rect 10997 13921 11007 13955
rect 10953 13905 11007 13921
rect 11059 13955 11113 13971
rect 11059 13921 11069 13955
rect 11103 13921 11113 13955
rect 11059 13905 11113 13921
rect 11155 13955 11219 13971
rect 11155 13921 11165 13955
rect 11199 13921 11219 13955
rect 11155 13905 11219 13921
rect 11266 13955 11351 13971
rect 12683 13955 12713 13987
rect 12779 13955 12809 13987
rect 11266 13921 11276 13955
rect 11310 13921 11351 13955
rect 11266 13905 11351 13921
rect 10953 13837 10983 13905
rect 11059 13837 11089 13905
rect 11155 13837 11185 13905
rect 11321 13883 11351 13905
rect 12629 13939 12713 13955
rect 12629 13905 12639 13939
rect 12673 13905 12713 13939
rect 12629 13889 12713 13905
rect 12755 13939 12809 13955
rect 12755 13905 12765 13939
rect 12799 13905 12809 13939
rect 12755 13889 12809 13905
rect 9845 13739 9875 13765
rect 12045 13829 12075 13855
rect 10865 13727 10895 13753
rect 10953 13727 10983 13753
rect 11059 13727 11089 13753
rect 11155 13727 11185 13753
rect 11321 13727 11351 13753
rect 11876 13713 11906 13739
rect 11948 13713 11978 13739
rect 12683 13827 12713 13889
rect 12779 13827 12809 13889
rect 12851 13872 12881 13987
rect 12947 13955 12977 13987
rect 13045 13955 13075 13987
rect 12931 13939 12985 13955
rect 12931 13905 12941 13939
rect 12975 13905 12985 13939
rect 12931 13889 12985 13905
rect 13027 13939 13082 13955
rect 13027 13905 13037 13939
rect 13071 13905 13082 13939
rect 13027 13889 13082 13905
rect 12851 13871 12892 13872
rect 12851 13842 12893 13871
rect 12863 13827 12893 13842
rect 12947 13827 12977 13889
rect 13045 13867 13075 13889
rect 12683 13717 12713 13743
rect 12779 13717 12809 13743
rect 12863 13717 12893 13743
rect 12947 13717 12977 13743
rect 13045 13711 13075 13737
rect 11876 13597 11906 13629
rect 11806 13581 11906 13597
rect 11806 13547 11822 13581
rect 11856 13547 11906 13581
rect 11806 13531 11906 13547
rect 11948 13597 11978 13629
rect 12045 13597 12075 13629
rect 11948 13581 12002 13597
rect 11948 13547 11958 13581
rect 11992 13547 12002 13581
rect 11948 13531 12002 13547
rect 12045 13581 12111 13597
rect 12045 13547 12061 13581
rect 12095 13547 12111 13581
rect 12045 13531 12111 13547
rect 11864 13463 11894 13531
rect 11948 13463 11978 13531
rect 12045 13509 12075 13531
rect 11261 13361 11291 13387
rect 11073 13340 11127 13356
rect 9519 13291 9549 13317
rect 9603 13291 9633 13317
rect 9687 13291 9717 13317
rect 9771 13291 9801 13317
rect 9959 13291 9989 13317
rect 11073 13306 11083 13340
rect 11117 13306 11127 13340
rect 11073 13290 11127 13306
rect 10989 13248 11019 13289
rect 11073 13248 11103 13290
rect 11166 13248 11196 13274
rect 10989 13115 11019 13164
rect 11073 13146 11103 13164
rect 9519 13059 9549 13091
rect 9603 13059 9633 13091
rect 9687 13059 9717 13091
rect 9771 13059 9801 13091
rect 9959 13059 9989 13091
rect 9507 13043 9561 13059
rect 9507 13009 9517 13043
rect 9551 13009 9561 13043
rect 9507 12993 9561 13009
rect 9603 13043 9717 13059
rect 9603 13009 9634 13043
rect 9668 13009 9717 13043
rect 9603 12993 9717 13009
rect 9759 13043 9813 13059
rect 9759 13009 9769 13043
rect 9803 13009 9813 13043
rect 9759 12993 9813 13009
rect 9855 13043 9989 13059
rect 9855 13009 9865 13043
rect 9899 13026 9989 13043
rect 10935 13067 11019 13115
rect 10935 13033 10945 13067
rect 10979 13033 11019 13067
rect 9899 13009 9985 13026
rect 10935 13010 11019 13033
rect 9855 12993 9985 13009
rect 10989 12995 11019 13010
rect 11061 13121 11103 13146
rect 11166 13123 11196 13164
rect 11864 13353 11894 13379
rect 11948 13353 11978 13379
rect 12045 13353 12075 13379
rect 11261 13129 11291 13161
rect 11061 12995 11091 13121
rect 11145 13107 11199 13123
rect 11145 13090 11155 13107
rect 11133 13073 11155 13090
rect 11189 13073 11199 13107
rect 11133 13057 11199 13073
rect 11241 13113 11295 13129
rect 11241 13079 11251 13113
rect 11285 13079 11295 13113
rect 11241 13063 11295 13079
rect 11133 13034 11175 13057
rect 11261 13041 11291 13063
rect 11133 13010 11170 13034
rect 11133 12995 11163 13010
rect 9519 12971 9549 12993
rect 9603 12971 9633 12993
rect 9687 12971 9717 12993
rect 9771 12971 9801 12993
rect 9955 12971 9985 12993
rect 10989 12885 11019 12911
rect 11061 12885 11091 12911
rect 11133 12885 11163 12911
rect 11261 12885 11291 12911
rect 9519 12815 9549 12841
rect 9603 12815 9633 12841
rect 9687 12815 9717 12841
rect 9771 12815 9801 12841
rect 9955 12815 9985 12841
rect 9837 12547 9867 12573
rect 9645 12505 9675 12531
rect 9729 12505 9759 12531
rect 9645 12315 9675 12421
rect 9588 12299 9675 12315
rect 9588 12265 9604 12299
rect 9638 12265 9675 12299
rect 9588 12249 9675 12265
rect 9645 12209 9675 12249
rect 9729 12315 9759 12421
rect 9837 12315 9867 12347
rect 11213 12341 11243 12367
rect 9729 12299 9795 12315
rect 9729 12265 9745 12299
rect 9779 12265 9795 12299
rect 9729 12249 9795 12265
rect 9837 12299 9903 12315
rect 11021 12299 11051 12325
rect 11105 12299 11135 12325
rect 9837 12265 9853 12299
rect 9887 12265 9903 12299
rect 9837 12249 9903 12265
rect 9729 12209 9759 12249
rect 9837 12227 9867 12249
rect 9645 12099 9675 12125
rect 9729 12099 9759 12125
rect 11021 12109 11051 12215
rect 9837 12071 9867 12097
rect 10964 12093 11051 12109
rect 10964 12059 10980 12093
rect 11014 12059 11051 12093
rect 10964 12043 11051 12059
rect 11021 12003 11051 12043
rect 11105 12109 11135 12215
rect 11213 12109 11243 12141
rect 11105 12093 11171 12109
rect 11105 12059 11121 12093
rect 11155 12059 11171 12093
rect 11105 12043 11171 12059
rect 11213 12093 11279 12109
rect 11213 12059 11229 12093
rect 11263 12059 11279 12093
rect 11213 12043 11279 12059
rect 11105 12003 11135 12043
rect 11213 12021 11243 12043
rect 11021 11893 11051 11919
rect 11105 11893 11135 11919
rect 11213 11865 11243 11891
rect 9529 11727 9559 11753
rect 9613 11727 9643 11753
rect 9697 11727 9727 11753
rect 9781 11727 9811 11753
rect 9969 11727 9999 11753
rect 9529 11495 9559 11527
rect 9613 11495 9643 11527
rect 9697 11495 9727 11527
rect 9781 11495 9811 11527
rect 9969 11495 9999 11527
rect 9517 11479 9571 11495
rect 9517 11445 9527 11479
rect 9561 11445 9571 11479
rect 9517 11429 9571 11445
rect 9613 11479 9727 11495
rect 9613 11445 9644 11479
rect 9678 11445 9727 11479
rect 9613 11429 9727 11445
rect 9769 11479 9823 11495
rect 9769 11445 9779 11479
rect 9813 11445 9823 11479
rect 9769 11429 9823 11445
rect 9865 11479 9999 11495
rect 9865 11445 9875 11479
rect 9909 11462 9999 11479
rect 9909 11445 9995 11462
rect 9865 11429 9995 11445
rect 9529 11407 9559 11429
rect 9613 11407 9643 11429
rect 9697 11407 9727 11429
rect 9781 11407 9811 11429
rect 9965 11407 9995 11429
rect 9529 11251 9559 11277
rect 9613 11251 9643 11277
rect 9697 11251 9727 11277
rect 9781 11251 9811 11277
rect 9965 11251 9995 11277
rect 9847 10983 9877 11009
rect 9655 10941 9685 10967
rect 9739 10941 9769 10967
rect 9655 10751 9685 10857
rect 9598 10735 9685 10751
rect 9598 10701 9614 10735
rect 9648 10701 9685 10735
rect 9598 10685 9685 10701
rect 9655 10645 9685 10685
rect 9739 10751 9769 10857
rect 9847 10751 9877 10783
rect 9739 10735 9805 10751
rect 9739 10701 9755 10735
rect 9789 10701 9805 10735
rect 9739 10685 9805 10701
rect 9847 10735 9913 10751
rect 9847 10701 9863 10735
rect 9897 10701 9913 10735
rect 9847 10685 9913 10701
rect 9739 10645 9769 10685
rect 9847 10663 9877 10685
rect 9655 10535 9685 10561
rect 9739 10535 9769 10561
rect 9847 10507 9877 10533
rect 6238 6553 6268 6579
rect 6238 6401 6268 6423
rect 6238 6385 6324 6401
rect 6238 6351 6274 6385
rect 6308 6351 6324 6385
rect 6238 6335 6324 6351
rect 6238 6303 6268 6335
rect 6238 6077 6268 6103
rect 9332 5921 9362 5947
rect 9431 5921 9461 5947
rect 9527 5921 9557 5947
rect 9599 5921 9629 5947
rect 9695 5921 9725 5947
rect 9784 5921 9814 5947
rect 9868 5921 9898 5947
rect 9952 5921 9982 5947
rect 10140 5921 10170 5947
rect 10224 5921 10254 5947
rect 10308 5921 10338 5947
rect 10392 5921 10422 5947
rect 10482 5921 10512 5947
rect 10581 5921 10611 5947
rect 9332 5769 9362 5791
rect 9431 5777 9461 5837
rect 9332 5753 9386 5769
rect 9332 5719 9342 5753
rect 9376 5719 9386 5753
rect 9332 5703 9386 5719
rect 9431 5761 9485 5777
rect 9431 5727 9441 5761
rect 9475 5727 9485 5761
rect 9431 5711 9485 5727
rect 9332 5671 9362 5703
rect 1950 5501 1980 5527
rect 2049 5501 2079 5527
rect 2145 5501 2175 5527
rect 2217 5501 2247 5527
rect 2313 5501 2343 5527
rect 2402 5501 2432 5527
rect 2486 5501 2516 5527
rect 2570 5501 2600 5527
rect 2758 5501 2788 5527
rect 2842 5501 2872 5527
rect 2926 5501 2956 5527
rect 3010 5501 3040 5527
rect 3100 5501 3130 5527
rect 3199 5501 3229 5527
rect 1950 5349 1980 5371
rect 2049 5357 2079 5417
rect 1950 5333 2004 5349
rect 1950 5299 1960 5333
rect 1994 5299 2004 5333
rect 1950 5283 2004 5299
rect 2049 5341 2103 5357
rect 2049 5307 2059 5341
rect 2093 5307 2103 5341
rect 2049 5291 2103 5307
rect 1950 5251 1980 5283
rect 2049 5135 2079 5291
rect 2145 5245 2175 5417
rect 2121 5229 2175 5245
rect 2121 5195 2131 5229
rect 2165 5195 2175 5229
rect 2121 5179 2175 5195
rect 2145 5135 2175 5179
rect 2217 5245 2247 5417
rect 2313 5373 2343 5417
rect 2402 5373 2432 5417
rect 2486 5402 2516 5417
rect 2289 5357 2343 5373
rect 2289 5323 2299 5357
rect 2333 5323 2343 5357
rect 2289 5307 2343 5323
rect 2389 5357 2443 5373
rect 2389 5323 2399 5357
rect 2433 5323 2443 5357
rect 2389 5307 2443 5323
rect 2485 5372 2516 5402
rect 2570 5402 2600 5417
rect 2758 5402 2788 5417
rect 2570 5372 2788 5402
rect 2217 5229 2271 5245
rect 2217 5195 2227 5229
rect 2261 5195 2271 5229
rect 2217 5179 2271 5195
rect 2217 5135 2247 5179
rect 2313 5135 2343 5307
rect 2402 5135 2432 5307
rect 2485 5261 2515 5372
rect 2570 5357 2611 5372
rect 2581 5261 2611 5357
rect 2842 5342 2872 5417
rect 2926 5343 2956 5417
rect 2818 5326 2872 5342
rect 2818 5292 2828 5326
rect 2862 5292 2872 5326
rect 2818 5276 2872 5292
rect 2914 5327 2968 5343
rect 2914 5293 2924 5327
rect 2958 5293 2968 5327
rect 2914 5277 2968 5293
rect 2474 5245 2528 5261
rect 2474 5211 2484 5245
rect 2518 5211 2528 5245
rect 2474 5195 2528 5211
rect 2581 5245 2645 5261
rect 2581 5211 2601 5245
rect 2635 5211 2645 5245
rect 2486 5135 2516 5195
rect 2581 5180 2645 5211
rect 2570 5150 2788 5180
rect 2570 5135 2600 5150
rect 2758 5135 2788 5150
rect 2842 5135 2872 5276
rect 2926 5135 2956 5277
rect 3010 5238 3040 5417
rect 3100 5349 3130 5417
rect 3820 5497 3850 5523
rect 3919 5497 3949 5523
rect 4015 5497 4045 5523
rect 4087 5497 4117 5523
rect 4183 5497 4213 5523
rect 4272 5497 4302 5523
rect 4356 5497 4386 5523
rect 4440 5497 4470 5523
rect 4628 5497 4658 5523
rect 4712 5497 4742 5523
rect 4796 5497 4826 5523
rect 4880 5497 4910 5523
rect 4970 5497 5000 5523
rect 5069 5497 5099 5523
rect 3199 5349 3229 5371
rect 3082 5333 3136 5349
rect 3082 5299 3092 5333
rect 3126 5299 3136 5333
rect 3082 5283 3136 5299
rect 3178 5333 3232 5349
rect 3178 5299 3188 5333
rect 3222 5299 3232 5333
rect 3178 5283 3232 5299
rect 3820 5345 3850 5367
rect 3919 5353 3949 5413
rect 3820 5329 3874 5345
rect 3820 5295 3830 5329
rect 3864 5295 3874 5329
rect 3004 5222 3058 5238
rect 3004 5188 3014 5222
rect 3048 5188 3058 5222
rect 3004 5172 3058 5188
rect 3010 5135 3040 5172
rect 3100 5135 3130 5283
rect 3199 5251 3229 5283
rect 3820 5279 3874 5295
rect 3919 5337 3973 5353
rect 3919 5303 3929 5337
rect 3963 5303 3973 5337
rect 3919 5287 3973 5303
rect 3820 5247 3850 5279
rect 1950 5025 1980 5051
rect 2049 5025 2079 5051
rect 2145 5025 2175 5051
rect 2217 5025 2247 5051
rect 2313 5025 2343 5051
rect 2402 5025 2432 5051
rect 2486 5025 2516 5051
rect 2570 5025 2600 5051
rect 2758 5025 2788 5051
rect 2842 5025 2872 5051
rect 2926 5025 2956 5051
rect 3010 5025 3040 5051
rect 3100 5025 3130 5051
rect 3199 5025 3229 5051
rect 3919 5131 3949 5287
rect 4015 5241 4045 5413
rect 3991 5225 4045 5241
rect 3991 5191 4001 5225
rect 4035 5191 4045 5225
rect 3991 5175 4045 5191
rect 4015 5131 4045 5175
rect 4087 5241 4117 5413
rect 4183 5369 4213 5413
rect 4272 5369 4302 5413
rect 4356 5398 4386 5413
rect 4159 5353 4213 5369
rect 4159 5319 4169 5353
rect 4203 5319 4213 5353
rect 4159 5303 4213 5319
rect 4259 5353 4313 5369
rect 4259 5319 4269 5353
rect 4303 5319 4313 5353
rect 4259 5303 4313 5319
rect 4355 5368 4386 5398
rect 4440 5398 4470 5413
rect 4628 5398 4658 5413
rect 4440 5368 4658 5398
rect 4087 5225 4141 5241
rect 4087 5191 4097 5225
rect 4131 5191 4141 5225
rect 4087 5175 4141 5191
rect 4087 5131 4117 5175
rect 4183 5131 4213 5303
rect 4272 5131 4302 5303
rect 4355 5257 4385 5368
rect 4440 5353 4481 5368
rect 4451 5257 4481 5353
rect 4712 5338 4742 5413
rect 4796 5339 4826 5413
rect 4688 5322 4742 5338
rect 4688 5288 4698 5322
rect 4732 5288 4742 5322
rect 4688 5272 4742 5288
rect 4784 5323 4838 5339
rect 4784 5289 4794 5323
rect 4828 5289 4838 5323
rect 4784 5273 4838 5289
rect 4344 5241 4398 5257
rect 4344 5207 4354 5241
rect 4388 5207 4398 5241
rect 4344 5191 4398 5207
rect 4451 5241 4515 5257
rect 4451 5207 4471 5241
rect 4505 5207 4515 5241
rect 4356 5131 4386 5191
rect 4451 5176 4515 5207
rect 4440 5146 4658 5176
rect 4440 5131 4470 5146
rect 4628 5131 4658 5146
rect 4712 5131 4742 5272
rect 4796 5131 4826 5273
rect 4880 5234 4910 5413
rect 4970 5345 5000 5413
rect 5636 5493 5666 5519
rect 5735 5493 5765 5519
rect 5831 5493 5861 5519
rect 5903 5493 5933 5519
rect 5999 5493 6029 5519
rect 6088 5493 6118 5519
rect 6172 5493 6202 5519
rect 6256 5493 6286 5519
rect 6444 5493 6474 5519
rect 6528 5493 6558 5519
rect 6612 5493 6642 5519
rect 6696 5493 6726 5519
rect 6786 5493 6816 5519
rect 6885 5493 6915 5519
rect 5069 5345 5099 5367
rect 4952 5329 5006 5345
rect 4952 5295 4962 5329
rect 4996 5295 5006 5329
rect 4952 5279 5006 5295
rect 5048 5329 5102 5345
rect 5048 5295 5058 5329
rect 5092 5295 5102 5329
rect 5048 5279 5102 5295
rect 5636 5341 5666 5363
rect 5735 5349 5765 5409
rect 5636 5325 5690 5341
rect 5636 5291 5646 5325
rect 5680 5291 5690 5325
rect 4874 5218 4928 5234
rect 4874 5184 4884 5218
rect 4918 5184 4928 5218
rect 4874 5168 4928 5184
rect 4880 5131 4910 5168
rect 4970 5131 5000 5279
rect 5069 5247 5099 5279
rect 5636 5275 5690 5291
rect 5735 5333 5789 5349
rect 5735 5299 5745 5333
rect 5779 5299 5789 5333
rect 5735 5283 5789 5299
rect 5636 5243 5666 5275
rect 3820 5021 3850 5047
rect 3919 5021 3949 5047
rect 4015 5021 4045 5047
rect 4087 5021 4117 5047
rect 4183 5021 4213 5047
rect 4272 5021 4302 5047
rect 4356 5021 4386 5047
rect 4440 5021 4470 5047
rect 4628 5021 4658 5047
rect 4712 5021 4742 5047
rect 4796 5021 4826 5047
rect 4880 5021 4910 5047
rect 4970 5021 5000 5047
rect 5069 5021 5099 5047
rect 5735 5127 5765 5283
rect 5831 5237 5861 5409
rect 5807 5221 5861 5237
rect 5807 5187 5817 5221
rect 5851 5187 5861 5221
rect 5807 5171 5861 5187
rect 5831 5127 5861 5171
rect 5903 5237 5933 5409
rect 5999 5365 6029 5409
rect 6088 5365 6118 5409
rect 6172 5394 6202 5409
rect 5975 5349 6029 5365
rect 5975 5315 5985 5349
rect 6019 5315 6029 5349
rect 5975 5299 6029 5315
rect 6075 5349 6129 5365
rect 6075 5315 6085 5349
rect 6119 5315 6129 5349
rect 6075 5299 6129 5315
rect 6171 5364 6202 5394
rect 6256 5394 6286 5409
rect 6444 5394 6474 5409
rect 6256 5364 6474 5394
rect 5903 5221 5957 5237
rect 5903 5187 5913 5221
rect 5947 5187 5957 5221
rect 5903 5171 5957 5187
rect 5903 5127 5933 5171
rect 5999 5127 6029 5299
rect 6088 5127 6118 5299
rect 6171 5253 6201 5364
rect 6256 5349 6297 5364
rect 6267 5253 6297 5349
rect 6528 5334 6558 5409
rect 6612 5335 6642 5409
rect 6504 5318 6558 5334
rect 6504 5284 6514 5318
rect 6548 5284 6558 5318
rect 6504 5268 6558 5284
rect 6600 5319 6654 5335
rect 6600 5285 6610 5319
rect 6644 5285 6654 5319
rect 6600 5269 6654 5285
rect 6160 5237 6214 5253
rect 6160 5203 6170 5237
rect 6204 5203 6214 5237
rect 6160 5187 6214 5203
rect 6267 5237 6331 5253
rect 6267 5203 6287 5237
rect 6321 5203 6331 5237
rect 6172 5127 6202 5187
rect 6267 5172 6331 5203
rect 6256 5142 6474 5172
rect 6256 5127 6286 5142
rect 6444 5127 6474 5142
rect 6528 5127 6558 5268
rect 6612 5127 6642 5269
rect 6696 5230 6726 5409
rect 6786 5341 6816 5409
rect 7506 5489 7536 5515
rect 7605 5489 7635 5515
rect 7701 5489 7731 5515
rect 7773 5489 7803 5515
rect 7869 5489 7899 5515
rect 7958 5489 7988 5515
rect 8042 5489 8072 5515
rect 8126 5489 8156 5515
rect 8314 5489 8344 5515
rect 8398 5489 8428 5515
rect 8482 5489 8512 5515
rect 8566 5489 8596 5515
rect 8656 5489 8686 5515
rect 8755 5489 8785 5515
rect 6885 5341 6915 5363
rect 6768 5325 6822 5341
rect 6768 5291 6778 5325
rect 6812 5291 6822 5325
rect 6768 5275 6822 5291
rect 6864 5325 6918 5341
rect 6864 5291 6874 5325
rect 6908 5291 6918 5325
rect 6864 5275 6918 5291
rect 7506 5337 7536 5359
rect 7605 5345 7635 5405
rect 7506 5321 7560 5337
rect 7506 5287 7516 5321
rect 7550 5287 7560 5321
rect 6690 5214 6744 5230
rect 6690 5180 6700 5214
rect 6734 5180 6744 5214
rect 6690 5164 6744 5180
rect 6696 5127 6726 5164
rect 6786 5127 6816 5275
rect 6885 5243 6915 5275
rect 7506 5271 7560 5287
rect 7605 5329 7659 5345
rect 7605 5295 7615 5329
rect 7649 5295 7659 5329
rect 7605 5279 7659 5295
rect 7506 5239 7536 5271
rect 5636 5017 5666 5043
rect 5735 5017 5765 5043
rect 5831 5017 5861 5043
rect 5903 5017 5933 5043
rect 5999 5017 6029 5043
rect 6088 5017 6118 5043
rect 6172 5017 6202 5043
rect 6256 5017 6286 5043
rect 6444 5017 6474 5043
rect 6528 5017 6558 5043
rect 6612 5017 6642 5043
rect 6696 5017 6726 5043
rect 6786 5017 6816 5043
rect 6885 5017 6915 5043
rect 7605 5123 7635 5279
rect 7701 5233 7731 5405
rect 7677 5217 7731 5233
rect 7677 5183 7687 5217
rect 7721 5183 7731 5217
rect 7677 5167 7731 5183
rect 7701 5123 7731 5167
rect 7773 5233 7803 5405
rect 7869 5361 7899 5405
rect 7958 5361 7988 5405
rect 8042 5390 8072 5405
rect 7845 5345 7899 5361
rect 7845 5311 7855 5345
rect 7889 5311 7899 5345
rect 7845 5295 7899 5311
rect 7945 5345 7999 5361
rect 7945 5311 7955 5345
rect 7989 5311 7999 5345
rect 7945 5295 7999 5311
rect 8041 5360 8072 5390
rect 8126 5390 8156 5405
rect 8314 5390 8344 5405
rect 8126 5360 8344 5390
rect 7773 5217 7827 5233
rect 7773 5183 7783 5217
rect 7817 5183 7827 5217
rect 7773 5167 7827 5183
rect 7773 5123 7803 5167
rect 7869 5123 7899 5295
rect 7958 5123 7988 5295
rect 8041 5249 8071 5360
rect 8126 5345 8167 5360
rect 8137 5249 8167 5345
rect 8398 5330 8428 5405
rect 8482 5331 8512 5405
rect 8374 5314 8428 5330
rect 8374 5280 8384 5314
rect 8418 5280 8428 5314
rect 8374 5264 8428 5280
rect 8470 5315 8524 5331
rect 8470 5281 8480 5315
rect 8514 5281 8524 5315
rect 8470 5265 8524 5281
rect 8030 5233 8084 5249
rect 8030 5199 8040 5233
rect 8074 5199 8084 5233
rect 8030 5183 8084 5199
rect 8137 5233 8201 5249
rect 8137 5199 8157 5233
rect 8191 5199 8201 5233
rect 8042 5123 8072 5183
rect 8137 5168 8201 5199
rect 8126 5138 8344 5168
rect 8126 5123 8156 5138
rect 8314 5123 8344 5138
rect 8398 5123 8428 5264
rect 8482 5123 8512 5265
rect 8566 5226 8596 5405
rect 8656 5337 8686 5405
rect 9431 5555 9461 5711
rect 9527 5665 9557 5837
rect 9503 5649 9557 5665
rect 9503 5615 9513 5649
rect 9547 5615 9557 5649
rect 9503 5599 9557 5615
rect 9527 5555 9557 5599
rect 9599 5665 9629 5837
rect 9695 5793 9725 5837
rect 9784 5793 9814 5837
rect 9868 5822 9898 5837
rect 9671 5777 9725 5793
rect 9671 5743 9681 5777
rect 9715 5743 9725 5777
rect 9671 5727 9725 5743
rect 9771 5777 9825 5793
rect 9771 5743 9781 5777
rect 9815 5743 9825 5777
rect 9771 5727 9825 5743
rect 9867 5792 9898 5822
rect 9952 5822 9982 5837
rect 10140 5822 10170 5837
rect 9952 5792 10170 5822
rect 9599 5649 9653 5665
rect 9599 5615 9609 5649
rect 9643 5615 9653 5649
rect 9599 5599 9653 5615
rect 9599 5555 9629 5599
rect 9695 5555 9725 5727
rect 9784 5555 9814 5727
rect 9867 5681 9897 5792
rect 9952 5777 9993 5792
rect 9963 5681 9993 5777
rect 10224 5762 10254 5837
rect 10308 5763 10338 5837
rect 10200 5746 10254 5762
rect 10200 5712 10210 5746
rect 10244 5712 10254 5746
rect 10200 5696 10254 5712
rect 10296 5747 10350 5763
rect 10296 5713 10306 5747
rect 10340 5713 10350 5747
rect 10296 5697 10350 5713
rect 9856 5665 9910 5681
rect 9856 5631 9866 5665
rect 9900 5631 9910 5665
rect 9856 5615 9910 5631
rect 9963 5665 10027 5681
rect 9963 5631 9983 5665
rect 10017 5631 10027 5665
rect 9868 5555 9898 5615
rect 9963 5600 10027 5631
rect 9952 5570 10170 5600
rect 9952 5555 9982 5570
rect 10140 5555 10170 5570
rect 10224 5555 10254 5696
rect 10308 5555 10338 5697
rect 10392 5658 10422 5837
rect 10482 5769 10512 5837
rect 11202 5917 11232 5943
rect 11301 5917 11331 5943
rect 11397 5917 11427 5943
rect 11469 5917 11499 5943
rect 11565 5917 11595 5943
rect 11654 5917 11684 5943
rect 11738 5917 11768 5943
rect 11822 5917 11852 5943
rect 12010 5917 12040 5943
rect 12094 5917 12124 5943
rect 12178 5917 12208 5943
rect 12262 5917 12292 5943
rect 12352 5917 12382 5943
rect 12451 5917 12481 5943
rect 10581 5769 10611 5791
rect 10464 5753 10518 5769
rect 10464 5719 10474 5753
rect 10508 5719 10518 5753
rect 10464 5703 10518 5719
rect 10560 5753 10614 5769
rect 10560 5719 10570 5753
rect 10604 5719 10614 5753
rect 10560 5703 10614 5719
rect 11202 5765 11232 5787
rect 11301 5773 11331 5833
rect 11202 5749 11256 5765
rect 11202 5715 11212 5749
rect 11246 5715 11256 5749
rect 10386 5642 10440 5658
rect 10386 5608 10396 5642
rect 10430 5608 10440 5642
rect 10386 5592 10440 5608
rect 10392 5555 10422 5592
rect 10482 5555 10512 5703
rect 10581 5671 10611 5703
rect 11202 5699 11256 5715
rect 11301 5757 11355 5773
rect 11301 5723 11311 5757
rect 11345 5723 11355 5757
rect 11301 5707 11355 5723
rect 11202 5667 11232 5699
rect 9332 5445 9362 5471
rect 9431 5445 9461 5471
rect 9527 5445 9557 5471
rect 9599 5445 9629 5471
rect 9695 5445 9725 5471
rect 9784 5445 9814 5471
rect 9868 5445 9898 5471
rect 9952 5445 9982 5471
rect 10140 5445 10170 5471
rect 10224 5445 10254 5471
rect 10308 5445 10338 5471
rect 10392 5445 10422 5471
rect 10482 5445 10512 5471
rect 10581 5445 10611 5471
rect 11301 5551 11331 5707
rect 11397 5661 11427 5833
rect 11373 5645 11427 5661
rect 11373 5611 11383 5645
rect 11417 5611 11427 5645
rect 11373 5595 11427 5611
rect 11397 5551 11427 5595
rect 11469 5661 11499 5833
rect 11565 5789 11595 5833
rect 11654 5789 11684 5833
rect 11738 5818 11768 5833
rect 11541 5773 11595 5789
rect 11541 5739 11551 5773
rect 11585 5739 11595 5773
rect 11541 5723 11595 5739
rect 11641 5773 11695 5789
rect 11641 5739 11651 5773
rect 11685 5739 11695 5773
rect 11641 5723 11695 5739
rect 11737 5788 11768 5818
rect 11822 5818 11852 5833
rect 12010 5818 12040 5833
rect 11822 5788 12040 5818
rect 11469 5645 11523 5661
rect 11469 5611 11479 5645
rect 11513 5611 11523 5645
rect 11469 5595 11523 5611
rect 11469 5551 11499 5595
rect 11565 5551 11595 5723
rect 11654 5551 11684 5723
rect 11737 5677 11767 5788
rect 11822 5773 11863 5788
rect 11833 5677 11863 5773
rect 12094 5758 12124 5833
rect 12178 5759 12208 5833
rect 12070 5742 12124 5758
rect 12070 5708 12080 5742
rect 12114 5708 12124 5742
rect 12070 5692 12124 5708
rect 12166 5743 12220 5759
rect 12166 5709 12176 5743
rect 12210 5709 12220 5743
rect 12166 5693 12220 5709
rect 11726 5661 11780 5677
rect 11726 5627 11736 5661
rect 11770 5627 11780 5661
rect 11726 5611 11780 5627
rect 11833 5661 11897 5677
rect 11833 5627 11853 5661
rect 11887 5627 11897 5661
rect 11738 5551 11768 5611
rect 11833 5596 11897 5627
rect 11822 5566 12040 5596
rect 11822 5551 11852 5566
rect 12010 5551 12040 5566
rect 12094 5551 12124 5692
rect 12178 5551 12208 5693
rect 12262 5654 12292 5833
rect 12352 5765 12382 5833
rect 13018 5913 13048 5939
rect 13117 5913 13147 5939
rect 13213 5913 13243 5939
rect 13285 5913 13315 5939
rect 13381 5913 13411 5939
rect 13470 5913 13500 5939
rect 13554 5913 13584 5939
rect 13638 5913 13668 5939
rect 13826 5913 13856 5939
rect 13910 5913 13940 5939
rect 13994 5913 14024 5939
rect 14078 5913 14108 5939
rect 14168 5913 14198 5939
rect 14267 5913 14297 5939
rect 12451 5765 12481 5787
rect 12334 5749 12388 5765
rect 12334 5715 12344 5749
rect 12378 5715 12388 5749
rect 12334 5699 12388 5715
rect 12430 5749 12484 5765
rect 12430 5715 12440 5749
rect 12474 5715 12484 5749
rect 12430 5699 12484 5715
rect 13018 5761 13048 5783
rect 13117 5769 13147 5829
rect 13018 5745 13072 5761
rect 13018 5711 13028 5745
rect 13062 5711 13072 5745
rect 12256 5638 12310 5654
rect 12256 5604 12266 5638
rect 12300 5604 12310 5638
rect 12256 5588 12310 5604
rect 12262 5551 12292 5588
rect 12352 5551 12382 5699
rect 12451 5667 12481 5699
rect 13018 5695 13072 5711
rect 13117 5753 13171 5769
rect 13117 5719 13127 5753
rect 13161 5719 13171 5753
rect 13117 5703 13171 5719
rect 13018 5663 13048 5695
rect 11202 5441 11232 5467
rect 11301 5441 11331 5467
rect 11397 5441 11427 5467
rect 11469 5441 11499 5467
rect 11565 5441 11595 5467
rect 11654 5441 11684 5467
rect 11738 5441 11768 5467
rect 11822 5441 11852 5467
rect 12010 5441 12040 5467
rect 12094 5441 12124 5467
rect 12178 5441 12208 5467
rect 12262 5441 12292 5467
rect 12352 5441 12382 5467
rect 12451 5441 12481 5467
rect 13117 5547 13147 5703
rect 13213 5657 13243 5829
rect 13189 5641 13243 5657
rect 13189 5607 13199 5641
rect 13233 5607 13243 5641
rect 13189 5591 13243 5607
rect 13213 5547 13243 5591
rect 13285 5657 13315 5829
rect 13381 5785 13411 5829
rect 13470 5785 13500 5829
rect 13554 5814 13584 5829
rect 13357 5769 13411 5785
rect 13357 5735 13367 5769
rect 13401 5735 13411 5769
rect 13357 5719 13411 5735
rect 13457 5769 13511 5785
rect 13457 5735 13467 5769
rect 13501 5735 13511 5769
rect 13457 5719 13511 5735
rect 13553 5784 13584 5814
rect 13638 5814 13668 5829
rect 13826 5814 13856 5829
rect 13638 5784 13856 5814
rect 13285 5641 13339 5657
rect 13285 5607 13295 5641
rect 13329 5607 13339 5641
rect 13285 5591 13339 5607
rect 13285 5547 13315 5591
rect 13381 5547 13411 5719
rect 13470 5547 13500 5719
rect 13553 5673 13583 5784
rect 13638 5769 13679 5784
rect 13649 5673 13679 5769
rect 13910 5754 13940 5829
rect 13994 5755 14024 5829
rect 13886 5738 13940 5754
rect 13886 5704 13896 5738
rect 13930 5704 13940 5738
rect 13886 5688 13940 5704
rect 13982 5739 14036 5755
rect 13982 5705 13992 5739
rect 14026 5705 14036 5739
rect 13982 5689 14036 5705
rect 13542 5657 13596 5673
rect 13542 5623 13552 5657
rect 13586 5623 13596 5657
rect 13542 5607 13596 5623
rect 13649 5657 13713 5673
rect 13649 5623 13669 5657
rect 13703 5623 13713 5657
rect 13554 5547 13584 5607
rect 13649 5592 13713 5623
rect 13638 5562 13856 5592
rect 13638 5547 13668 5562
rect 13826 5547 13856 5562
rect 13910 5547 13940 5688
rect 13994 5547 14024 5689
rect 14078 5650 14108 5829
rect 14168 5761 14198 5829
rect 14888 5909 14918 5935
rect 14987 5909 15017 5935
rect 15083 5909 15113 5935
rect 15155 5909 15185 5935
rect 15251 5909 15281 5935
rect 15340 5909 15370 5935
rect 15424 5909 15454 5935
rect 15508 5909 15538 5935
rect 15696 5909 15726 5935
rect 15780 5909 15810 5935
rect 15864 5909 15894 5935
rect 15948 5909 15978 5935
rect 16038 5909 16068 5935
rect 16137 5909 16167 5935
rect 14267 5761 14297 5783
rect 14150 5745 14204 5761
rect 14150 5711 14160 5745
rect 14194 5711 14204 5745
rect 14150 5695 14204 5711
rect 14246 5745 14300 5761
rect 14246 5711 14256 5745
rect 14290 5711 14300 5745
rect 14246 5695 14300 5711
rect 14888 5757 14918 5779
rect 14987 5765 15017 5825
rect 14888 5741 14942 5757
rect 14888 5707 14898 5741
rect 14932 5707 14942 5741
rect 14072 5634 14126 5650
rect 14072 5600 14082 5634
rect 14116 5600 14126 5634
rect 14072 5584 14126 5600
rect 14078 5547 14108 5584
rect 14168 5547 14198 5695
rect 14267 5663 14297 5695
rect 14888 5691 14942 5707
rect 14987 5749 15041 5765
rect 14987 5715 14997 5749
rect 15031 5715 15041 5749
rect 14987 5699 15041 5715
rect 14888 5659 14918 5691
rect 13018 5437 13048 5463
rect 13117 5437 13147 5463
rect 13213 5437 13243 5463
rect 13285 5437 13315 5463
rect 13381 5437 13411 5463
rect 13470 5437 13500 5463
rect 13554 5437 13584 5463
rect 13638 5437 13668 5463
rect 13826 5437 13856 5463
rect 13910 5437 13940 5463
rect 13994 5437 14024 5463
rect 14078 5437 14108 5463
rect 14168 5437 14198 5463
rect 14267 5437 14297 5463
rect 14987 5543 15017 5699
rect 15083 5653 15113 5825
rect 15059 5637 15113 5653
rect 15059 5603 15069 5637
rect 15103 5603 15113 5637
rect 15059 5587 15113 5603
rect 15083 5543 15113 5587
rect 15155 5653 15185 5825
rect 15251 5781 15281 5825
rect 15340 5781 15370 5825
rect 15424 5810 15454 5825
rect 15227 5765 15281 5781
rect 15227 5731 15237 5765
rect 15271 5731 15281 5765
rect 15227 5715 15281 5731
rect 15327 5765 15381 5781
rect 15327 5731 15337 5765
rect 15371 5731 15381 5765
rect 15327 5715 15381 5731
rect 15423 5780 15454 5810
rect 15508 5810 15538 5825
rect 15696 5810 15726 5825
rect 15508 5780 15726 5810
rect 15155 5637 15209 5653
rect 15155 5603 15165 5637
rect 15199 5603 15209 5637
rect 15155 5587 15209 5603
rect 15155 5543 15185 5587
rect 15251 5543 15281 5715
rect 15340 5543 15370 5715
rect 15423 5669 15453 5780
rect 15508 5765 15549 5780
rect 15519 5669 15549 5765
rect 15780 5750 15810 5825
rect 15864 5751 15894 5825
rect 15756 5734 15810 5750
rect 15756 5700 15766 5734
rect 15800 5700 15810 5734
rect 15756 5684 15810 5700
rect 15852 5735 15906 5751
rect 15852 5701 15862 5735
rect 15896 5701 15906 5735
rect 15852 5685 15906 5701
rect 15412 5653 15466 5669
rect 15412 5619 15422 5653
rect 15456 5619 15466 5653
rect 15412 5603 15466 5619
rect 15519 5653 15583 5669
rect 15519 5619 15539 5653
rect 15573 5619 15583 5653
rect 15424 5543 15454 5603
rect 15519 5588 15583 5619
rect 15508 5558 15726 5588
rect 15508 5543 15538 5558
rect 15696 5543 15726 5558
rect 15780 5543 15810 5684
rect 15864 5543 15894 5685
rect 15948 5646 15978 5825
rect 16038 5757 16068 5825
rect 16137 5757 16167 5779
rect 16020 5741 16074 5757
rect 16020 5707 16030 5741
rect 16064 5707 16074 5741
rect 16020 5691 16074 5707
rect 16116 5741 16170 5757
rect 16116 5707 16126 5741
rect 16160 5707 16170 5741
rect 16116 5691 16170 5707
rect 15942 5630 15996 5646
rect 15942 5596 15952 5630
rect 15986 5596 15996 5630
rect 15942 5580 15996 5596
rect 15948 5543 15978 5580
rect 16038 5543 16068 5691
rect 16137 5659 16167 5691
rect 14888 5433 14918 5459
rect 14987 5433 15017 5459
rect 15083 5433 15113 5459
rect 15155 5433 15185 5459
rect 15251 5433 15281 5459
rect 15340 5433 15370 5459
rect 15424 5433 15454 5459
rect 15508 5433 15538 5459
rect 15696 5433 15726 5459
rect 15780 5433 15810 5459
rect 15864 5433 15894 5459
rect 15948 5433 15978 5459
rect 16038 5433 16068 5459
rect 16137 5433 16167 5459
rect 8755 5337 8785 5359
rect 8638 5321 8692 5337
rect 8638 5287 8648 5321
rect 8682 5287 8692 5321
rect 8638 5271 8692 5287
rect 8734 5321 8788 5337
rect 8734 5287 8744 5321
rect 8778 5287 8788 5321
rect 8734 5271 8788 5287
rect 8560 5210 8614 5226
rect 8560 5176 8570 5210
rect 8604 5176 8614 5210
rect 8560 5160 8614 5176
rect 8566 5123 8596 5160
rect 8656 5123 8686 5271
rect 8755 5239 8785 5271
rect 9360 5047 9390 5073
rect 9459 5047 9489 5073
rect 9555 5047 9585 5073
rect 9627 5047 9657 5073
rect 9723 5047 9753 5073
rect 9812 5047 9842 5073
rect 9896 5047 9926 5073
rect 9980 5047 10010 5073
rect 10168 5047 10198 5073
rect 10252 5047 10282 5073
rect 10336 5047 10366 5073
rect 10420 5047 10450 5073
rect 10510 5047 10540 5073
rect 10609 5047 10639 5073
rect 7506 5013 7536 5039
rect 7605 5013 7635 5039
rect 7701 5013 7731 5039
rect 7773 5013 7803 5039
rect 7869 5013 7899 5039
rect 7958 5013 7988 5039
rect 8042 5013 8072 5039
rect 8126 5013 8156 5039
rect 8314 5013 8344 5039
rect 8398 5013 8428 5039
rect 8482 5013 8512 5039
rect 8566 5013 8596 5039
rect 8656 5013 8686 5039
rect 8755 5013 8785 5039
rect 9360 4895 9390 4917
rect 9459 4903 9489 4963
rect 9360 4879 9414 4895
rect 9360 4845 9370 4879
rect 9404 4845 9414 4879
rect 9360 4829 9414 4845
rect 9459 4887 9513 4903
rect 9459 4853 9469 4887
rect 9503 4853 9513 4887
rect 9459 4837 9513 4853
rect 9360 4797 9390 4829
rect 9459 4681 9489 4837
rect 9555 4791 9585 4963
rect 9531 4775 9585 4791
rect 9531 4741 9541 4775
rect 9575 4741 9585 4775
rect 9531 4725 9585 4741
rect 9555 4681 9585 4725
rect 9627 4791 9657 4963
rect 9723 4919 9753 4963
rect 9812 4919 9842 4963
rect 9896 4948 9926 4963
rect 9699 4903 9753 4919
rect 9699 4869 9709 4903
rect 9743 4869 9753 4903
rect 9699 4853 9753 4869
rect 9799 4903 9853 4919
rect 9799 4869 9809 4903
rect 9843 4869 9853 4903
rect 9799 4853 9853 4869
rect 9895 4918 9926 4948
rect 9980 4948 10010 4963
rect 10168 4948 10198 4963
rect 9980 4918 10198 4948
rect 9627 4775 9681 4791
rect 9627 4741 9637 4775
rect 9671 4741 9681 4775
rect 9627 4725 9681 4741
rect 9627 4681 9657 4725
rect 9723 4681 9753 4853
rect 9812 4681 9842 4853
rect 9895 4807 9925 4918
rect 9980 4903 10021 4918
rect 9991 4807 10021 4903
rect 10252 4888 10282 4963
rect 10336 4889 10366 4963
rect 10228 4872 10282 4888
rect 10228 4838 10238 4872
rect 10272 4838 10282 4872
rect 10228 4822 10282 4838
rect 10324 4873 10378 4889
rect 10324 4839 10334 4873
rect 10368 4839 10378 4873
rect 10324 4823 10378 4839
rect 9884 4791 9938 4807
rect 9884 4757 9894 4791
rect 9928 4757 9938 4791
rect 9884 4741 9938 4757
rect 9991 4791 10055 4807
rect 9991 4757 10011 4791
rect 10045 4757 10055 4791
rect 9896 4681 9926 4741
rect 9991 4726 10055 4757
rect 9980 4696 10198 4726
rect 9980 4681 10010 4696
rect 10168 4681 10198 4696
rect 10252 4681 10282 4822
rect 10336 4681 10366 4823
rect 10420 4784 10450 4963
rect 10510 4895 10540 4963
rect 11230 5043 11260 5069
rect 11329 5043 11359 5069
rect 11425 5043 11455 5069
rect 11497 5043 11527 5069
rect 11593 5043 11623 5069
rect 11682 5043 11712 5069
rect 11766 5043 11796 5069
rect 11850 5043 11880 5069
rect 12038 5043 12068 5069
rect 12122 5043 12152 5069
rect 12206 5043 12236 5069
rect 12290 5043 12320 5069
rect 12380 5043 12410 5069
rect 12479 5043 12509 5069
rect 10609 4895 10639 4917
rect 10492 4879 10546 4895
rect 10492 4845 10502 4879
rect 10536 4845 10546 4879
rect 10492 4829 10546 4845
rect 10588 4879 10642 4895
rect 10588 4845 10598 4879
rect 10632 4845 10642 4879
rect 10588 4829 10642 4845
rect 11230 4891 11260 4913
rect 11329 4899 11359 4959
rect 11230 4875 11284 4891
rect 11230 4841 11240 4875
rect 11274 4841 11284 4875
rect 10414 4768 10468 4784
rect 10414 4734 10424 4768
rect 10458 4734 10468 4768
rect 10414 4718 10468 4734
rect 10420 4681 10450 4718
rect 10510 4681 10540 4829
rect 10609 4797 10639 4829
rect 11230 4825 11284 4841
rect 11329 4883 11383 4899
rect 11329 4849 11339 4883
rect 11373 4849 11383 4883
rect 11329 4833 11383 4849
rect 11230 4793 11260 4825
rect 9360 4571 9390 4597
rect 9459 4571 9489 4597
rect 9555 4571 9585 4597
rect 9627 4571 9657 4597
rect 9723 4571 9753 4597
rect 9812 4571 9842 4597
rect 9896 4571 9926 4597
rect 9980 4571 10010 4597
rect 10168 4571 10198 4597
rect 10252 4571 10282 4597
rect 10336 4571 10366 4597
rect 10420 4571 10450 4597
rect 10510 4571 10540 4597
rect 10609 4571 10639 4597
rect 11329 4677 11359 4833
rect 11425 4787 11455 4959
rect 11401 4771 11455 4787
rect 11401 4737 11411 4771
rect 11445 4737 11455 4771
rect 11401 4721 11455 4737
rect 11425 4677 11455 4721
rect 11497 4787 11527 4959
rect 11593 4915 11623 4959
rect 11682 4915 11712 4959
rect 11766 4944 11796 4959
rect 11569 4899 11623 4915
rect 11569 4865 11579 4899
rect 11613 4865 11623 4899
rect 11569 4849 11623 4865
rect 11669 4899 11723 4915
rect 11669 4865 11679 4899
rect 11713 4865 11723 4899
rect 11669 4849 11723 4865
rect 11765 4914 11796 4944
rect 11850 4944 11880 4959
rect 12038 4944 12068 4959
rect 11850 4914 12068 4944
rect 11497 4771 11551 4787
rect 11497 4737 11507 4771
rect 11541 4737 11551 4771
rect 11497 4721 11551 4737
rect 11497 4677 11527 4721
rect 11593 4677 11623 4849
rect 11682 4677 11712 4849
rect 11765 4803 11795 4914
rect 11850 4899 11891 4914
rect 11861 4803 11891 4899
rect 12122 4884 12152 4959
rect 12206 4885 12236 4959
rect 12098 4868 12152 4884
rect 12098 4834 12108 4868
rect 12142 4834 12152 4868
rect 12098 4818 12152 4834
rect 12194 4869 12248 4885
rect 12194 4835 12204 4869
rect 12238 4835 12248 4869
rect 12194 4819 12248 4835
rect 11754 4787 11808 4803
rect 11754 4753 11764 4787
rect 11798 4753 11808 4787
rect 11754 4737 11808 4753
rect 11861 4787 11925 4803
rect 11861 4753 11881 4787
rect 11915 4753 11925 4787
rect 11766 4677 11796 4737
rect 11861 4722 11925 4753
rect 11850 4692 12068 4722
rect 11850 4677 11880 4692
rect 12038 4677 12068 4692
rect 12122 4677 12152 4818
rect 12206 4677 12236 4819
rect 12290 4780 12320 4959
rect 12380 4891 12410 4959
rect 13046 5039 13076 5065
rect 13145 5039 13175 5065
rect 13241 5039 13271 5065
rect 13313 5039 13343 5065
rect 13409 5039 13439 5065
rect 13498 5039 13528 5065
rect 13582 5039 13612 5065
rect 13666 5039 13696 5065
rect 13854 5039 13884 5065
rect 13938 5039 13968 5065
rect 14022 5039 14052 5065
rect 14106 5039 14136 5065
rect 14196 5039 14226 5065
rect 14295 5039 14325 5065
rect 12479 4891 12509 4913
rect 12362 4875 12416 4891
rect 12362 4841 12372 4875
rect 12406 4841 12416 4875
rect 12362 4825 12416 4841
rect 12458 4875 12512 4891
rect 12458 4841 12468 4875
rect 12502 4841 12512 4875
rect 12458 4825 12512 4841
rect 13046 4887 13076 4909
rect 13145 4895 13175 4955
rect 13046 4871 13100 4887
rect 13046 4837 13056 4871
rect 13090 4837 13100 4871
rect 12284 4764 12338 4780
rect 12284 4730 12294 4764
rect 12328 4730 12338 4764
rect 12284 4714 12338 4730
rect 12290 4677 12320 4714
rect 12380 4677 12410 4825
rect 12479 4793 12509 4825
rect 13046 4821 13100 4837
rect 13145 4879 13199 4895
rect 13145 4845 13155 4879
rect 13189 4845 13199 4879
rect 13145 4829 13199 4845
rect 13046 4789 13076 4821
rect 11230 4567 11260 4593
rect 11329 4567 11359 4593
rect 11425 4567 11455 4593
rect 11497 4567 11527 4593
rect 11593 4567 11623 4593
rect 11682 4567 11712 4593
rect 11766 4567 11796 4593
rect 11850 4567 11880 4593
rect 12038 4567 12068 4593
rect 12122 4567 12152 4593
rect 12206 4567 12236 4593
rect 12290 4567 12320 4593
rect 12380 4567 12410 4593
rect 12479 4567 12509 4593
rect 13145 4673 13175 4829
rect 13241 4783 13271 4955
rect 13217 4767 13271 4783
rect 13217 4733 13227 4767
rect 13261 4733 13271 4767
rect 13217 4717 13271 4733
rect 13241 4673 13271 4717
rect 13313 4783 13343 4955
rect 13409 4911 13439 4955
rect 13498 4911 13528 4955
rect 13582 4940 13612 4955
rect 13385 4895 13439 4911
rect 13385 4861 13395 4895
rect 13429 4861 13439 4895
rect 13385 4845 13439 4861
rect 13485 4895 13539 4911
rect 13485 4861 13495 4895
rect 13529 4861 13539 4895
rect 13485 4845 13539 4861
rect 13581 4910 13612 4940
rect 13666 4940 13696 4955
rect 13854 4940 13884 4955
rect 13666 4910 13884 4940
rect 13313 4767 13367 4783
rect 13313 4733 13323 4767
rect 13357 4733 13367 4767
rect 13313 4717 13367 4733
rect 13313 4673 13343 4717
rect 13409 4673 13439 4845
rect 13498 4673 13528 4845
rect 13581 4799 13611 4910
rect 13666 4895 13707 4910
rect 13677 4799 13707 4895
rect 13938 4880 13968 4955
rect 14022 4881 14052 4955
rect 13914 4864 13968 4880
rect 13914 4830 13924 4864
rect 13958 4830 13968 4864
rect 13914 4814 13968 4830
rect 14010 4865 14064 4881
rect 14010 4831 14020 4865
rect 14054 4831 14064 4865
rect 14010 4815 14064 4831
rect 13570 4783 13624 4799
rect 13570 4749 13580 4783
rect 13614 4749 13624 4783
rect 13570 4733 13624 4749
rect 13677 4783 13741 4799
rect 13677 4749 13697 4783
rect 13731 4749 13741 4783
rect 13582 4673 13612 4733
rect 13677 4718 13741 4749
rect 13666 4688 13884 4718
rect 13666 4673 13696 4688
rect 13854 4673 13884 4688
rect 13938 4673 13968 4814
rect 14022 4673 14052 4815
rect 14106 4776 14136 4955
rect 14196 4887 14226 4955
rect 14916 5035 14946 5061
rect 15015 5035 15045 5061
rect 15111 5035 15141 5061
rect 15183 5035 15213 5061
rect 15279 5035 15309 5061
rect 15368 5035 15398 5061
rect 15452 5035 15482 5061
rect 15536 5035 15566 5061
rect 15724 5035 15754 5061
rect 15808 5035 15838 5061
rect 15892 5035 15922 5061
rect 15976 5035 16006 5061
rect 16066 5035 16096 5061
rect 16165 5035 16195 5061
rect 14295 4887 14325 4909
rect 14178 4871 14232 4887
rect 14178 4837 14188 4871
rect 14222 4837 14232 4871
rect 14178 4821 14232 4837
rect 14274 4871 14328 4887
rect 14274 4837 14284 4871
rect 14318 4837 14328 4871
rect 14274 4821 14328 4837
rect 14916 4883 14946 4905
rect 15015 4891 15045 4951
rect 14916 4867 14970 4883
rect 14916 4833 14926 4867
rect 14960 4833 14970 4867
rect 14100 4760 14154 4776
rect 14100 4726 14110 4760
rect 14144 4726 14154 4760
rect 14100 4710 14154 4726
rect 14106 4673 14136 4710
rect 14196 4673 14226 4821
rect 14295 4789 14325 4821
rect 14916 4817 14970 4833
rect 15015 4875 15069 4891
rect 15015 4841 15025 4875
rect 15059 4841 15069 4875
rect 15015 4825 15069 4841
rect 14916 4785 14946 4817
rect 13046 4563 13076 4589
rect 13145 4563 13175 4589
rect 13241 4563 13271 4589
rect 13313 4563 13343 4589
rect 13409 4563 13439 4589
rect 13498 4563 13528 4589
rect 13582 4563 13612 4589
rect 13666 4563 13696 4589
rect 13854 4563 13884 4589
rect 13938 4563 13968 4589
rect 14022 4563 14052 4589
rect 14106 4563 14136 4589
rect 14196 4563 14226 4589
rect 14295 4563 14325 4589
rect 15015 4669 15045 4825
rect 15111 4779 15141 4951
rect 15087 4763 15141 4779
rect 15087 4729 15097 4763
rect 15131 4729 15141 4763
rect 15087 4713 15141 4729
rect 15111 4669 15141 4713
rect 15183 4779 15213 4951
rect 15279 4907 15309 4951
rect 15368 4907 15398 4951
rect 15452 4936 15482 4951
rect 15255 4891 15309 4907
rect 15255 4857 15265 4891
rect 15299 4857 15309 4891
rect 15255 4841 15309 4857
rect 15355 4891 15409 4907
rect 15355 4857 15365 4891
rect 15399 4857 15409 4891
rect 15355 4841 15409 4857
rect 15451 4906 15482 4936
rect 15536 4936 15566 4951
rect 15724 4936 15754 4951
rect 15536 4906 15754 4936
rect 15183 4763 15237 4779
rect 15183 4729 15193 4763
rect 15227 4729 15237 4763
rect 15183 4713 15237 4729
rect 15183 4669 15213 4713
rect 15279 4669 15309 4841
rect 15368 4669 15398 4841
rect 15451 4795 15481 4906
rect 15536 4891 15577 4906
rect 15547 4795 15577 4891
rect 15808 4876 15838 4951
rect 15892 4877 15922 4951
rect 15784 4860 15838 4876
rect 15784 4826 15794 4860
rect 15828 4826 15838 4860
rect 15784 4810 15838 4826
rect 15880 4861 15934 4877
rect 15880 4827 15890 4861
rect 15924 4827 15934 4861
rect 15880 4811 15934 4827
rect 15440 4779 15494 4795
rect 15440 4745 15450 4779
rect 15484 4745 15494 4779
rect 15440 4729 15494 4745
rect 15547 4779 15611 4795
rect 15547 4745 15567 4779
rect 15601 4745 15611 4779
rect 15452 4669 15482 4729
rect 15547 4714 15611 4745
rect 15536 4684 15754 4714
rect 15536 4669 15566 4684
rect 15724 4669 15754 4684
rect 15808 4669 15838 4810
rect 15892 4669 15922 4811
rect 15976 4772 16006 4951
rect 16066 4883 16096 4951
rect 16165 4883 16195 4905
rect 16048 4867 16102 4883
rect 16048 4833 16058 4867
rect 16092 4833 16102 4867
rect 16048 4817 16102 4833
rect 16144 4867 16198 4883
rect 16144 4833 16154 4867
rect 16188 4833 16198 4867
rect 16144 4817 16198 4833
rect 15970 4756 16024 4772
rect 15970 4722 15980 4756
rect 16014 4722 16024 4756
rect 15970 4706 16024 4722
rect 15976 4669 16006 4706
rect 16066 4669 16096 4817
rect 16165 4785 16195 4817
rect 14916 4559 14946 4585
rect 15015 4559 15045 4585
rect 15111 4559 15141 4585
rect 15183 4559 15213 4585
rect 15279 4559 15309 4585
rect 15368 4559 15398 4585
rect 15452 4559 15482 4585
rect 15536 4559 15566 4585
rect 15724 4559 15754 4585
rect 15808 4559 15838 4585
rect 15892 4559 15922 4585
rect 15976 4559 16006 4585
rect 16066 4559 16096 4585
rect 16165 4559 16195 4585
rect 1920 2241 1950 2267
rect 2019 2241 2049 2267
rect 2115 2241 2145 2267
rect 2187 2241 2217 2267
rect 2283 2241 2313 2267
rect 2372 2241 2402 2267
rect 2456 2241 2486 2267
rect 2540 2241 2570 2267
rect 2728 2241 2758 2267
rect 2812 2241 2842 2267
rect 2896 2241 2926 2267
rect 2980 2241 3010 2267
rect 3070 2241 3100 2267
rect 3169 2241 3199 2267
rect 1920 2089 1950 2111
rect 2019 2097 2049 2157
rect 1920 2073 1974 2089
rect 1920 2039 1930 2073
rect 1964 2039 1974 2073
rect 1920 2023 1974 2039
rect 2019 2081 2073 2097
rect 2019 2047 2029 2081
rect 2063 2047 2073 2081
rect 2019 2031 2073 2047
rect 1920 1991 1950 2023
rect 2019 1875 2049 2031
rect 2115 1985 2145 2157
rect 2091 1969 2145 1985
rect 2091 1935 2101 1969
rect 2135 1935 2145 1969
rect 2091 1919 2145 1935
rect 2115 1875 2145 1919
rect 2187 1985 2217 2157
rect 2283 2113 2313 2157
rect 2372 2113 2402 2157
rect 2456 2142 2486 2157
rect 2259 2097 2313 2113
rect 2259 2063 2269 2097
rect 2303 2063 2313 2097
rect 2259 2047 2313 2063
rect 2359 2097 2413 2113
rect 2359 2063 2369 2097
rect 2403 2063 2413 2097
rect 2359 2047 2413 2063
rect 2455 2112 2486 2142
rect 2540 2142 2570 2157
rect 2728 2142 2758 2157
rect 2540 2112 2758 2142
rect 2187 1969 2241 1985
rect 2187 1935 2197 1969
rect 2231 1935 2241 1969
rect 2187 1919 2241 1935
rect 2187 1875 2217 1919
rect 2283 1875 2313 2047
rect 2372 1875 2402 2047
rect 2455 2001 2485 2112
rect 2540 2097 2581 2112
rect 2551 2001 2581 2097
rect 2812 2082 2842 2157
rect 2896 2083 2926 2157
rect 2788 2066 2842 2082
rect 2788 2032 2798 2066
rect 2832 2032 2842 2066
rect 2788 2016 2842 2032
rect 2884 2067 2938 2083
rect 2884 2033 2894 2067
rect 2928 2033 2938 2067
rect 2884 2017 2938 2033
rect 2444 1985 2498 2001
rect 2444 1951 2454 1985
rect 2488 1951 2498 1985
rect 2444 1935 2498 1951
rect 2551 1985 2615 2001
rect 2551 1951 2571 1985
rect 2605 1951 2615 1985
rect 2456 1875 2486 1935
rect 2551 1920 2615 1951
rect 2540 1890 2758 1920
rect 2540 1875 2570 1890
rect 2728 1875 2758 1890
rect 2812 1875 2842 2016
rect 2896 1875 2926 2017
rect 2980 1978 3010 2157
rect 3070 2089 3100 2157
rect 3790 2237 3820 2263
rect 3889 2237 3919 2263
rect 3985 2237 4015 2263
rect 4057 2237 4087 2263
rect 4153 2237 4183 2263
rect 4242 2237 4272 2263
rect 4326 2237 4356 2263
rect 4410 2237 4440 2263
rect 4598 2237 4628 2263
rect 4682 2237 4712 2263
rect 4766 2237 4796 2263
rect 4850 2237 4880 2263
rect 4940 2237 4970 2263
rect 5039 2237 5069 2263
rect 3169 2089 3199 2111
rect 3052 2073 3106 2089
rect 3052 2039 3062 2073
rect 3096 2039 3106 2073
rect 3052 2023 3106 2039
rect 3148 2073 3202 2089
rect 3148 2039 3158 2073
rect 3192 2039 3202 2073
rect 3148 2023 3202 2039
rect 3790 2085 3820 2107
rect 3889 2093 3919 2153
rect 3790 2069 3844 2085
rect 3790 2035 3800 2069
rect 3834 2035 3844 2069
rect 2974 1962 3028 1978
rect 2974 1928 2984 1962
rect 3018 1928 3028 1962
rect 2974 1912 3028 1928
rect 2980 1875 3010 1912
rect 3070 1875 3100 2023
rect 3169 1991 3199 2023
rect 3790 2019 3844 2035
rect 3889 2077 3943 2093
rect 3889 2043 3899 2077
rect 3933 2043 3943 2077
rect 3889 2027 3943 2043
rect 3790 1987 3820 2019
rect 1920 1765 1950 1791
rect 2019 1765 2049 1791
rect 2115 1765 2145 1791
rect 2187 1765 2217 1791
rect 2283 1765 2313 1791
rect 2372 1765 2402 1791
rect 2456 1765 2486 1791
rect 2540 1765 2570 1791
rect 2728 1765 2758 1791
rect 2812 1765 2842 1791
rect 2896 1765 2926 1791
rect 2980 1765 3010 1791
rect 3070 1765 3100 1791
rect 3169 1765 3199 1791
rect 3889 1871 3919 2027
rect 3985 1981 4015 2153
rect 3961 1965 4015 1981
rect 3961 1931 3971 1965
rect 4005 1931 4015 1965
rect 3961 1915 4015 1931
rect 3985 1871 4015 1915
rect 4057 1981 4087 2153
rect 4153 2109 4183 2153
rect 4242 2109 4272 2153
rect 4326 2138 4356 2153
rect 4129 2093 4183 2109
rect 4129 2059 4139 2093
rect 4173 2059 4183 2093
rect 4129 2043 4183 2059
rect 4229 2093 4283 2109
rect 4229 2059 4239 2093
rect 4273 2059 4283 2093
rect 4229 2043 4283 2059
rect 4325 2108 4356 2138
rect 4410 2138 4440 2153
rect 4598 2138 4628 2153
rect 4410 2108 4628 2138
rect 4057 1965 4111 1981
rect 4057 1931 4067 1965
rect 4101 1931 4111 1965
rect 4057 1915 4111 1931
rect 4057 1871 4087 1915
rect 4153 1871 4183 2043
rect 4242 1871 4272 2043
rect 4325 1997 4355 2108
rect 4410 2093 4451 2108
rect 4421 1997 4451 2093
rect 4682 2078 4712 2153
rect 4766 2079 4796 2153
rect 4658 2062 4712 2078
rect 4658 2028 4668 2062
rect 4702 2028 4712 2062
rect 4658 2012 4712 2028
rect 4754 2063 4808 2079
rect 4754 2029 4764 2063
rect 4798 2029 4808 2063
rect 4754 2013 4808 2029
rect 4314 1981 4368 1997
rect 4314 1947 4324 1981
rect 4358 1947 4368 1981
rect 4314 1931 4368 1947
rect 4421 1981 4485 1997
rect 4421 1947 4441 1981
rect 4475 1947 4485 1981
rect 4326 1871 4356 1931
rect 4421 1916 4485 1947
rect 4410 1886 4628 1916
rect 4410 1871 4440 1886
rect 4598 1871 4628 1886
rect 4682 1871 4712 2012
rect 4766 1871 4796 2013
rect 4850 1974 4880 2153
rect 4940 2085 4970 2153
rect 5606 2233 5636 2259
rect 5705 2233 5735 2259
rect 5801 2233 5831 2259
rect 5873 2233 5903 2259
rect 5969 2233 5999 2259
rect 6058 2233 6088 2259
rect 6142 2233 6172 2259
rect 6226 2233 6256 2259
rect 6414 2233 6444 2259
rect 6498 2233 6528 2259
rect 6582 2233 6612 2259
rect 6666 2233 6696 2259
rect 6756 2233 6786 2259
rect 6855 2233 6885 2259
rect 5039 2085 5069 2107
rect 4922 2069 4976 2085
rect 4922 2035 4932 2069
rect 4966 2035 4976 2069
rect 4922 2019 4976 2035
rect 5018 2069 5072 2085
rect 5018 2035 5028 2069
rect 5062 2035 5072 2069
rect 5018 2019 5072 2035
rect 5606 2081 5636 2103
rect 5705 2089 5735 2149
rect 5606 2065 5660 2081
rect 5606 2031 5616 2065
rect 5650 2031 5660 2065
rect 4844 1958 4898 1974
rect 4844 1924 4854 1958
rect 4888 1924 4898 1958
rect 4844 1908 4898 1924
rect 4850 1871 4880 1908
rect 4940 1871 4970 2019
rect 5039 1987 5069 2019
rect 5606 2015 5660 2031
rect 5705 2073 5759 2089
rect 5705 2039 5715 2073
rect 5749 2039 5759 2073
rect 5705 2023 5759 2039
rect 5606 1983 5636 2015
rect 3790 1761 3820 1787
rect 3889 1761 3919 1787
rect 3985 1761 4015 1787
rect 4057 1761 4087 1787
rect 4153 1761 4183 1787
rect 4242 1761 4272 1787
rect 4326 1761 4356 1787
rect 4410 1761 4440 1787
rect 4598 1761 4628 1787
rect 4682 1761 4712 1787
rect 4766 1761 4796 1787
rect 4850 1761 4880 1787
rect 4940 1761 4970 1787
rect 5039 1761 5069 1787
rect 5705 1867 5735 2023
rect 5801 1977 5831 2149
rect 5777 1961 5831 1977
rect 5777 1927 5787 1961
rect 5821 1927 5831 1961
rect 5777 1911 5831 1927
rect 5801 1867 5831 1911
rect 5873 1977 5903 2149
rect 5969 2105 5999 2149
rect 6058 2105 6088 2149
rect 6142 2134 6172 2149
rect 5945 2089 5999 2105
rect 5945 2055 5955 2089
rect 5989 2055 5999 2089
rect 5945 2039 5999 2055
rect 6045 2089 6099 2105
rect 6045 2055 6055 2089
rect 6089 2055 6099 2089
rect 6045 2039 6099 2055
rect 6141 2104 6172 2134
rect 6226 2134 6256 2149
rect 6414 2134 6444 2149
rect 6226 2104 6444 2134
rect 5873 1961 5927 1977
rect 5873 1927 5883 1961
rect 5917 1927 5927 1961
rect 5873 1911 5927 1927
rect 5873 1867 5903 1911
rect 5969 1867 5999 2039
rect 6058 1867 6088 2039
rect 6141 1993 6171 2104
rect 6226 2089 6267 2104
rect 6237 1993 6267 2089
rect 6498 2074 6528 2149
rect 6582 2075 6612 2149
rect 6474 2058 6528 2074
rect 6474 2024 6484 2058
rect 6518 2024 6528 2058
rect 6474 2008 6528 2024
rect 6570 2059 6624 2075
rect 6570 2025 6580 2059
rect 6614 2025 6624 2059
rect 6570 2009 6624 2025
rect 6130 1977 6184 1993
rect 6130 1943 6140 1977
rect 6174 1943 6184 1977
rect 6130 1927 6184 1943
rect 6237 1977 6301 1993
rect 6237 1943 6257 1977
rect 6291 1943 6301 1977
rect 6142 1867 6172 1927
rect 6237 1912 6301 1943
rect 6226 1882 6444 1912
rect 6226 1867 6256 1882
rect 6414 1867 6444 1882
rect 6498 1867 6528 2008
rect 6582 1867 6612 2009
rect 6666 1970 6696 2149
rect 6756 2081 6786 2149
rect 7476 2229 7506 2255
rect 7575 2229 7605 2255
rect 7671 2229 7701 2255
rect 7743 2229 7773 2255
rect 7839 2229 7869 2255
rect 7928 2229 7958 2255
rect 8012 2229 8042 2255
rect 8096 2229 8126 2255
rect 8284 2229 8314 2255
rect 8368 2229 8398 2255
rect 8452 2229 8482 2255
rect 8536 2229 8566 2255
rect 8626 2229 8656 2255
rect 8725 2229 8755 2255
rect 6855 2081 6885 2103
rect 6738 2065 6792 2081
rect 6738 2031 6748 2065
rect 6782 2031 6792 2065
rect 6738 2015 6792 2031
rect 6834 2065 6888 2081
rect 6834 2031 6844 2065
rect 6878 2031 6888 2065
rect 6834 2015 6888 2031
rect 7476 2077 7506 2099
rect 7575 2085 7605 2145
rect 7476 2061 7530 2077
rect 7476 2027 7486 2061
rect 7520 2027 7530 2061
rect 6660 1954 6714 1970
rect 6660 1920 6670 1954
rect 6704 1920 6714 1954
rect 6660 1904 6714 1920
rect 6666 1867 6696 1904
rect 6756 1867 6786 2015
rect 6855 1983 6885 2015
rect 7476 2011 7530 2027
rect 7575 2069 7629 2085
rect 7575 2035 7585 2069
rect 7619 2035 7629 2069
rect 7575 2019 7629 2035
rect 7476 1979 7506 2011
rect 5606 1757 5636 1783
rect 5705 1757 5735 1783
rect 5801 1757 5831 1783
rect 5873 1757 5903 1783
rect 5969 1757 5999 1783
rect 6058 1757 6088 1783
rect 6142 1757 6172 1783
rect 6226 1757 6256 1783
rect 6414 1757 6444 1783
rect 6498 1757 6528 1783
rect 6582 1757 6612 1783
rect 6666 1757 6696 1783
rect 6756 1757 6786 1783
rect 6855 1757 6885 1783
rect 7575 1863 7605 2019
rect 7671 1973 7701 2145
rect 7647 1957 7701 1973
rect 7647 1923 7657 1957
rect 7691 1923 7701 1957
rect 7647 1907 7701 1923
rect 7671 1863 7701 1907
rect 7743 1973 7773 2145
rect 7839 2101 7869 2145
rect 7928 2101 7958 2145
rect 8012 2130 8042 2145
rect 7815 2085 7869 2101
rect 7815 2051 7825 2085
rect 7859 2051 7869 2085
rect 7815 2035 7869 2051
rect 7915 2085 7969 2101
rect 7915 2051 7925 2085
rect 7959 2051 7969 2085
rect 7915 2035 7969 2051
rect 8011 2100 8042 2130
rect 8096 2130 8126 2145
rect 8284 2130 8314 2145
rect 8096 2100 8314 2130
rect 7743 1957 7797 1973
rect 7743 1923 7753 1957
rect 7787 1923 7797 1957
rect 7743 1907 7797 1923
rect 7743 1863 7773 1907
rect 7839 1863 7869 2035
rect 7928 1863 7958 2035
rect 8011 1989 8041 2100
rect 8096 2085 8137 2100
rect 8107 1989 8137 2085
rect 8368 2070 8398 2145
rect 8452 2071 8482 2145
rect 8344 2054 8398 2070
rect 8344 2020 8354 2054
rect 8388 2020 8398 2054
rect 8344 2004 8398 2020
rect 8440 2055 8494 2071
rect 8440 2021 8450 2055
rect 8484 2021 8494 2055
rect 8440 2005 8494 2021
rect 8000 1973 8054 1989
rect 8000 1939 8010 1973
rect 8044 1939 8054 1973
rect 8000 1923 8054 1939
rect 8107 1973 8171 1989
rect 8107 1939 8127 1973
rect 8161 1939 8171 1973
rect 8012 1863 8042 1923
rect 8107 1908 8171 1939
rect 8096 1878 8314 1908
rect 8096 1863 8126 1878
rect 8284 1863 8314 1878
rect 8368 1863 8398 2004
rect 8452 1863 8482 2005
rect 8536 1966 8566 2145
rect 8626 2077 8656 2145
rect 9290 2227 9320 2253
rect 9389 2227 9419 2253
rect 9485 2227 9515 2253
rect 9557 2227 9587 2253
rect 9653 2227 9683 2253
rect 9742 2227 9772 2253
rect 9826 2227 9856 2253
rect 9910 2227 9940 2253
rect 10098 2227 10128 2253
rect 10182 2227 10212 2253
rect 10266 2227 10296 2253
rect 10350 2227 10380 2253
rect 10440 2227 10470 2253
rect 10539 2227 10569 2253
rect 8725 2077 8755 2099
rect 8608 2061 8662 2077
rect 8608 2027 8618 2061
rect 8652 2027 8662 2061
rect 8608 2011 8662 2027
rect 8704 2061 8758 2077
rect 8704 2027 8714 2061
rect 8748 2027 8758 2061
rect 8704 2011 8758 2027
rect 9290 2075 9320 2097
rect 9389 2083 9419 2143
rect 9290 2059 9344 2075
rect 9290 2025 9300 2059
rect 9334 2025 9344 2059
rect 8530 1950 8584 1966
rect 8530 1916 8540 1950
rect 8574 1916 8584 1950
rect 8530 1900 8584 1916
rect 8536 1863 8566 1900
rect 8626 1863 8656 2011
rect 8725 1979 8755 2011
rect 9290 2009 9344 2025
rect 9389 2067 9443 2083
rect 9389 2033 9399 2067
rect 9433 2033 9443 2067
rect 9389 2017 9443 2033
rect 9290 1977 9320 2009
rect 7476 1753 7506 1779
rect 7575 1753 7605 1779
rect 7671 1753 7701 1779
rect 7743 1753 7773 1779
rect 7839 1753 7869 1779
rect 7928 1753 7958 1779
rect 8012 1753 8042 1779
rect 8096 1753 8126 1779
rect 8284 1753 8314 1779
rect 8368 1753 8398 1779
rect 8452 1753 8482 1779
rect 8536 1753 8566 1779
rect 8626 1753 8656 1779
rect 8725 1753 8755 1779
rect 9389 1861 9419 2017
rect 9485 1971 9515 2143
rect 9461 1955 9515 1971
rect 9461 1921 9471 1955
rect 9505 1921 9515 1955
rect 9461 1905 9515 1921
rect 9485 1861 9515 1905
rect 9557 1971 9587 2143
rect 9653 2099 9683 2143
rect 9742 2099 9772 2143
rect 9826 2128 9856 2143
rect 9629 2083 9683 2099
rect 9629 2049 9639 2083
rect 9673 2049 9683 2083
rect 9629 2033 9683 2049
rect 9729 2083 9783 2099
rect 9729 2049 9739 2083
rect 9773 2049 9783 2083
rect 9729 2033 9783 2049
rect 9825 2098 9856 2128
rect 9910 2128 9940 2143
rect 10098 2128 10128 2143
rect 9910 2098 10128 2128
rect 9557 1955 9611 1971
rect 9557 1921 9567 1955
rect 9601 1921 9611 1955
rect 9557 1905 9611 1921
rect 9557 1861 9587 1905
rect 9653 1861 9683 2033
rect 9742 1861 9772 2033
rect 9825 1987 9855 2098
rect 9910 2083 9951 2098
rect 9921 1987 9951 2083
rect 10182 2068 10212 2143
rect 10266 2069 10296 2143
rect 10158 2052 10212 2068
rect 10158 2018 10168 2052
rect 10202 2018 10212 2052
rect 10158 2002 10212 2018
rect 10254 2053 10308 2069
rect 10254 2019 10264 2053
rect 10298 2019 10308 2053
rect 10254 2003 10308 2019
rect 9814 1971 9868 1987
rect 9814 1937 9824 1971
rect 9858 1937 9868 1971
rect 9814 1921 9868 1937
rect 9921 1971 9985 1987
rect 9921 1937 9941 1971
rect 9975 1937 9985 1971
rect 9826 1861 9856 1921
rect 9921 1906 9985 1937
rect 9910 1876 10128 1906
rect 9910 1861 9940 1876
rect 10098 1861 10128 1876
rect 10182 1861 10212 2002
rect 10266 1861 10296 2003
rect 10350 1964 10380 2143
rect 10440 2075 10470 2143
rect 11160 2223 11190 2249
rect 11259 2223 11289 2249
rect 11355 2223 11385 2249
rect 11427 2223 11457 2249
rect 11523 2223 11553 2249
rect 11612 2223 11642 2249
rect 11696 2223 11726 2249
rect 11780 2223 11810 2249
rect 11968 2223 11998 2249
rect 12052 2223 12082 2249
rect 12136 2223 12166 2249
rect 12220 2223 12250 2249
rect 12310 2223 12340 2249
rect 12409 2223 12439 2249
rect 10539 2075 10569 2097
rect 10422 2059 10476 2075
rect 10422 2025 10432 2059
rect 10466 2025 10476 2059
rect 10422 2009 10476 2025
rect 10518 2059 10572 2075
rect 10518 2025 10528 2059
rect 10562 2025 10572 2059
rect 10518 2009 10572 2025
rect 11160 2071 11190 2093
rect 11259 2079 11289 2139
rect 11160 2055 11214 2071
rect 11160 2021 11170 2055
rect 11204 2021 11214 2055
rect 10344 1948 10398 1964
rect 10344 1914 10354 1948
rect 10388 1914 10398 1948
rect 10344 1898 10398 1914
rect 10350 1861 10380 1898
rect 10440 1861 10470 2009
rect 10539 1977 10569 2009
rect 11160 2005 11214 2021
rect 11259 2063 11313 2079
rect 11259 2029 11269 2063
rect 11303 2029 11313 2063
rect 11259 2013 11313 2029
rect 11160 1973 11190 2005
rect 9290 1751 9320 1777
rect 9389 1751 9419 1777
rect 9485 1751 9515 1777
rect 9557 1751 9587 1777
rect 9653 1751 9683 1777
rect 9742 1751 9772 1777
rect 9826 1751 9856 1777
rect 9910 1751 9940 1777
rect 10098 1751 10128 1777
rect 10182 1751 10212 1777
rect 10266 1751 10296 1777
rect 10350 1751 10380 1777
rect 10440 1751 10470 1777
rect 10539 1751 10569 1777
rect 11259 1857 11289 2013
rect 11355 1967 11385 2139
rect 11331 1951 11385 1967
rect 11331 1917 11341 1951
rect 11375 1917 11385 1951
rect 11331 1901 11385 1917
rect 11355 1857 11385 1901
rect 11427 1967 11457 2139
rect 11523 2095 11553 2139
rect 11612 2095 11642 2139
rect 11696 2124 11726 2139
rect 11499 2079 11553 2095
rect 11499 2045 11509 2079
rect 11543 2045 11553 2079
rect 11499 2029 11553 2045
rect 11599 2079 11653 2095
rect 11599 2045 11609 2079
rect 11643 2045 11653 2079
rect 11599 2029 11653 2045
rect 11695 2094 11726 2124
rect 11780 2124 11810 2139
rect 11968 2124 11998 2139
rect 11780 2094 11998 2124
rect 11427 1951 11481 1967
rect 11427 1917 11437 1951
rect 11471 1917 11481 1951
rect 11427 1901 11481 1917
rect 11427 1857 11457 1901
rect 11523 1857 11553 2029
rect 11612 1857 11642 2029
rect 11695 1983 11725 2094
rect 11780 2079 11821 2094
rect 11791 1983 11821 2079
rect 12052 2064 12082 2139
rect 12136 2065 12166 2139
rect 12028 2048 12082 2064
rect 12028 2014 12038 2048
rect 12072 2014 12082 2048
rect 12028 1998 12082 2014
rect 12124 2049 12178 2065
rect 12124 2015 12134 2049
rect 12168 2015 12178 2049
rect 12124 1999 12178 2015
rect 11684 1967 11738 1983
rect 11684 1933 11694 1967
rect 11728 1933 11738 1967
rect 11684 1917 11738 1933
rect 11791 1967 11855 1983
rect 11791 1933 11811 1967
rect 11845 1933 11855 1967
rect 11696 1857 11726 1917
rect 11791 1902 11855 1933
rect 11780 1872 11998 1902
rect 11780 1857 11810 1872
rect 11968 1857 11998 1872
rect 12052 1857 12082 1998
rect 12136 1857 12166 1999
rect 12220 1960 12250 2139
rect 12310 2071 12340 2139
rect 12976 2219 13006 2245
rect 13075 2219 13105 2245
rect 13171 2219 13201 2245
rect 13243 2219 13273 2245
rect 13339 2219 13369 2245
rect 13428 2219 13458 2245
rect 13512 2219 13542 2245
rect 13596 2219 13626 2245
rect 13784 2219 13814 2245
rect 13868 2219 13898 2245
rect 13952 2219 13982 2245
rect 14036 2219 14066 2245
rect 14126 2219 14156 2245
rect 14225 2219 14255 2245
rect 12409 2071 12439 2093
rect 12292 2055 12346 2071
rect 12292 2021 12302 2055
rect 12336 2021 12346 2055
rect 12292 2005 12346 2021
rect 12388 2055 12442 2071
rect 12388 2021 12398 2055
rect 12432 2021 12442 2055
rect 12388 2005 12442 2021
rect 12976 2067 13006 2089
rect 13075 2075 13105 2135
rect 12976 2051 13030 2067
rect 12976 2017 12986 2051
rect 13020 2017 13030 2051
rect 12214 1944 12268 1960
rect 12214 1910 12224 1944
rect 12258 1910 12268 1944
rect 12214 1894 12268 1910
rect 12220 1857 12250 1894
rect 12310 1857 12340 2005
rect 12409 1973 12439 2005
rect 12976 2001 13030 2017
rect 13075 2059 13129 2075
rect 13075 2025 13085 2059
rect 13119 2025 13129 2059
rect 13075 2009 13129 2025
rect 12976 1969 13006 2001
rect 11160 1747 11190 1773
rect 11259 1747 11289 1773
rect 11355 1747 11385 1773
rect 11427 1747 11457 1773
rect 11523 1747 11553 1773
rect 11612 1747 11642 1773
rect 11696 1747 11726 1773
rect 11780 1747 11810 1773
rect 11968 1747 11998 1773
rect 12052 1747 12082 1773
rect 12136 1747 12166 1773
rect 12220 1747 12250 1773
rect 12310 1747 12340 1773
rect 12409 1747 12439 1773
rect 13075 1853 13105 2009
rect 13171 1963 13201 2135
rect 13147 1947 13201 1963
rect 13147 1913 13157 1947
rect 13191 1913 13201 1947
rect 13147 1897 13201 1913
rect 13171 1853 13201 1897
rect 13243 1963 13273 2135
rect 13339 2091 13369 2135
rect 13428 2091 13458 2135
rect 13512 2120 13542 2135
rect 13315 2075 13369 2091
rect 13315 2041 13325 2075
rect 13359 2041 13369 2075
rect 13315 2025 13369 2041
rect 13415 2075 13469 2091
rect 13415 2041 13425 2075
rect 13459 2041 13469 2075
rect 13415 2025 13469 2041
rect 13511 2090 13542 2120
rect 13596 2120 13626 2135
rect 13784 2120 13814 2135
rect 13596 2090 13814 2120
rect 13243 1947 13297 1963
rect 13243 1913 13253 1947
rect 13287 1913 13297 1947
rect 13243 1897 13297 1913
rect 13243 1853 13273 1897
rect 13339 1853 13369 2025
rect 13428 1853 13458 2025
rect 13511 1979 13541 2090
rect 13596 2075 13637 2090
rect 13607 1979 13637 2075
rect 13868 2060 13898 2135
rect 13952 2061 13982 2135
rect 13844 2044 13898 2060
rect 13844 2010 13854 2044
rect 13888 2010 13898 2044
rect 13844 1994 13898 2010
rect 13940 2045 13994 2061
rect 13940 2011 13950 2045
rect 13984 2011 13994 2045
rect 13940 1995 13994 2011
rect 13500 1963 13554 1979
rect 13500 1929 13510 1963
rect 13544 1929 13554 1963
rect 13500 1913 13554 1929
rect 13607 1963 13671 1979
rect 13607 1929 13627 1963
rect 13661 1929 13671 1963
rect 13512 1853 13542 1913
rect 13607 1898 13671 1929
rect 13596 1868 13814 1898
rect 13596 1853 13626 1868
rect 13784 1853 13814 1868
rect 13868 1853 13898 1994
rect 13952 1853 13982 1995
rect 14036 1956 14066 2135
rect 14126 2067 14156 2135
rect 14846 2215 14876 2241
rect 14945 2215 14975 2241
rect 15041 2215 15071 2241
rect 15113 2215 15143 2241
rect 15209 2215 15239 2241
rect 15298 2215 15328 2241
rect 15382 2215 15412 2241
rect 15466 2215 15496 2241
rect 15654 2215 15684 2241
rect 15738 2215 15768 2241
rect 15822 2215 15852 2241
rect 15906 2215 15936 2241
rect 15996 2215 16026 2241
rect 16095 2215 16125 2241
rect 14225 2067 14255 2089
rect 14108 2051 14162 2067
rect 14108 2017 14118 2051
rect 14152 2017 14162 2051
rect 14108 2001 14162 2017
rect 14204 2051 14258 2067
rect 14204 2017 14214 2051
rect 14248 2017 14258 2051
rect 14204 2001 14258 2017
rect 14846 2063 14876 2085
rect 14945 2071 14975 2131
rect 14846 2047 14900 2063
rect 14846 2013 14856 2047
rect 14890 2013 14900 2047
rect 14030 1940 14084 1956
rect 14030 1906 14040 1940
rect 14074 1906 14084 1940
rect 14030 1890 14084 1906
rect 14036 1853 14066 1890
rect 14126 1853 14156 2001
rect 14225 1969 14255 2001
rect 14846 1997 14900 2013
rect 14945 2055 14999 2071
rect 14945 2021 14955 2055
rect 14989 2021 14999 2055
rect 14945 2005 14999 2021
rect 14846 1965 14876 1997
rect 12976 1743 13006 1769
rect 13075 1743 13105 1769
rect 13171 1743 13201 1769
rect 13243 1743 13273 1769
rect 13339 1743 13369 1769
rect 13428 1743 13458 1769
rect 13512 1743 13542 1769
rect 13596 1743 13626 1769
rect 13784 1743 13814 1769
rect 13868 1743 13898 1769
rect 13952 1743 13982 1769
rect 14036 1743 14066 1769
rect 14126 1743 14156 1769
rect 14225 1743 14255 1769
rect 14945 1849 14975 2005
rect 15041 1959 15071 2131
rect 15017 1943 15071 1959
rect 15017 1909 15027 1943
rect 15061 1909 15071 1943
rect 15017 1893 15071 1909
rect 15041 1849 15071 1893
rect 15113 1959 15143 2131
rect 15209 2087 15239 2131
rect 15298 2087 15328 2131
rect 15382 2116 15412 2131
rect 15185 2071 15239 2087
rect 15185 2037 15195 2071
rect 15229 2037 15239 2071
rect 15185 2021 15239 2037
rect 15285 2071 15339 2087
rect 15285 2037 15295 2071
rect 15329 2037 15339 2071
rect 15285 2021 15339 2037
rect 15381 2086 15412 2116
rect 15466 2116 15496 2131
rect 15654 2116 15684 2131
rect 15466 2086 15684 2116
rect 15113 1943 15167 1959
rect 15113 1909 15123 1943
rect 15157 1909 15167 1943
rect 15113 1893 15167 1909
rect 15113 1849 15143 1893
rect 15209 1849 15239 2021
rect 15298 1849 15328 2021
rect 15381 1975 15411 2086
rect 15466 2071 15507 2086
rect 15477 1975 15507 2071
rect 15738 2056 15768 2131
rect 15822 2057 15852 2131
rect 15714 2040 15768 2056
rect 15714 2006 15724 2040
rect 15758 2006 15768 2040
rect 15714 1990 15768 2006
rect 15810 2041 15864 2057
rect 15810 2007 15820 2041
rect 15854 2007 15864 2041
rect 15810 1991 15864 2007
rect 15370 1959 15424 1975
rect 15370 1925 15380 1959
rect 15414 1925 15424 1959
rect 15370 1909 15424 1925
rect 15477 1959 15541 1975
rect 15477 1925 15497 1959
rect 15531 1925 15541 1959
rect 15382 1849 15412 1909
rect 15477 1894 15541 1925
rect 15466 1864 15684 1894
rect 15466 1849 15496 1864
rect 15654 1849 15684 1864
rect 15738 1849 15768 1990
rect 15822 1849 15852 1991
rect 15906 1952 15936 2131
rect 15996 2063 16026 2131
rect 16095 2063 16125 2085
rect 15978 2047 16032 2063
rect 15978 2013 15988 2047
rect 16022 2013 16032 2047
rect 15978 1997 16032 2013
rect 16074 2047 16128 2063
rect 16074 2013 16084 2047
rect 16118 2013 16128 2047
rect 16074 1997 16128 2013
rect 15900 1936 15954 1952
rect 15900 1902 15910 1936
rect 15944 1902 15954 1936
rect 15900 1886 15954 1902
rect 15906 1849 15936 1886
rect 15996 1849 16026 1997
rect 16095 1965 16125 1997
rect 14846 1739 14876 1765
rect 14945 1739 14975 1765
rect 15041 1739 15071 1765
rect 15113 1739 15143 1765
rect 15209 1739 15239 1765
rect 15298 1739 15328 1765
rect 15382 1739 15412 1765
rect 15466 1739 15496 1765
rect 15654 1739 15684 1765
rect 15738 1739 15768 1765
rect 15822 1739 15852 1765
rect 15906 1739 15936 1765
rect 15996 1739 16026 1765
rect 16095 1739 16125 1765
<< polycont >>
rect 9515 16241 9549 16275
rect 9632 16241 9666 16275
rect 9767 16241 9801 16275
rect 9863 16241 9897 16275
rect 9602 15497 9636 15531
rect 9743 15497 9777 15531
rect 9851 15497 9885 15531
rect 11601 15387 11635 15421
rect 11747 15387 11781 15421
rect 11853 15387 11887 15421
rect 11949 15387 11983 15421
rect 12060 15387 12094 15421
rect 10786 14887 10820 14921
rect 10927 14887 10961 14921
rect 11035 14887 11069 14921
rect 9525 14677 9559 14711
rect 9642 14677 9676 14711
rect 9777 14677 9811 14711
rect 9873 14677 9907 14711
rect 9612 13933 9646 13967
rect 9753 13933 9787 13967
rect 12861 14129 12895 14163
rect 9861 13933 9895 13967
rect 10817 13921 10851 13955
rect 10963 13921 10997 13955
rect 11069 13921 11103 13955
rect 11165 13921 11199 13955
rect 11276 13921 11310 13955
rect 12639 13905 12673 13939
rect 12765 13905 12799 13939
rect 12941 13905 12975 13939
rect 13037 13905 13071 13939
rect 11822 13547 11856 13581
rect 11958 13547 11992 13581
rect 12061 13547 12095 13581
rect 11083 13306 11117 13340
rect 9517 13009 9551 13043
rect 9634 13009 9668 13043
rect 9769 13009 9803 13043
rect 9865 13009 9899 13043
rect 10945 13033 10979 13067
rect 11155 13073 11189 13107
rect 11251 13079 11285 13113
rect 9604 12265 9638 12299
rect 9745 12265 9779 12299
rect 9853 12265 9887 12299
rect 10980 12059 11014 12093
rect 11121 12059 11155 12093
rect 11229 12059 11263 12093
rect 9527 11445 9561 11479
rect 9644 11445 9678 11479
rect 9779 11445 9813 11479
rect 9875 11445 9909 11479
rect 9614 10701 9648 10735
rect 9755 10701 9789 10735
rect 9863 10701 9897 10735
rect 6274 6351 6308 6385
rect 9342 5719 9376 5753
rect 9441 5727 9475 5761
rect 1960 5299 1994 5333
rect 2059 5307 2093 5341
rect 2131 5195 2165 5229
rect 2299 5323 2333 5357
rect 2399 5323 2433 5357
rect 2227 5195 2261 5229
rect 2828 5292 2862 5326
rect 2924 5293 2958 5327
rect 2484 5211 2518 5245
rect 2601 5211 2635 5245
rect 3092 5299 3126 5333
rect 3188 5299 3222 5333
rect 3830 5295 3864 5329
rect 3014 5188 3048 5222
rect 3929 5303 3963 5337
rect 4001 5191 4035 5225
rect 4169 5319 4203 5353
rect 4269 5319 4303 5353
rect 4097 5191 4131 5225
rect 4698 5288 4732 5322
rect 4794 5289 4828 5323
rect 4354 5207 4388 5241
rect 4471 5207 4505 5241
rect 4962 5295 4996 5329
rect 5058 5295 5092 5329
rect 5646 5291 5680 5325
rect 4884 5184 4918 5218
rect 5745 5299 5779 5333
rect 5817 5187 5851 5221
rect 5985 5315 6019 5349
rect 6085 5315 6119 5349
rect 5913 5187 5947 5221
rect 6514 5284 6548 5318
rect 6610 5285 6644 5319
rect 6170 5203 6204 5237
rect 6287 5203 6321 5237
rect 6778 5291 6812 5325
rect 6874 5291 6908 5325
rect 7516 5287 7550 5321
rect 6700 5180 6734 5214
rect 7615 5295 7649 5329
rect 7687 5183 7721 5217
rect 7855 5311 7889 5345
rect 7955 5311 7989 5345
rect 7783 5183 7817 5217
rect 8384 5280 8418 5314
rect 8480 5281 8514 5315
rect 8040 5199 8074 5233
rect 8157 5199 8191 5233
rect 9513 5615 9547 5649
rect 9681 5743 9715 5777
rect 9781 5743 9815 5777
rect 9609 5615 9643 5649
rect 10210 5712 10244 5746
rect 10306 5713 10340 5747
rect 9866 5631 9900 5665
rect 9983 5631 10017 5665
rect 10474 5719 10508 5753
rect 10570 5719 10604 5753
rect 11212 5715 11246 5749
rect 10396 5608 10430 5642
rect 11311 5723 11345 5757
rect 11383 5611 11417 5645
rect 11551 5739 11585 5773
rect 11651 5739 11685 5773
rect 11479 5611 11513 5645
rect 12080 5708 12114 5742
rect 12176 5709 12210 5743
rect 11736 5627 11770 5661
rect 11853 5627 11887 5661
rect 12344 5715 12378 5749
rect 12440 5715 12474 5749
rect 13028 5711 13062 5745
rect 12266 5604 12300 5638
rect 13127 5719 13161 5753
rect 13199 5607 13233 5641
rect 13367 5735 13401 5769
rect 13467 5735 13501 5769
rect 13295 5607 13329 5641
rect 13896 5704 13930 5738
rect 13992 5705 14026 5739
rect 13552 5623 13586 5657
rect 13669 5623 13703 5657
rect 14160 5711 14194 5745
rect 14256 5711 14290 5745
rect 14898 5707 14932 5741
rect 14082 5600 14116 5634
rect 14997 5715 15031 5749
rect 15069 5603 15103 5637
rect 15237 5731 15271 5765
rect 15337 5731 15371 5765
rect 15165 5603 15199 5637
rect 15766 5700 15800 5734
rect 15862 5701 15896 5735
rect 15422 5619 15456 5653
rect 15539 5619 15573 5653
rect 16030 5707 16064 5741
rect 16126 5707 16160 5741
rect 15952 5596 15986 5630
rect 8648 5287 8682 5321
rect 8744 5287 8778 5321
rect 8570 5176 8604 5210
rect 9370 4845 9404 4879
rect 9469 4853 9503 4887
rect 9541 4741 9575 4775
rect 9709 4869 9743 4903
rect 9809 4869 9843 4903
rect 9637 4741 9671 4775
rect 10238 4838 10272 4872
rect 10334 4839 10368 4873
rect 9894 4757 9928 4791
rect 10011 4757 10045 4791
rect 10502 4845 10536 4879
rect 10598 4845 10632 4879
rect 11240 4841 11274 4875
rect 10424 4734 10458 4768
rect 11339 4849 11373 4883
rect 11411 4737 11445 4771
rect 11579 4865 11613 4899
rect 11679 4865 11713 4899
rect 11507 4737 11541 4771
rect 12108 4834 12142 4868
rect 12204 4835 12238 4869
rect 11764 4753 11798 4787
rect 11881 4753 11915 4787
rect 12372 4841 12406 4875
rect 12468 4841 12502 4875
rect 13056 4837 13090 4871
rect 12294 4730 12328 4764
rect 13155 4845 13189 4879
rect 13227 4733 13261 4767
rect 13395 4861 13429 4895
rect 13495 4861 13529 4895
rect 13323 4733 13357 4767
rect 13924 4830 13958 4864
rect 14020 4831 14054 4865
rect 13580 4749 13614 4783
rect 13697 4749 13731 4783
rect 14188 4837 14222 4871
rect 14284 4837 14318 4871
rect 14926 4833 14960 4867
rect 14110 4726 14144 4760
rect 15025 4841 15059 4875
rect 15097 4729 15131 4763
rect 15265 4857 15299 4891
rect 15365 4857 15399 4891
rect 15193 4729 15227 4763
rect 15794 4826 15828 4860
rect 15890 4827 15924 4861
rect 15450 4745 15484 4779
rect 15567 4745 15601 4779
rect 16058 4833 16092 4867
rect 16154 4833 16188 4867
rect 15980 4722 16014 4756
rect 1930 2039 1964 2073
rect 2029 2047 2063 2081
rect 2101 1935 2135 1969
rect 2269 2063 2303 2097
rect 2369 2063 2403 2097
rect 2197 1935 2231 1969
rect 2798 2032 2832 2066
rect 2894 2033 2928 2067
rect 2454 1951 2488 1985
rect 2571 1951 2605 1985
rect 3062 2039 3096 2073
rect 3158 2039 3192 2073
rect 3800 2035 3834 2069
rect 2984 1928 3018 1962
rect 3899 2043 3933 2077
rect 3971 1931 4005 1965
rect 4139 2059 4173 2093
rect 4239 2059 4273 2093
rect 4067 1931 4101 1965
rect 4668 2028 4702 2062
rect 4764 2029 4798 2063
rect 4324 1947 4358 1981
rect 4441 1947 4475 1981
rect 4932 2035 4966 2069
rect 5028 2035 5062 2069
rect 5616 2031 5650 2065
rect 4854 1924 4888 1958
rect 5715 2039 5749 2073
rect 5787 1927 5821 1961
rect 5955 2055 5989 2089
rect 6055 2055 6089 2089
rect 5883 1927 5917 1961
rect 6484 2024 6518 2058
rect 6580 2025 6614 2059
rect 6140 1943 6174 1977
rect 6257 1943 6291 1977
rect 6748 2031 6782 2065
rect 6844 2031 6878 2065
rect 7486 2027 7520 2061
rect 6670 1920 6704 1954
rect 7585 2035 7619 2069
rect 7657 1923 7691 1957
rect 7825 2051 7859 2085
rect 7925 2051 7959 2085
rect 7753 1923 7787 1957
rect 8354 2020 8388 2054
rect 8450 2021 8484 2055
rect 8010 1939 8044 1973
rect 8127 1939 8161 1973
rect 8618 2027 8652 2061
rect 8714 2027 8748 2061
rect 9300 2025 9334 2059
rect 8540 1916 8574 1950
rect 9399 2033 9433 2067
rect 9471 1921 9505 1955
rect 9639 2049 9673 2083
rect 9739 2049 9773 2083
rect 9567 1921 9601 1955
rect 10168 2018 10202 2052
rect 10264 2019 10298 2053
rect 9824 1937 9858 1971
rect 9941 1937 9975 1971
rect 10432 2025 10466 2059
rect 10528 2025 10562 2059
rect 11170 2021 11204 2055
rect 10354 1914 10388 1948
rect 11269 2029 11303 2063
rect 11341 1917 11375 1951
rect 11509 2045 11543 2079
rect 11609 2045 11643 2079
rect 11437 1917 11471 1951
rect 12038 2014 12072 2048
rect 12134 2015 12168 2049
rect 11694 1933 11728 1967
rect 11811 1933 11845 1967
rect 12302 2021 12336 2055
rect 12398 2021 12432 2055
rect 12986 2017 13020 2051
rect 12224 1910 12258 1944
rect 13085 2025 13119 2059
rect 13157 1913 13191 1947
rect 13325 2041 13359 2075
rect 13425 2041 13459 2075
rect 13253 1913 13287 1947
rect 13854 2010 13888 2044
rect 13950 2011 13984 2045
rect 13510 1929 13544 1963
rect 13627 1929 13661 1963
rect 14118 2017 14152 2051
rect 14214 2017 14248 2051
rect 14856 2013 14890 2047
rect 14040 1906 14074 1940
rect 14955 2021 14989 2055
rect 15027 1909 15061 1943
rect 15195 2037 15229 2071
rect 15295 2037 15329 2071
rect 15123 1909 15157 1943
rect 15724 2006 15758 2040
rect 15820 2007 15854 2041
rect 15380 1925 15414 1959
rect 15497 1925 15531 1959
rect 15988 2013 16022 2047
rect 16084 2013 16118 2047
rect 15910 1902 15944 1936
<< locali >>
rect 9430 16553 9459 16587
rect 9493 16553 9551 16587
rect 9585 16553 9643 16587
rect 9677 16553 9735 16587
rect 9769 16553 9827 16587
rect 9861 16553 9919 16587
rect 9953 16553 10011 16587
rect 10045 16553 10074 16587
rect 9447 16511 9523 16519
rect 9447 16477 9473 16511
rect 9507 16477 9523 16511
rect 9447 16443 9523 16477
rect 9447 16409 9473 16443
rect 9507 16409 9523 16443
rect 9447 16383 9523 16409
rect 9641 16501 9675 16553
rect 9641 16433 9675 16467
rect 9641 16383 9675 16399
rect 9709 16501 9775 16519
rect 9709 16467 9725 16501
rect 9759 16467 9775 16501
rect 9709 16433 9775 16467
rect 9809 16501 9843 16553
rect 9809 16451 9843 16467
rect 9877 16501 9957 16519
rect 9877 16467 9913 16501
rect 9947 16467 9957 16501
rect 9709 16399 9725 16433
rect 9759 16417 9775 16433
rect 9877 16433 9957 16467
rect 9877 16417 9913 16433
rect 9759 16399 9913 16417
rect 9947 16399 9957 16433
rect 9709 16383 9957 16399
rect 9993 16503 10057 16519
rect 9993 16469 9997 16503
rect 10031 16469 10057 16503
rect 9993 16435 10057 16469
rect 9993 16401 9997 16435
rect 10031 16401 10057 16435
rect 9447 16191 9481 16383
rect 9993 16374 10057 16401
rect 9993 16367 10006 16374
rect 9515 16315 9776 16349
rect 9993 16333 9997 16367
rect 10040 16336 10057 16374
rect 10031 16333 10057 16336
rect 9515 16276 9564 16315
rect 9515 16275 9516 16276
rect 9550 16242 9564 16276
rect 9549 16241 9564 16242
rect 9598 16278 9708 16281
rect 9598 16275 9636 16278
rect 9598 16241 9632 16275
rect 9670 16244 9708 16278
rect 9666 16241 9708 16244
rect 9742 16275 9776 16315
rect 9931 16299 10057 16333
rect 9851 16275 9897 16291
rect 9742 16241 9767 16275
rect 9801 16241 9817 16275
rect 9851 16241 9863 16275
rect 9515 16225 9564 16241
rect 9851 16191 9897 16241
rect 9447 16157 9897 16191
rect 9557 16143 9591 16157
rect 9457 16087 9473 16121
rect 9507 16087 9523 16121
rect 9931 16123 9965 16299
rect 9557 16093 9591 16109
rect 9457 16043 9523 16087
rect 9625 16087 9641 16121
rect 9675 16087 9691 16121
rect 9774 16089 9809 16123
rect 9843 16089 9909 16123
rect 9943 16089 9965 16123
rect 9999 16194 10057 16210
rect 10033 16160 10057 16194
rect 9999 16126 10057 16160
rect 10033 16092 10057 16126
rect 9625 16043 9691 16087
rect 9999 16043 10057 16092
rect 9430 16009 9459 16043
rect 9493 16009 9551 16043
rect 9585 16009 9643 16043
rect 9677 16009 9735 16043
rect 9769 16009 9827 16043
rect 9861 16009 9919 16043
rect 9953 16009 10011 16043
rect 10045 16009 10074 16043
rect 9528 15809 9557 15843
rect 9591 15809 9649 15843
rect 9683 15809 9741 15843
rect 9775 15809 9833 15843
rect 9867 15809 9925 15843
rect 9959 15809 9988 15843
rect 9585 15725 9641 15809
rect 9775 15767 9841 15809
rect 9585 15691 9599 15725
rect 9633 15691 9641 15725
rect 9585 15675 9641 15691
rect 9675 15725 9735 15741
rect 9675 15691 9683 15725
rect 9717 15691 9735 15725
rect 9675 15631 9735 15691
rect 9775 15733 9791 15767
rect 9825 15733 9841 15767
rect 9775 15699 9841 15733
rect 9775 15665 9791 15699
rect 9825 15665 9841 15699
rect 9879 15767 9971 15775
rect 9879 15733 9895 15767
rect 9929 15733 9971 15767
rect 9879 15699 9971 15733
rect 11570 15699 11599 15733
rect 11633 15699 11691 15733
rect 11725 15699 11783 15733
rect 11817 15699 11875 15733
rect 11909 15699 11967 15733
rect 12001 15699 12059 15733
rect 12093 15699 12151 15733
rect 12185 15699 12214 15733
rect 9879 15665 9895 15699
rect 9929 15665 9971 15699
rect 9548 15554 9601 15619
rect 9675 15597 9863 15631
rect 9548 15514 9550 15554
rect 9592 15547 9601 15554
rect 9829 15547 9863 15597
rect 9592 15531 9683 15547
rect 9592 15514 9602 15531
rect 9548 15497 9602 15514
rect 9636 15497 9683 15531
rect 9727 15544 9795 15547
rect 9727 15504 9740 15544
rect 9782 15504 9795 15544
rect 9727 15497 9743 15504
rect 9777 15497 9795 15504
rect 9829 15531 9887 15547
rect 9829 15497 9851 15531
rect 9885 15497 9887 15531
rect 9829 15481 9887 15497
rect 9829 15463 9863 15481
rect 9585 15425 9863 15463
rect 9921 15474 9971 15665
rect 11588 15657 11655 15699
rect 11588 15623 11605 15657
rect 11639 15623 11655 15657
rect 11689 15649 11739 15665
rect 11689 15615 11697 15649
rect 11731 15615 11739 15649
rect 9921 15440 9932 15474
rect 9968 15440 9971 15474
rect 9585 15403 9651 15425
rect 9585 15369 9599 15403
rect 9633 15369 9651 15403
rect 9921 15391 9971 15440
rect 9585 15353 9651 15369
rect 9775 15375 9825 15391
rect 9775 15341 9791 15375
rect 9775 15299 9825 15341
rect 9859 15375 9971 15391
rect 9859 15341 9875 15375
rect 9909 15341 9971 15375
rect 9859 15333 9971 15341
rect 11587 15421 11635 15587
rect 11689 15505 11739 15615
rect 11783 15657 11849 15699
rect 11783 15623 11799 15657
rect 11833 15623 11849 15657
rect 11783 15555 11849 15623
rect 11886 15649 11936 15665
rect 11886 15615 11894 15649
rect 11928 15615 11936 15649
rect 11886 15505 11936 15615
rect 12029 15657 12095 15699
rect 12029 15623 12045 15657
rect 12079 15623 12095 15657
rect 12029 15589 12095 15623
rect 12129 15657 12197 15665
rect 12129 15623 12145 15657
rect 12179 15623 12197 15657
rect 12129 15613 12197 15623
rect 12029 15555 12045 15589
rect 12079 15555 12095 15589
rect 12029 15539 12095 15555
rect 12145 15589 12197 15613
rect 12179 15555 12197 15589
rect 12145 15521 12197 15555
rect 11587 15387 11601 15421
rect 11587 15384 11635 15387
rect 11587 15348 11594 15384
rect 11630 15348 11635 15384
rect 11587 15325 11635 15348
rect 11669 15471 12107 15505
rect 9528 15265 9557 15299
rect 9591 15265 9649 15299
rect 9683 15265 9741 15299
rect 9775 15265 9833 15299
rect 9867 15265 9925 15299
rect 9959 15265 9988 15299
rect 11669 15289 11703 15471
rect 12044 15437 12107 15471
rect 12179 15487 12197 15521
rect 11604 15273 11703 15289
rect 11604 15239 11605 15273
rect 11639 15239 11703 15273
rect 11747 15421 11817 15437
rect 11781 15418 11817 15421
rect 11747 15382 11766 15387
rect 11800 15382 11817 15418
rect 11747 15244 11817 15382
rect 11853 15421 11913 15437
rect 11887 15387 11913 15421
rect 11853 15294 11913 15387
rect 11853 15260 11864 15294
rect 11898 15260 11913 15294
rect 11853 15243 11913 15260
rect 11949 15421 12005 15437
rect 11983 15387 12005 15421
rect 12044 15421 12110 15437
rect 12044 15387 12060 15421
rect 12094 15387 12110 15421
rect 12145 15416 12197 15487
rect 11949 15364 12005 15387
rect 11949 15328 11960 15364
rect 11994 15328 12005 15364
rect 12145 15382 12152 15416
rect 12186 15382 12197 15416
rect 11949 15243 12005 15328
rect 12041 15333 12095 15349
rect 12145 15333 12197 15382
rect 12041 15299 12046 15333
rect 12080 15299 12095 15333
rect 12041 15265 12095 15299
rect 10712 15199 10741 15233
rect 10775 15199 10833 15233
rect 10867 15199 10925 15233
rect 10959 15199 11017 15233
rect 11051 15199 11109 15233
rect 11143 15199 11172 15233
rect 11604 15223 11703 15239
rect 12041 15231 12046 15265
rect 12080 15231 12095 15265
rect 12129 15299 12145 15333
rect 12179 15299 12197 15333
rect 12129 15265 12197 15299
rect 12129 15231 12145 15265
rect 12179 15231 12197 15265
rect 10769 15115 10825 15199
rect 10959 15157 11025 15199
rect 12041 15189 12095 15231
rect 10769 15081 10783 15115
rect 10817 15081 10825 15115
rect 10769 15065 10825 15081
rect 10859 15115 10919 15131
rect 10859 15081 10867 15115
rect 10901 15081 10919 15115
rect 9440 14989 9469 15023
rect 9503 14989 9561 15023
rect 9595 14989 9653 15023
rect 9687 14989 9745 15023
rect 9779 14989 9837 15023
rect 9871 14989 9929 15023
rect 9963 14989 10021 15023
rect 10055 14989 10084 15023
rect 10859 15021 10919 15081
rect 10959 15123 10975 15157
rect 11009 15123 11025 15157
rect 10959 15089 11025 15123
rect 10959 15055 10975 15089
rect 11009 15055 11025 15089
rect 11063 15157 11155 15165
rect 11063 15123 11079 15157
rect 11113 15132 11155 15157
rect 11570 15155 11599 15189
rect 11633 15155 11691 15189
rect 11725 15155 11783 15189
rect 11817 15155 11875 15189
rect 11909 15155 11967 15189
rect 12001 15155 12059 15189
rect 12093 15155 12151 15189
rect 12185 15155 12214 15189
rect 11063 15096 11106 15123
rect 11146 15096 11155 15132
rect 11063 15089 11155 15096
rect 11063 15055 11079 15089
rect 11113 15055 11155 15089
rect 9457 14947 9533 14955
rect 9457 14913 9483 14947
rect 9517 14913 9533 14947
rect 9457 14879 9533 14913
rect 9457 14845 9483 14879
rect 9517 14845 9533 14879
rect 9457 14819 9533 14845
rect 9651 14937 9685 14989
rect 9651 14869 9685 14903
rect 9651 14819 9685 14835
rect 9719 14937 9785 14955
rect 9719 14903 9735 14937
rect 9769 14903 9785 14937
rect 9719 14869 9785 14903
rect 9819 14937 9853 14989
rect 9819 14887 9853 14903
rect 9887 14937 9967 14955
rect 9887 14903 9923 14937
rect 9957 14903 9967 14937
rect 9719 14835 9735 14869
rect 9769 14853 9785 14869
rect 9887 14869 9967 14903
rect 9887 14853 9923 14869
rect 9769 14835 9923 14853
rect 9957 14835 9967 14869
rect 9719 14819 9967 14835
rect 10003 14939 10067 14955
rect 10003 14905 10007 14939
rect 10041 14914 10067 14939
rect 10003 14880 10018 14905
rect 10052 14880 10067 14914
rect 10732 14937 10785 15009
rect 10859 14987 11047 15021
rect 11013 14937 11047 14987
rect 10732 14922 10867 14937
rect 10732 14887 10786 14922
rect 10820 14887 10867 14922
rect 10911 14922 10979 14937
rect 10911 14888 10926 14922
rect 10962 14888 10979 14922
rect 10911 14887 10927 14888
rect 10961 14887 10979 14888
rect 11013 14921 11071 14937
rect 11013 14887 11035 14921
rect 11069 14887 11071 14921
rect 10003 14871 10067 14880
rect 10003 14837 10007 14871
rect 10041 14837 10067 14871
rect 11013 14871 11071 14887
rect 11013 14853 11047 14871
rect 9457 14627 9491 14819
rect 10003 14803 10067 14837
rect 9525 14751 9786 14785
rect 10003 14769 10007 14803
rect 10041 14769 10067 14803
rect 9525 14712 9574 14751
rect 9525 14711 9526 14712
rect 9560 14678 9574 14712
rect 9559 14677 9574 14678
rect 9608 14714 9718 14717
rect 9608 14711 9646 14714
rect 9608 14677 9642 14711
rect 9680 14680 9718 14714
rect 9676 14677 9718 14680
rect 9752 14711 9786 14751
rect 9941 14735 10067 14769
rect 10769 14815 11047 14853
rect 10769 14793 10835 14815
rect 10769 14759 10783 14793
rect 10817 14759 10835 14793
rect 11105 14781 11155 15055
rect 10769 14743 10835 14759
rect 10959 14765 11009 14781
rect 9861 14711 9907 14727
rect 9752 14677 9777 14711
rect 9811 14677 9827 14711
rect 9861 14677 9873 14711
rect 9525 14661 9574 14677
rect 9861 14627 9907 14677
rect 9457 14593 9907 14627
rect 9567 14579 9601 14593
rect 9467 14523 9483 14557
rect 9517 14523 9533 14557
rect 9941 14559 9975 14735
rect 10959 14731 10975 14765
rect 10959 14689 11009 14731
rect 11043 14765 11155 14781
rect 11043 14731 11059 14765
rect 11093 14731 11155 14765
rect 11043 14723 11155 14731
rect 10712 14655 10741 14689
rect 10775 14655 10833 14689
rect 10867 14655 10925 14689
rect 10959 14655 11017 14689
rect 11051 14655 11109 14689
rect 11143 14655 11172 14689
rect 9567 14529 9601 14545
rect 9467 14479 9533 14523
rect 9635 14523 9651 14557
rect 9685 14523 9701 14557
rect 9784 14525 9819 14559
rect 9853 14525 9919 14559
rect 9953 14525 9975 14559
rect 10009 14630 10067 14646
rect 10043 14596 10067 14630
rect 10009 14562 10067 14596
rect 10043 14528 10067 14562
rect 9635 14479 9701 14523
rect 10009 14479 10067 14528
rect 9440 14445 9469 14479
rect 9503 14445 9561 14479
rect 9595 14445 9653 14479
rect 9687 14445 9745 14479
rect 9779 14445 9837 14479
rect 9871 14445 9929 14479
rect 9963 14445 10021 14479
rect 10055 14445 10084 14479
rect 9538 14245 9567 14279
rect 9601 14245 9659 14279
rect 9693 14245 9751 14279
rect 9785 14245 9843 14279
rect 9877 14245 9935 14279
rect 9969 14245 9998 14279
rect 9595 14161 9651 14245
rect 9785 14203 9851 14245
rect 10786 14233 10815 14267
rect 10849 14233 10907 14267
rect 10941 14233 10999 14267
rect 11033 14233 11091 14267
rect 11125 14233 11183 14267
rect 11217 14233 11275 14267
rect 11309 14233 11367 14267
rect 11401 14233 11430 14267
rect 9595 14127 9609 14161
rect 9643 14127 9651 14161
rect 9595 14111 9651 14127
rect 9685 14161 9745 14177
rect 9685 14127 9693 14161
rect 9727 14127 9745 14161
rect 9685 14067 9745 14127
rect 9785 14169 9801 14203
rect 9835 14169 9851 14203
rect 9785 14135 9851 14169
rect 9785 14101 9801 14135
rect 9835 14101 9851 14135
rect 9889 14203 9981 14211
rect 9889 14169 9905 14203
rect 9939 14169 9981 14203
rect 9889 14135 9981 14169
rect 10804 14191 10871 14233
rect 10804 14157 10821 14191
rect 10855 14157 10871 14191
rect 10905 14183 10955 14199
rect 9889 14101 9905 14135
rect 9939 14101 9981 14135
rect 10905 14149 10913 14183
rect 10947 14149 10955 14183
rect 9558 13990 9611 14055
rect 9685 14033 9873 14067
rect 9558 13950 9560 13990
rect 9602 13983 9611 13990
rect 9839 13983 9873 14033
rect 9602 13967 9693 13983
rect 9602 13950 9612 13967
rect 9558 13933 9612 13950
rect 9646 13933 9693 13967
rect 9737 13980 9805 13983
rect 9737 13940 9750 13980
rect 9792 13940 9805 13980
rect 9737 13933 9753 13940
rect 9787 13933 9805 13940
rect 9839 13967 9897 13983
rect 9839 13933 9861 13967
rect 9895 13933 9897 13967
rect 9839 13917 9897 13933
rect 9839 13899 9873 13917
rect 9595 13861 9873 13899
rect 9931 13868 9981 14101
rect 9595 13839 9661 13861
rect 9595 13805 9609 13839
rect 9643 13805 9661 13839
rect 9931 13834 9940 13868
rect 9976 13834 9981 13868
rect 10803 13960 10851 14121
rect 10905 14039 10955 14149
rect 10999 14191 11065 14233
rect 10999 14157 11015 14191
rect 11049 14157 11065 14191
rect 10999 14089 11065 14157
rect 11102 14183 11152 14199
rect 11102 14149 11110 14183
rect 11144 14149 11152 14183
rect 11102 14039 11152 14149
rect 11245 14191 11311 14233
rect 12604 14217 12633 14251
rect 12667 14217 12725 14251
rect 12759 14217 12817 14251
rect 12851 14217 12909 14251
rect 12943 14217 13001 14251
rect 13035 14217 13093 14251
rect 13127 14217 13156 14251
rect 11245 14157 11261 14191
rect 11295 14157 11311 14191
rect 11245 14123 11311 14157
rect 11345 14191 11413 14199
rect 11345 14157 11361 14191
rect 11395 14157 11413 14191
rect 12987 14175 13043 14217
rect 11345 14147 11413 14157
rect 11245 14089 11261 14123
rect 11295 14089 11311 14123
rect 11245 14073 11311 14089
rect 11361 14123 11413 14147
rect 11395 14089 11413 14123
rect 12622 14163 12953 14173
rect 12622 14150 12861 14163
rect 12622 14116 12778 14150
rect 12814 14129 12861 14150
rect 12895 14129 12953 14163
rect 12814 14116 12953 14129
rect 12622 14115 12953 14116
rect 12987 14141 13000 14175
rect 13034 14141 13043 14175
rect 11361 14055 11413 14089
rect 12987 14107 13043 14141
rect 10803 13926 10812 13960
rect 10846 13955 10851 13960
rect 10803 13921 10817 13926
rect 10803 13859 10851 13921
rect 10885 14005 11323 14039
rect 9931 13827 9981 13834
rect 9595 13789 9661 13805
rect 9785 13811 9835 13827
rect 9785 13777 9801 13811
rect 9785 13735 9835 13777
rect 9869 13811 9981 13827
rect 10885 13823 10919 14005
rect 11260 13971 11323 14005
rect 11395 14021 11413 14055
rect 9869 13777 9885 13811
rect 9919 13777 9981 13811
rect 9869 13769 9981 13777
rect 10820 13807 10919 13823
rect 10820 13773 10821 13807
rect 10855 13773 10919 13807
rect 10963 13955 11033 13971
rect 10997 13921 11033 13955
rect 10963 13864 11033 13921
rect 10963 13830 10982 13864
rect 11016 13830 11033 13864
rect 10963 13778 11033 13830
rect 11069 13955 11129 13971
rect 11103 13921 11129 13955
rect 11069 13904 11129 13921
rect 11069 13870 11080 13904
rect 11114 13870 11129 13904
rect 11069 13777 11129 13870
rect 11165 13955 11221 13971
rect 11199 13954 11221 13955
rect 11165 13916 11174 13921
rect 11210 13916 11221 13954
rect 11260 13955 11326 13971
rect 11260 13921 11276 13955
rect 11310 13921 11326 13955
rect 11165 13777 11221 13916
rect 11257 13867 11311 13883
rect 11361 13867 11413 14021
rect 12622 14047 12940 14081
rect 12987 14073 13000 14107
rect 13034 14073 13043 14107
rect 12987 14057 13043 14073
rect 13085 14144 13139 14183
rect 13119 14110 13139 14144
rect 13085 14076 13139 14110
rect 12622 14044 12686 14047
rect 12622 14010 12639 14044
rect 12673 14010 12686 14044
rect 12906 14023 12940 14047
rect 13119 14056 13139 14076
rect 12622 13989 12686 14010
rect 12622 13939 12692 13955
rect 12622 13932 12639 13939
rect 12673 13932 12692 13939
rect 12622 13898 12636 13932
rect 12676 13898 12692 13932
rect 11257 13833 11262 13867
rect 11296 13833 11311 13867
rect 11257 13799 11311 13833
rect 10820 13757 10919 13773
rect 11257 13765 11262 13799
rect 11296 13765 11311 13799
rect 11345 13836 11361 13867
rect 11345 13798 11356 13836
rect 11395 13833 11413 13867
rect 11756 13859 11785 13893
rect 11819 13859 11877 13893
rect 11911 13859 11969 13893
rect 12003 13859 12061 13893
rect 12095 13859 12153 13893
rect 12187 13859 12216 13893
rect 11394 13799 11413 13833
rect 11345 13765 11361 13798
rect 11395 13765 11413 13799
rect 11985 13801 12051 13859
rect 12622 13841 12692 13898
rect 12726 13944 12868 14013
rect 12906 13989 13051 14023
rect 13085 14016 13092 14042
rect 13134 14016 13139 14056
rect 13085 13989 13139 14016
rect 13017 13955 13051 13989
rect 12726 13902 12762 13944
rect 12812 13902 12868 13944
rect 12726 13889 12868 13902
rect 12902 13940 12983 13955
rect 12902 13904 12934 13940
rect 12972 13939 12983 13940
rect 12975 13905 12983 13939
rect 12972 13904 12983 13905
rect 12902 13889 12983 13904
rect 13017 13939 13071 13955
rect 13017 13905 13037 13939
rect 13017 13889 13071 13905
rect 13017 13855 13051 13889
rect 11985 13767 12001 13801
rect 12035 13767 12051 13801
rect 9538 13701 9567 13735
rect 9601 13701 9659 13735
rect 9693 13701 9751 13735
rect 9785 13701 9843 13735
rect 9877 13701 9935 13735
rect 9969 13701 9998 13735
rect 11257 13723 11311 13765
rect 11985 13733 12051 13767
rect 10786 13689 10815 13723
rect 10849 13689 10907 13723
rect 10941 13689 10999 13723
rect 11033 13689 11091 13723
rect 11125 13689 11183 13723
rect 11217 13689 11275 13723
rect 11309 13689 11367 13723
rect 11401 13689 11430 13723
rect 11810 13681 11888 13700
rect 11985 13699 12001 13733
rect 12035 13699 12051 13733
rect 12085 13817 12192 13825
rect 12085 13783 12101 13817
rect 12135 13783 12192 13817
rect 12729 13821 13051 13855
rect 13105 13842 13139 13989
rect 13085 13825 13139 13842
rect 12085 13749 12192 13783
rect 12085 13715 12101 13749
rect 12135 13748 12192 13749
rect 12085 13714 12124 13715
rect 12158 13714 12192 13748
rect 12085 13701 12192 13714
rect 12623 13773 12639 13807
rect 12673 13773 12689 13807
rect 12623 13707 12689 13773
rect 12729 13801 12763 13821
rect 12903 13801 12937 13821
rect 12729 13751 12763 13767
rect 12803 13753 12819 13787
rect 12853 13753 12869 13787
rect 12803 13707 12869 13753
rect 13119 13791 13139 13825
rect 12903 13751 12937 13767
rect 12971 13753 12997 13787
rect 13031 13753 13047 13787
rect 13085 13773 13139 13791
rect 12971 13707 13047 13753
rect 11810 13647 11832 13681
rect 11866 13665 11888 13681
rect 11866 13647 12095 13665
rect 11810 13631 12095 13647
rect 11785 13581 11856 13597
rect 11785 13547 11822 13581
rect 11785 13538 11856 13547
rect 11785 13504 11796 13538
rect 11830 13504 11856 13538
rect 11785 13485 11856 13504
rect 11890 13451 11924 13631
rect 11958 13588 12011 13597
rect 11958 13581 11974 13588
rect 12008 13554 12011 13588
rect 11992 13547 12011 13554
rect 11958 13485 12011 13547
rect 12061 13581 12095 13631
rect 12061 13531 12095 13547
rect 12129 13497 12192 13701
rect 12604 13673 12633 13707
rect 12667 13673 12725 13707
rect 12759 13673 12817 13707
rect 12851 13673 12909 13707
rect 12943 13673 13001 13707
rect 13035 13673 13093 13707
rect 13127 13673 13156 13707
rect 12069 13495 12192 13497
rect 12069 13461 12085 13495
rect 12119 13461 12192 13495
rect 11806 13435 11854 13451
rect 10910 13391 10939 13425
rect 10973 13391 11031 13425
rect 11065 13391 11123 13425
rect 11157 13391 11215 13425
rect 11249 13391 11307 13425
rect 11341 13391 11370 13425
rect 11806 13401 11820 13435
rect 9432 13321 9461 13355
rect 9495 13321 9553 13355
rect 9587 13321 9645 13355
rect 9679 13321 9737 13355
rect 9771 13321 9829 13355
rect 9863 13321 9921 13355
rect 9955 13321 10013 13355
rect 10047 13321 10076 13355
rect 9449 13279 9525 13287
rect 9449 13245 9475 13279
rect 9509 13245 9525 13279
rect 9449 13211 9525 13245
rect 9449 13177 9475 13211
rect 9509 13177 9525 13211
rect 9449 13151 9525 13177
rect 9643 13269 9677 13321
rect 9643 13201 9677 13235
rect 9643 13151 9677 13167
rect 9711 13269 9777 13287
rect 9711 13235 9727 13269
rect 9761 13235 9777 13269
rect 9711 13201 9777 13235
rect 9811 13269 9845 13321
rect 9811 13219 9845 13235
rect 9879 13269 9959 13287
rect 9879 13235 9915 13269
rect 9949 13235 9959 13269
rect 9711 13167 9727 13201
rect 9761 13185 9777 13201
rect 9879 13201 9959 13235
rect 9879 13185 9915 13201
rect 9761 13167 9915 13185
rect 9949 13167 9959 13201
rect 9711 13151 9959 13167
rect 9995 13271 10059 13287
rect 9995 13237 9999 13271
rect 10033 13237 10059 13271
rect 10927 13280 11048 13391
rect 11083 13340 11179 13357
rect 11117 13318 11179 13340
rect 11083 13289 11108 13306
rect 11144 13289 11179 13318
rect 11213 13349 11264 13391
rect 11213 13315 11217 13349
rect 11251 13315 11264 13349
rect 11213 13282 11264 13315
rect 11298 13335 11353 13357
rect 11806 13349 11854 13401
rect 11890 13435 11946 13451
rect 11890 13401 11904 13435
rect 11938 13401 11946 13435
rect 11890 13385 11946 13401
rect 11992 13435 12035 13451
rect 11992 13401 12000 13435
rect 12034 13401 12035 13435
rect 11992 13349 12035 13401
rect 12069 13427 12192 13461
rect 12069 13393 12085 13427
rect 12119 13393 12192 13427
rect 12069 13383 12192 13393
rect 11298 13301 11301 13335
rect 11335 13301 11353 13335
rect 11756 13315 11785 13349
rect 11819 13315 11877 13349
rect 11911 13315 11969 13349
rect 12003 13315 12061 13349
rect 12095 13315 12153 13349
rect 12187 13315 12216 13349
rect 10927 13260 11050 13280
rect 9995 13204 10059 13237
rect 11013 13255 11050 13260
rect 11298 13267 11353 13301
rect 11013 13240 11079 13255
rect 9995 13203 10010 13204
rect 9995 13169 9999 13203
rect 10044 13170 10059 13204
rect 10033 13169 10059 13170
rect 9449 12959 9483 13151
rect 9995 13135 10059 13169
rect 9517 13083 9778 13117
rect 9995 13101 9999 13135
rect 10033 13101 10059 13135
rect 10927 13210 10979 13226
rect 10927 13176 10945 13210
rect 11013 13206 11029 13240
rect 11063 13206 11079 13240
rect 11113 13221 11264 13241
rect 11113 13191 11122 13221
rect 11110 13187 11122 13191
rect 11156 13187 11264 13221
rect 11298 13233 11301 13267
rect 11335 13262 11353 13267
rect 11298 13224 11304 13233
rect 11342 13224 11353 13262
rect 11298 13217 11353 13224
rect 11110 13184 11264 13187
rect 11107 13182 11264 13184
rect 11106 13179 11285 13182
rect 11102 13176 11285 13179
rect 10927 13136 10979 13176
rect 11098 13174 11285 13176
rect 11093 13172 11285 13174
rect 11079 13166 11285 13172
rect 11075 13160 11285 13166
rect 11071 13154 11285 13160
rect 11065 13149 11285 13154
rect 11058 13142 11285 13149
rect 11052 13141 11285 13142
rect 11052 13140 11130 13141
rect 11052 13138 11125 13140
rect 11052 13137 11122 13138
rect 11052 13136 11119 13137
rect 10927 13135 11119 13136
rect 10927 13133 11117 13135
rect 10927 13132 11115 13133
rect 10927 13130 11113 13132
rect 10927 13128 11112 13130
rect 10927 13127 11111 13128
rect 10927 13124 11109 13127
rect 10927 13121 11108 13124
rect 10927 13116 11106 13121
rect 10927 13102 11105 13116
rect 11239 13113 11285 13141
rect 9517 13044 9566 13083
rect 9517 13043 9518 13044
rect 9552 13010 9566 13044
rect 9551 13009 9566 13010
rect 9600 13046 9710 13049
rect 9600 13043 9638 13046
rect 9600 13009 9634 13043
rect 9672 13012 9710 13046
rect 9668 13009 9710 13012
rect 9744 13043 9778 13083
rect 9933 13067 10059 13101
rect 10927 13067 11037 13068
rect 9853 13043 9899 13059
rect 9744 13009 9769 13043
rect 9803 13009 9819 13043
rect 9853 13009 9865 13043
rect 9517 12993 9566 13009
rect 9853 12959 9899 13009
rect 9449 12925 9899 12959
rect 9559 12911 9593 12925
rect 9459 12855 9475 12889
rect 9509 12855 9525 12889
rect 9933 12891 9967 13067
rect 10927 13033 10945 13067
rect 10979 13044 11037 13067
rect 10927 13010 10956 13033
rect 10990 13010 11037 13044
rect 10927 12991 11037 13010
rect 9559 12861 9593 12877
rect 9459 12811 9525 12855
rect 9627 12855 9643 12889
rect 9677 12855 9693 12889
rect 9776 12857 9811 12891
rect 9845 12857 9911 12891
rect 9945 12857 9967 12891
rect 10001 12962 10059 12978
rect 10035 12928 10059 12962
rect 11071 12957 11105 13102
rect 10001 12894 10059 12928
rect 10927 12923 10945 12957
rect 10979 12923 11105 12957
rect 11139 13073 11155 13107
rect 11189 13073 11205 13107
rect 11139 13050 11205 13073
rect 11239 13079 11251 13113
rect 11239 13062 11285 13079
rect 11139 13016 11158 13050
rect 11194 13022 11205 13050
rect 11139 12925 11183 13016
rect 11319 13011 11353 13217
rect 11217 12973 11267 12989
rect 11251 12939 11267 12973
rect 10035 12860 10059 12894
rect 11217 12881 11267 12939
rect 11301 12983 11353 13011
rect 11335 12949 11353 12983
rect 11301 12915 11353 12949
rect 9627 12811 9693 12855
rect 10001 12811 10059 12860
rect 10910 12847 10939 12881
rect 10973 12847 11031 12881
rect 11065 12847 11123 12881
rect 11157 12847 11215 12881
rect 11249 12847 11307 12881
rect 11341 12847 11370 12881
rect 9432 12777 9461 12811
rect 9495 12777 9553 12811
rect 9587 12777 9645 12811
rect 9679 12777 9737 12811
rect 9771 12777 9829 12811
rect 9863 12777 9921 12811
rect 9955 12777 10013 12811
rect 10047 12777 10076 12811
rect 9530 12577 9559 12611
rect 9593 12577 9651 12611
rect 9685 12577 9743 12611
rect 9777 12577 9835 12611
rect 9869 12577 9927 12611
rect 9961 12577 9990 12611
rect 9587 12493 9643 12577
rect 9777 12535 9843 12577
rect 9587 12459 9601 12493
rect 9635 12459 9643 12493
rect 9587 12443 9643 12459
rect 9677 12493 9737 12509
rect 9677 12459 9685 12493
rect 9719 12459 9737 12493
rect 9677 12399 9737 12459
rect 9777 12501 9793 12535
rect 9827 12501 9843 12535
rect 9777 12467 9843 12501
rect 9777 12433 9793 12467
rect 9827 12433 9843 12467
rect 9881 12535 9973 12543
rect 9881 12501 9897 12535
rect 9931 12501 9973 12535
rect 9881 12467 9973 12501
rect 9881 12433 9897 12467
rect 9931 12433 9973 12467
rect 9550 12322 9603 12387
rect 9677 12365 9865 12399
rect 9550 12282 9552 12322
rect 9594 12315 9603 12322
rect 9831 12315 9865 12365
rect 9923 12354 9973 12433
rect 10906 12371 10935 12405
rect 10969 12371 11027 12405
rect 11061 12371 11119 12405
rect 11153 12371 11211 12405
rect 11245 12371 11303 12405
rect 11337 12371 11366 12405
rect 9923 12320 9932 12354
rect 9968 12320 9973 12354
rect 9594 12299 9685 12315
rect 9594 12282 9604 12299
rect 9550 12265 9604 12282
rect 9638 12265 9685 12299
rect 9729 12312 9797 12315
rect 9729 12272 9742 12312
rect 9784 12272 9797 12312
rect 9729 12265 9745 12272
rect 9779 12265 9797 12272
rect 9831 12299 9889 12315
rect 9831 12265 9853 12299
rect 9887 12265 9889 12299
rect 9831 12249 9889 12265
rect 9831 12231 9865 12249
rect 9587 12193 9865 12231
rect 9587 12171 9653 12193
rect 9587 12137 9601 12171
rect 9635 12137 9653 12171
rect 9923 12159 9973 12320
rect 10963 12287 11019 12371
rect 11153 12329 11219 12371
rect 10963 12253 10977 12287
rect 11011 12253 11019 12287
rect 10963 12237 11019 12253
rect 11053 12287 11113 12303
rect 11053 12253 11061 12287
rect 11095 12253 11113 12287
rect 11053 12193 11113 12253
rect 11153 12295 11169 12329
rect 11203 12295 11219 12329
rect 11153 12261 11219 12295
rect 11153 12227 11169 12261
rect 11203 12227 11219 12261
rect 11257 12329 11349 12337
rect 11257 12295 11273 12329
rect 11307 12295 11349 12329
rect 11257 12261 11349 12295
rect 11257 12227 11273 12261
rect 11307 12227 11349 12261
rect 9587 12121 9653 12137
rect 9777 12143 9827 12159
rect 9777 12109 9793 12143
rect 9777 12067 9827 12109
rect 9861 12143 9973 12159
rect 9861 12109 9877 12143
rect 9911 12109 9973 12143
rect 9861 12101 9973 12109
rect 10926 12109 10979 12181
rect 11053 12159 11241 12193
rect 11207 12109 11241 12159
rect 11299 12180 11349 12227
rect 11299 12146 11308 12180
rect 11342 12146 11349 12180
rect 10926 12096 11061 12109
rect 9530 12033 9559 12067
rect 9593 12033 9651 12067
rect 9685 12033 9743 12067
rect 9777 12033 9835 12067
rect 9869 12033 9927 12067
rect 9961 12033 9990 12067
rect 10926 12059 10980 12096
rect 11016 12062 11061 12096
rect 11014 12059 11061 12062
rect 11105 12094 11173 12109
rect 11105 12060 11120 12094
rect 11156 12060 11173 12094
rect 11105 12059 11121 12060
rect 11155 12059 11173 12060
rect 11207 12093 11265 12109
rect 11207 12059 11229 12093
rect 11263 12059 11265 12093
rect 11207 12043 11265 12059
rect 11207 12025 11241 12043
rect 10963 11987 11241 12025
rect 10963 11965 11029 11987
rect 10963 11931 10977 11965
rect 11011 11931 11029 11965
rect 11299 11953 11349 12146
rect 10963 11915 11029 11931
rect 11153 11937 11203 11953
rect 11153 11903 11169 11937
rect 11153 11861 11203 11903
rect 11237 11937 11349 11953
rect 11237 11903 11253 11937
rect 11287 11903 11349 11937
rect 11237 11895 11349 11903
rect 10906 11827 10935 11861
rect 10969 11827 11027 11861
rect 11061 11827 11119 11861
rect 11153 11827 11211 11861
rect 11245 11827 11303 11861
rect 11337 11827 11366 11861
rect 9442 11757 9471 11791
rect 9505 11757 9563 11791
rect 9597 11757 9655 11791
rect 9689 11757 9747 11791
rect 9781 11757 9839 11791
rect 9873 11757 9931 11791
rect 9965 11757 10023 11791
rect 10057 11757 10086 11791
rect 9459 11715 9535 11723
rect 9459 11681 9485 11715
rect 9519 11681 9535 11715
rect 9459 11647 9535 11681
rect 9459 11613 9485 11647
rect 9519 11613 9535 11647
rect 9459 11587 9535 11613
rect 9653 11705 9687 11757
rect 9653 11637 9687 11671
rect 9653 11587 9687 11603
rect 9721 11705 9787 11723
rect 9721 11671 9737 11705
rect 9771 11671 9787 11705
rect 9721 11637 9787 11671
rect 9821 11705 9855 11757
rect 9821 11655 9855 11671
rect 9889 11705 9969 11723
rect 9889 11671 9925 11705
rect 9959 11671 9969 11705
rect 9721 11603 9737 11637
rect 9771 11621 9787 11637
rect 9889 11637 9969 11671
rect 9889 11621 9925 11637
rect 9771 11603 9925 11621
rect 9959 11603 9969 11637
rect 9721 11587 9969 11603
rect 10005 11707 10069 11723
rect 10005 11673 10009 11707
rect 10043 11673 10069 11707
rect 10005 11640 10069 11673
rect 10005 11639 10010 11640
rect 10005 11605 10009 11639
rect 10046 11606 10069 11640
rect 10043 11605 10069 11606
rect 9459 11395 9493 11587
rect 10005 11571 10069 11605
rect 9527 11519 9788 11553
rect 10005 11537 10009 11571
rect 10043 11537 10069 11571
rect 9527 11480 9576 11519
rect 9527 11479 9528 11480
rect 9562 11446 9576 11480
rect 9561 11445 9576 11446
rect 9610 11482 9720 11485
rect 9610 11479 9648 11482
rect 9610 11445 9644 11479
rect 9682 11448 9720 11482
rect 9678 11445 9720 11448
rect 9754 11479 9788 11519
rect 9943 11503 10069 11537
rect 9863 11479 9909 11495
rect 9754 11445 9779 11479
rect 9813 11445 9829 11479
rect 9863 11445 9875 11479
rect 9527 11429 9576 11445
rect 9863 11395 9909 11445
rect 9459 11361 9909 11395
rect 9569 11347 9603 11361
rect 9469 11291 9485 11325
rect 9519 11291 9535 11325
rect 9943 11327 9977 11503
rect 9569 11297 9603 11313
rect 9469 11247 9535 11291
rect 9637 11291 9653 11325
rect 9687 11291 9703 11325
rect 9786 11293 9821 11327
rect 9855 11293 9921 11327
rect 9955 11293 9977 11327
rect 10011 11398 10069 11414
rect 10045 11364 10069 11398
rect 10011 11330 10069 11364
rect 10045 11296 10069 11330
rect 9637 11247 9703 11291
rect 10011 11247 10069 11296
rect 9442 11213 9471 11247
rect 9505 11213 9563 11247
rect 9597 11213 9655 11247
rect 9689 11213 9747 11247
rect 9781 11213 9839 11247
rect 9873 11213 9931 11247
rect 9965 11213 10023 11247
rect 10057 11213 10086 11247
rect 9540 11013 9569 11047
rect 9603 11013 9661 11047
rect 9695 11013 9753 11047
rect 9787 11013 9845 11047
rect 9879 11013 9937 11047
rect 9971 11013 10000 11047
rect 9597 10929 9653 11013
rect 9787 10971 9853 11013
rect 9597 10895 9611 10929
rect 9645 10895 9653 10929
rect 9597 10879 9653 10895
rect 9687 10929 9747 10945
rect 9687 10895 9695 10929
rect 9729 10895 9747 10929
rect 9687 10835 9747 10895
rect 9787 10937 9803 10971
rect 9837 10937 9853 10971
rect 9787 10903 9853 10937
rect 9787 10869 9803 10903
rect 9837 10869 9853 10903
rect 9891 10971 9983 10979
rect 9891 10937 9907 10971
rect 9941 10937 9983 10971
rect 9891 10903 9983 10937
rect 9891 10869 9907 10903
rect 9941 10869 9983 10903
rect 9560 10758 9613 10823
rect 9687 10801 9875 10835
rect 9560 10718 9562 10758
rect 9604 10751 9613 10758
rect 9841 10751 9875 10801
rect 9604 10735 9695 10751
rect 9604 10718 9614 10735
rect 9560 10701 9614 10718
rect 9648 10701 9695 10735
rect 9739 10748 9807 10751
rect 9739 10708 9752 10748
rect 9794 10708 9807 10748
rect 9739 10701 9755 10708
rect 9789 10701 9807 10708
rect 9841 10735 9899 10751
rect 9841 10701 9863 10735
rect 9897 10701 9899 10735
rect 9841 10685 9899 10701
rect 9933 10714 9983 10869
rect 9841 10667 9875 10685
rect 9597 10629 9875 10667
rect 9933 10678 9944 10714
rect 9978 10678 9983 10714
rect 9597 10607 9663 10629
rect 9597 10573 9611 10607
rect 9645 10573 9663 10607
rect 9933 10595 9983 10678
rect 9597 10557 9663 10573
rect 9787 10579 9837 10595
rect 9787 10545 9803 10579
rect 9787 10503 9837 10545
rect 9871 10579 9983 10595
rect 9871 10545 9887 10579
rect 9921 10545 9983 10579
rect 9871 10537 9983 10545
rect 9540 10469 9569 10503
rect 9603 10469 9661 10503
rect 9695 10469 9753 10503
rect 9787 10469 9845 10503
rect 9879 10469 9937 10503
rect 9971 10469 10000 10503
rect 6112 6583 6141 6617
rect 6175 6583 6233 6617
rect 6267 6583 6325 6617
rect 6359 6583 6388 6617
rect 6178 6537 6244 6549
rect 6178 6503 6194 6537
rect 6228 6503 6244 6537
rect 6178 6469 6244 6503
rect 6178 6435 6194 6469
rect 6228 6435 6244 6469
rect 6178 6423 6244 6435
rect 6278 6537 6324 6583
rect 6312 6503 6324 6537
rect 6278 6469 6324 6503
rect 6312 6435 6324 6469
rect 6178 6382 6224 6423
rect 6278 6419 6324 6435
rect 6212 6348 6224 6382
rect 6178 6303 6224 6348
rect 6258 6350 6274 6385
rect 6308 6350 6324 6385
rect 6258 6337 6324 6350
rect 6178 6285 6244 6303
rect 6178 6251 6194 6285
rect 6228 6251 6244 6285
rect 6178 6217 6244 6251
rect 6178 6183 6194 6217
rect 6228 6183 6244 6217
rect 6178 6149 6244 6183
rect 6178 6115 6194 6149
rect 6228 6115 6244 6149
rect 6178 6107 6244 6115
rect 6278 6285 6320 6301
rect 6312 6251 6320 6285
rect 6278 6217 6320 6251
rect 6312 6183 6320 6217
rect 6278 6149 6320 6183
rect 6312 6115 6320 6149
rect 6278 6073 6320 6115
rect 6112 6039 6141 6073
rect 6175 6039 6233 6073
rect 6267 6039 6325 6073
rect 6359 6039 6388 6073
rect 9218 5951 9247 5985
rect 9281 5951 9339 5985
rect 9373 5951 9431 5985
rect 9465 5951 9523 5985
rect 9557 5951 9615 5985
rect 9649 5951 9707 5985
rect 9741 5951 9799 5985
rect 9833 5951 9891 5985
rect 9925 5951 9983 5985
rect 10017 5951 10075 5985
rect 10109 5951 10167 5985
rect 10201 5951 10259 5985
rect 10293 5951 10351 5985
rect 10385 5951 10443 5985
rect 10477 5951 10535 5985
rect 10569 5951 10627 5985
rect 10661 5951 10690 5985
rect 9242 5873 9322 5917
rect 9371 5913 9437 5951
rect 9371 5879 9387 5913
rect 9421 5879 9437 5913
rect 9471 5901 9673 5917
rect 9242 5839 9288 5873
rect 9471 5867 9639 5901
rect 9471 5845 9505 5867
rect 9639 5849 9673 5867
rect 9740 5896 9774 5917
rect 9808 5913 9874 5951
rect 9808 5879 9824 5913
rect 9858 5879 9874 5913
rect 9908 5896 9942 5917
rect 9242 5806 9322 5839
rect 9357 5811 9505 5845
rect 9740 5845 9774 5862
rect 9976 5904 10042 5951
rect 9976 5870 9992 5904
rect 10026 5870 10042 5904
rect 10096 5896 10130 5917
rect 9908 5845 9942 5862
rect 9242 5671 9308 5806
rect 9357 5769 9391 5811
rect 9342 5753 9391 5769
rect 9598 5781 9610 5815
rect 9644 5781 9697 5815
rect 9740 5811 9942 5845
rect 10164 5913 10230 5951
rect 10164 5879 10180 5913
rect 10214 5879 10230 5913
rect 10264 5896 10298 5917
rect 10096 5845 10130 5862
rect 10264 5845 10298 5862
rect 10096 5811 10298 5845
rect 10348 5896 10468 5917
rect 10382 5862 10468 5896
rect 10521 5909 10587 5951
rect 11088 5947 11117 5981
rect 11151 5947 11209 5981
rect 11243 5947 11301 5981
rect 11335 5947 11393 5981
rect 11427 5947 11485 5981
rect 11519 5947 11577 5981
rect 11611 5947 11669 5981
rect 11703 5947 11761 5981
rect 11795 5947 11853 5981
rect 11887 5947 11945 5981
rect 11979 5947 12037 5981
rect 12071 5947 12129 5981
rect 12163 5947 12221 5981
rect 12255 5947 12313 5981
rect 12347 5947 12405 5981
rect 12439 5947 12497 5981
rect 12531 5947 12560 5981
rect 10521 5875 10537 5909
rect 10571 5875 10587 5909
rect 10348 5841 10468 5862
rect 10621 5873 10673 5917
rect 10348 5815 10587 5841
rect 10348 5781 10350 5815
rect 10384 5807 10587 5815
rect 10384 5781 10396 5807
rect 9598 5777 9697 5781
rect 9376 5719 9391 5753
rect 9342 5703 9391 5719
rect 9425 5747 9441 5761
rect 9425 5713 9426 5747
rect 9475 5727 9513 5761
rect 9598 5743 9681 5777
rect 9715 5743 9731 5777
rect 9765 5743 9781 5777
rect 9815 5747 9840 5777
rect 9460 5713 9513 5727
rect 9765 5713 9794 5743
rect 9828 5713 9840 5747
rect 9899 5718 10132 5775
rect 10553 5769 10587 5807
rect 10655 5839 10673 5873
rect 10621 5802 10673 5839
rect 9242 5633 9322 5671
rect 9242 5599 9288 5633
rect 1836 5531 1865 5565
rect 1899 5531 1957 5565
rect 1991 5531 2049 5565
rect 2083 5531 2141 5565
rect 2175 5531 2233 5565
rect 2267 5531 2325 5565
rect 2359 5531 2417 5565
rect 2451 5531 2509 5565
rect 2543 5531 2601 5565
rect 2635 5531 2693 5565
rect 2727 5531 2785 5565
rect 2819 5531 2877 5565
rect 2911 5531 2969 5565
rect 3003 5531 3061 5565
rect 3095 5531 3153 5565
rect 3187 5531 3245 5565
rect 3279 5531 3308 5565
rect 1860 5453 1940 5497
rect 1989 5493 2055 5531
rect 1989 5459 2005 5493
rect 2039 5459 2055 5493
rect 2089 5481 2291 5497
rect 1860 5419 1906 5453
rect 2089 5447 2257 5481
rect 2089 5425 2123 5447
rect 2257 5429 2291 5447
rect 2358 5476 2392 5497
rect 2426 5493 2492 5531
rect 2426 5459 2442 5493
rect 2476 5459 2492 5493
rect 2526 5476 2560 5497
rect 1860 5386 1940 5419
rect 1975 5391 2123 5425
rect 2358 5425 2392 5442
rect 2594 5484 2660 5531
rect 2594 5450 2610 5484
rect 2644 5450 2660 5484
rect 2714 5476 2748 5497
rect 2526 5425 2560 5442
rect 1860 5251 1926 5386
rect 1975 5349 2009 5391
rect 1960 5333 2009 5349
rect 2216 5361 2228 5395
rect 2262 5361 2315 5395
rect 2358 5391 2560 5425
rect 2782 5493 2848 5531
rect 2782 5459 2798 5493
rect 2832 5459 2848 5493
rect 2882 5476 2916 5497
rect 2714 5425 2748 5442
rect 2882 5425 2916 5442
rect 2714 5391 2916 5425
rect 2966 5476 3086 5497
rect 3000 5442 3086 5476
rect 3139 5489 3205 5531
rect 3706 5527 3735 5561
rect 3769 5527 3827 5561
rect 3861 5527 3919 5561
rect 3953 5527 4011 5561
rect 4045 5527 4103 5561
rect 4137 5527 4195 5561
rect 4229 5527 4287 5561
rect 4321 5527 4379 5561
rect 4413 5527 4471 5561
rect 4505 5527 4563 5561
rect 4597 5527 4655 5561
rect 4689 5527 4747 5561
rect 4781 5527 4839 5561
rect 4873 5527 4931 5561
rect 4965 5527 5023 5561
rect 5057 5527 5115 5561
rect 5149 5527 5178 5561
rect 3139 5455 3155 5489
rect 3189 5455 3205 5489
rect 2966 5421 3086 5442
rect 3239 5453 3291 5497
rect 2966 5395 3205 5421
rect 2966 5361 2968 5395
rect 3002 5387 3205 5395
rect 3002 5361 3014 5387
rect 2216 5357 2315 5361
rect 1994 5299 2009 5333
rect 1960 5283 2009 5299
rect 2043 5327 2059 5341
rect 2043 5293 2044 5327
rect 2093 5307 2131 5341
rect 2216 5323 2299 5357
rect 2333 5323 2349 5357
rect 2383 5323 2399 5357
rect 2433 5327 2458 5357
rect 2078 5293 2131 5307
rect 2383 5293 2412 5323
rect 2446 5293 2458 5327
rect 2517 5298 2750 5355
rect 3171 5349 3205 5387
rect 3273 5419 3291 5453
rect 3239 5382 3291 5419
rect 1860 5213 1940 5251
rect 1860 5179 1906 5213
rect 1860 5123 1940 5179
rect 1975 5161 2009 5283
rect 2097 5229 2136 5259
rect 2097 5195 2131 5229
rect 2170 5225 2181 5259
rect 2517 5245 2551 5298
rect 2165 5195 2181 5225
rect 2227 5229 2484 5245
rect 2261 5211 2484 5229
rect 2518 5211 2551 5245
rect 2596 5259 2668 5261
rect 2630 5245 2668 5259
rect 2596 5211 2601 5225
rect 2635 5211 2668 5245
rect 2261 5195 2277 5211
rect 2596 5195 2668 5211
rect 2716 5229 2750 5298
rect 2784 5327 2862 5342
rect 3060 5333 3126 5349
rect 3060 5327 3092 5333
rect 2818 5326 2862 5327
rect 2818 5293 2828 5326
rect 2784 5292 2828 5293
rect 2784 5276 2862 5292
rect 2900 5293 2924 5327
rect 2958 5293 2974 5327
rect 3094 5293 3126 5299
rect 2900 5229 2934 5293
rect 3092 5283 3126 5293
rect 3171 5333 3222 5349
rect 3171 5299 3188 5333
rect 3171 5283 3222 5299
rect 2716 5195 2934 5229
rect 3002 5225 3048 5259
rect 2968 5222 3048 5225
rect 3171 5223 3205 5283
rect 3256 5251 3291 5382
rect 2227 5194 2277 5195
rect 1975 5127 2108 5161
rect 2227 5160 2236 5194
rect 2270 5160 2277 5194
rect 2968 5188 3014 5222
rect 2968 5172 3048 5188
rect 2227 5157 2277 5160
rect 1860 5089 1906 5123
rect 2074 5123 2108 5127
rect 2358 5127 2560 5161
rect 2074 5105 2291 5123
rect 1860 5055 1940 5089
rect 1974 5059 1990 5093
rect 2024 5059 2040 5093
rect 1974 5021 2040 5059
rect 2074 5071 2257 5105
rect 2074 5055 2291 5071
rect 2358 5110 2392 5127
rect 2526 5110 2560 5127
rect 2358 5055 2392 5076
rect 2426 5059 2442 5093
rect 2476 5059 2492 5093
rect 2426 5021 2492 5059
rect 2701 5127 2916 5161
rect 3087 5159 3205 5223
rect 3239 5210 3291 5251
rect 3273 5186 3291 5210
rect 3087 5135 3121 5159
rect 2701 5110 2748 5127
rect 2526 5055 2560 5076
rect 2594 5063 2610 5097
rect 2644 5063 2660 5097
rect 2594 5021 2660 5063
rect 2701 5076 2714 5110
rect 2882 5110 2916 5127
rect 2701 5055 2748 5076
rect 2782 5059 2798 5093
rect 2832 5059 2848 5093
rect 2782 5021 2848 5059
rect 2882 5055 2916 5076
rect 2966 5110 3121 5135
rect 3239 5150 3244 5176
rect 3284 5150 3291 5186
rect 3000 5076 3121 5110
rect 2966 5055 3121 5076
rect 3155 5101 3205 5118
rect 3189 5067 3205 5101
rect 3155 5021 3205 5067
rect 3239 5116 3291 5150
rect 3273 5082 3291 5116
rect 3239 5055 3291 5082
rect 3730 5449 3810 5493
rect 3859 5489 3925 5527
rect 3859 5455 3875 5489
rect 3909 5455 3925 5489
rect 3959 5477 4161 5493
rect 3730 5415 3776 5449
rect 3959 5443 4127 5477
rect 3959 5421 3993 5443
rect 4127 5425 4161 5443
rect 4228 5472 4262 5493
rect 4296 5489 4362 5527
rect 4296 5455 4312 5489
rect 4346 5455 4362 5489
rect 4396 5472 4430 5493
rect 3730 5382 3810 5415
rect 3845 5387 3993 5421
rect 4228 5421 4262 5438
rect 4464 5480 4530 5527
rect 4464 5446 4480 5480
rect 4514 5446 4530 5480
rect 4584 5472 4618 5493
rect 4396 5421 4430 5438
rect 3730 5247 3796 5382
rect 3845 5345 3879 5387
rect 3830 5329 3879 5345
rect 4086 5357 4098 5391
rect 4132 5357 4185 5391
rect 4228 5387 4430 5421
rect 4652 5489 4718 5527
rect 4652 5455 4668 5489
rect 4702 5455 4718 5489
rect 4752 5472 4786 5493
rect 4584 5421 4618 5438
rect 4752 5421 4786 5438
rect 4584 5387 4786 5421
rect 4836 5472 4956 5493
rect 4870 5438 4956 5472
rect 5009 5485 5075 5527
rect 5522 5523 5551 5557
rect 5585 5523 5643 5557
rect 5677 5523 5735 5557
rect 5769 5523 5827 5557
rect 5861 5523 5919 5557
rect 5953 5523 6011 5557
rect 6045 5523 6103 5557
rect 6137 5523 6195 5557
rect 6229 5523 6287 5557
rect 6321 5523 6379 5557
rect 6413 5523 6471 5557
rect 6505 5523 6563 5557
rect 6597 5523 6655 5557
rect 6689 5523 6747 5557
rect 6781 5523 6839 5557
rect 6873 5523 6931 5557
rect 6965 5523 6994 5557
rect 5009 5451 5025 5485
rect 5059 5451 5075 5485
rect 4836 5417 4956 5438
rect 5109 5449 5161 5493
rect 4836 5391 5075 5417
rect 4836 5357 4838 5391
rect 4872 5383 5075 5391
rect 4872 5357 4884 5383
rect 4086 5353 4185 5357
rect 3864 5295 3879 5329
rect 3830 5279 3879 5295
rect 3913 5323 3929 5337
rect 3913 5289 3914 5323
rect 3963 5303 4001 5337
rect 4086 5319 4169 5353
rect 4203 5319 4219 5353
rect 4253 5319 4269 5353
rect 4303 5323 4328 5353
rect 3948 5289 4001 5303
rect 4253 5289 4282 5319
rect 4316 5289 4328 5323
rect 4387 5294 4620 5351
rect 5041 5345 5075 5383
rect 5143 5415 5161 5449
rect 5109 5378 5161 5415
rect 3730 5209 3810 5247
rect 3730 5175 3776 5209
rect 3730 5119 3810 5175
rect 3845 5157 3879 5279
rect 3967 5225 4006 5255
rect 3967 5191 4001 5225
rect 4040 5221 4051 5255
rect 4387 5241 4421 5294
rect 4035 5191 4051 5221
rect 4097 5225 4354 5241
rect 4131 5207 4354 5225
rect 4388 5207 4421 5241
rect 4466 5255 4538 5257
rect 4500 5241 4538 5255
rect 4466 5207 4471 5221
rect 4505 5207 4538 5241
rect 4131 5191 4147 5207
rect 4466 5191 4538 5207
rect 4586 5225 4620 5294
rect 4654 5323 4732 5338
rect 4930 5329 4996 5345
rect 4930 5323 4962 5329
rect 4688 5322 4732 5323
rect 4688 5289 4698 5322
rect 4654 5288 4698 5289
rect 4654 5272 4732 5288
rect 4770 5289 4794 5323
rect 4828 5289 4844 5323
rect 4964 5289 4996 5295
rect 4770 5225 4804 5289
rect 4962 5279 4996 5289
rect 5041 5329 5092 5345
rect 5041 5295 5058 5329
rect 5041 5279 5092 5295
rect 4586 5191 4804 5225
rect 4872 5221 4918 5255
rect 4838 5218 4918 5221
rect 5041 5219 5075 5279
rect 5126 5247 5161 5378
rect 4097 5188 4147 5191
rect 3845 5123 3978 5157
rect 4097 5154 4104 5188
rect 4138 5154 4147 5188
rect 4838 5184 4884 5218
rect 4838 5168 4918 5184
rect 4097 5153 4147 5154
rect 3730 5085 3776 5119
rect 3944 5119 3978 5123
rect 4228 5123 4430 5157
rect 3944 5101 4161 5119
rect 3730 5051 3810 5085
rect 3844 5055 3860 5089
rect 3894 5055 3910 5089
rect 1836 4987 1865 5021
rect 1899 4987 1957 5021
rect 1991 4987 2049 5021
rect 2083 4987 2141 5021
rect 2175 4987 2233 5021
rect 2267 4987 2325 5021
rect 2359 4987 2417 5021
rect 2451 4987 2509 5021
rect 2543 4987 2601 5021
rect 2635 4987 2693 5021
rect 2727 4987 2785 5021
rect 2819 4987 2877 5021
rect 2911 4987 2969 5021
rect 3003 4987 3061 5021
rect 3095 4987 3153 5021
rect 3187 4987 3245 5021
rect 3279 4987 3308 5021
rect 3844 5017 3910 5055
rect 3944 5067 4127 5101
rect 3944 5051 4161 5067
rect 4228 5106 4262 5123
rect 4396 5106 4430 5123
rect 4228 5051 4262 5072
rect 4296 5055 4312 5089
rect 4346 5055 4362 5089
rect 4296 5017 4362 5055
rect 4571 5123 4786 5157
rect 4957 5155 5075 5219
rect 5109 5206 5161 5247
rect 5143 5182 5161 5206
rect 4957 5131 4991 5155
rect 4571 5106 4618 5123
rect 4396 5051 4430 5072
rect 4464 5059 4480 5093
rect 4514 5059 4530 5093
rect 4464 5017 4530 5059
rect 4571 5072 4584 5106
rect 4752 5106 4786 5123
rect 4571 5051 4618 5072
rect 4652 5055 4668 5089
rect 4702 5055 4718 5089
rect 4652 5017 4718 5055
rect 4752 5051 4786 5072
rect 4836 5106 4991 5131
rect 5109 5144 5120 5172
rect 5156 5144 5161 5182
rect 4870 5072 4991 5106
rect 4836 5051 4991 5072
rect 5025 5097 5075 5114
rect 5059 5063 5075 5097
rect 5025 5017 5075 5063
rect 5109 5112 5161 5144
rect 5143 5078 5161 5112
rect 5109 5051 5161 5078
rect 5546 5445 5626 5489
rect 5675 5485 5741 5523
rect 5675 5451 5691 5485
rect 5725 5451 5741 5485
rect 5775 5473 5977 5489
rect 5546 5411 5592 5445
rect 5775 5439 5943 5473
rect 5775 5417 5809 5439
rect 5943 5421 5977 5439
rect 6044 5468 6078 5489
rect 6112 5485 6178 5523
rect 6112 5451 6128 5485
rect 6162 5451 6178 5485
rect 6212 5468 6246 5489
rect 5546 5378 5626 5411
rect 5661 5383 5809 5417
rect 6044 5417 6078 5434
rect 6280 5476 6346 5523
rect 6280 5442 6296 5476
rect 6330 5442 6346 5476
rect 6400 5468 6434 5489
rect 6212 5417 6246 5434
rect 5546 5243 5612 5378
rect 5661 5341 5695 5383
rect 5646 5325 5695 5341
rect 5902 5353 5914 5387
rect 5948 5353 6001 5387
rect 6044 5383 6246 5417
rect 6468 5485 6534 5523
rect 6468 5451 6484 5485
rect 6518 5451 6534 5485
rect 6568 5468 6602 5489
rect 6400 5417 6434 5434
rect 6568 5417 6602 5434
rect 6400 5383 6602 5417
rect 6652 5468 6772 5489
rect 6686 5434 6772 5468
rect 6825 5481 6891 5523
rect 7392 5519 7421 5553
rect 7455 5519 7513 5553
rect 7547 5519 7605 5553
rect 7639 5519 7697 5553
rect 7731 5519 7789 5553
rect 7823 5519 7881 5553
rect 7915 5519 7973 5553
rect 8007 5519 8065 5553
rect 8099 5519 8157 5553
rect 8191 5519 8249 5553
rect 8283 5519 8341 5553
rect 8375 5519 8433 5553
rect 8467 5519 8525 5553
rect 8559 5519 8617 5553
rect 8651 5519 8709 5553
rect 8743 5519 8801 5553
rect 8835 5519 8864 5553
rect 9242 5543 9322 5599
rect 9357 5581 9391 5703
rect 9479 5649 9518 5679
rect 9479 5615 9513 5649
rect 9552 5645 9563 5679
rect 9899 5665 9933 5718
rect 9547 5615 9563 5645
rect 9609 5649 9866 5665
rect 9643 5631 9866 5649
rect 9900 5631 9933 5665
rect 9978 5679 10050 5681
rect 10012 5665 10050 5679
rect 9978 5631 9983 5645
rect 10017 5631 10050 5665
rect 9643 5615 9659 5631
rect 9978 5615 10050 5631
rect 10098 5649 10132 5718
rect 10166 5747 10244 5762
rect 10442 5753 10508 5769
rect 10442 5747 10474 5753
rect 10200 5746 10244 5747
rect 10200 5713 10210 5746
rect 10166 5712 10210 5713
rect 10166 5696 10244 5712
rect 10282 5713 10306 5747
rect 10340 5713 10356 5747
rect 10476 5713 10508 5719
rect 10282 5649 10316 5713
rect 10474 5703 10508 5713
rect 10553 5753 10604 5769
rect 10553 5719 10570 5753
rect 10553 5703 10604 5719
rect 10098 5615 10316 5649
rect 10384 5645 10430 5679
rect 10350 5642 10430 5645
rect 10553 5643 10587 5703
rect 10638 5671 10673 5802
rect 9609 5614 9659 5615
rect 9357 5547 9490 5581
rect 9609 5580 9618 5614
rect 9652 5580 9659 5614
rect 10350 5608 10396 5642
rect 10350 5592 10430 5608
rect 9609 5577 9659 5580
rect 6825 5447 6841 5481
rect 6875 5447 6891 5481
rect 6652 5413 6772 5434
rect 6925 5445 6977 5489
rect 6652 5387 6891 5413
rect 6652 5353 6654 5387
rect 6688 5379 6891 5387
rect 6688 5353 6700 5379
rect 5902 5349 6001 5353
rect 5680 5291 5695 5325
rect 5646 5275 5695 5291
rect 5729 5319 5745 5333
rect 5729 5285 5730 5319
rect 5779 5299 5817 5333
rect 5902 5315 5985 5349
rect 6019 5315 6035 5349
rect 6069 5315 6085 5349
rect 6119 5319 6144 5349
rect 5764 5285 5817 5299
rect 6069 5285 6098 5315
rect 6132 5285 6144 5319
rect 6203 5290 6436 5347
rect 6857 5341 6891 5379
rect 6959 5411 6977 5445
rect 6925 5374 6977 5411
rect 5546 5205 5626 5243
rect 5546 5171 5592 5205
rect 5546 5115 5626 5171
rect 5661 5153 5695 5275
rect 5783 5221 5822 5251
rect 5783 5187 5817 5221
rect 5856 5217 5867 5251
rect 6203 5237 6237 5290
rect 5851 5187 5867 5217
rect 5913 5221 6170 5237
rect 5947 5203 6170 5221
rect 6204 5203 6237 5237
rect 6282 5251 6354 5253
rect 6316 5237 6354 5251
rect 6282 5203 6287 5217
rect 6321 5203 6354 5237
rect 5947 5187 5963 5203
rect 6282 5187 6354 5203
rect 6402 5221 6436 5290
rect 6470 5319 6548 5334
rect 6746 5325 6812 5341
rect 6746 5319 6778 5325
rect 6504 5318 6548 5319
rect 6504 5285 6514 5318
rect 6470 5284 6514 5285
rect 6470 5268 6548 5284
rect 6586 5285 6610 5319
rect 6644 5285 6660 5319
rect 6780 5285 6812 5291
rect 6586 5221 6620 5285
rect 6778 5275 6812 5285
rect 6857 5325 6908 5341
rect 6857 5291 6874 5325
rect 6857 5275 6908 5291
rect 6402 5187 6620 5221
rect 6688 5217 6734 5251
rect 6654 5214 6734 5217
rect 6857 5215 6891 5275
rect 6942 5243 6977 5374
rect 5913 5184 5963 5187
rect 5661 5119 5794 5153
rect 5913 5150 5920 5184
rect 5954 5150 5963 5184
rect 6654 5180 6700 5214
rect 6654 5164 6734 5180
rect 5913 5149 5963 5150
rect 5546 5081 5592 5115
rect 5760 5115 5794 5119
rect 6044 5119 6246 5153
rect 5760 5097 5977 5115
rect 5546 5047 5626 5081
rect 5660 5051 5676 5085
rect 5710 5051 5726 5085
rect 3706 4983 3735 5017
rect 3769 4983 3827 5017
rect 3861 4983 3919 5017
rect 3953 4983 4011 5017
rect 4045 4983 4103 5017
rect 4137 4983 4195 5017
rect 4229 4983 4287 5017
rect 4321 4983 4379 5017
rect 4413 4983 4471 5017
rect 4505 4983 4563 5017
rect 4597 4983 4655 5017
rect 4689 4983 4747 5017
rect 4781 4983 4839 5017
rect 4873 4983 4931 5017
rect 4965 4983 5023 5017
rect 5057 4983 5115 5017
rect 5149 4983 5178 5017
rect 5660 5013 5726 5051
rect 5760 5063 5943 5097
rect 5760 5047 5977 5063
rect 6044 5102 6078 5119
rect 6212 5102 6246 5119
rect 6044 5047 6078 5068
rect 6112 5051 6128 5085
rect 6162 5051 6178 5085
rect 6112 5013 6178 5051
rect 6387 5119 6602 5153
rect 6773 5151 6891 5215
rect 6925 5202 6977 5243
rect 6959 5178 6977 5202
rect 6773 5127 6807 5151
rect 6387 5102 6434 5119
rect 6212 5047 6246 5068
rect 6280 5055 6296 5089
rect 6330 5055 6346 5089
rect 6280 5013 6346 5055
rect 6387 5068 6400 5102
rect 6568 5102 6602 5119
rect 6387 5047 6434 5068
rect 6468 5051 6484 5085
rect 6518 5051 6534 5085
rect 6468 5013 6534 5051
rect 6568 5047 6602 5068
rect 6652 5102 6807 5127
rect 6925 5142 6930 5168
rect 6970 5142 6977 5178
rect 6686 5068 6807 5102
rect 6652 5047 6807 5068
rect 6841 5093 6891 5110
rect 6875 5059 6891 5093
rect 6841 5013 6891 5059
rect 6925 5108 6977 5142
rect 6959 5074 6977 5108
rect 6925 5047 6977 5074
rect 7416 5441 7496 5485
rect 7545 5481 7611 5519
rect 7545 5447 7561 5481
rect 7595 5447 7611 5481
rect 7645 5469 7847 5485
rect 7416 5407 7462 5441
rect 7645 5435 7813 5469
rect 7645 5413 7679 5435
rect 7813 5417 7847 5435
rect 7914 5464 7948 5485
rect 7982 5481 8048 5519
rect 7982 5447 7998 5481
rect 8032 5447 8048 5481
rect 8082 5464 8116 5485
rect 7416 5374 7496 5407
rect 7531 5379 7679 5413
rect 7914 5413 7948 5430
rect 8150 5472 8216 5519
rect 8150 5438 8166 5472
rect 8200 5438 8216 5472
rect 8270 5464 8304 5485
rect 8082 5413 8116 5430
rect 7416 5239 7482 5374
rect 7531 5337 7565 5379
rect 7516 5321 7565 5337
rect 7772 5349 7784 5383
rect 7818 5349 7871 5383
rect 7914 5379 8116 5413
rect 8338 5481 8404 5519
rect 8338 5447 8354 5481
rect 8388 5447 8404 5481
rect 8438 5464 8472 5485
rect 8270 5413 8304 5430
rect 8438 5413 8472 5430
rect 8270 5379 8472 5413
rect 8522 5464 8642 5485
rect 8556 5430 8642 5464
rect 8695 5477 8761 5519
rect 9242 5509 9288 5543
rect 9456 5543 9490 5547
rect 9740 5547 9942 5581
rect 9456 5525 9673 5543
rect 8695 5443 8711 5477
rect 8745 5443 8761 5477
rect 8522 5409 8642 5430
rect 8795 5441 8847 5485
rect 9242 5475 9322 5509
rect 9356 5479 9372 5513
rect 9406 5479 9422 5513
rect 9356 5441 9422 5479
rect 9456 5491 9639 5525
rect 9456 5475 9673 5491
rect 9740 5530 9774 5547
rect 9908 5530 9942 5547
rect 9740 5475 9774 5496
rect 9808 5479 9824 5513
rect 9858 5479 9874 5513
rect 9808 5441 9874 5479
rect 10083 5547 10298 5581
rect 10469 5579 10587 5643
rect 10621 5630 10673 5671
rect 10655 5606 10673 5630
rect 10469 5555 10503 5579
rect 10083 5530 10130 5547
rect 9908 5475 9942 5496
rect 9976 5483 9992 5517
rect 10026 5483 10042 5517
rect 9976 5441 10042 5483
rect 10083 5496 10096 5530
rect 10264 5530 10298 5547
rect 10083 5475 10130 5496
rect 10164 5479 10180 5513
rect 10214 5479 10230 5513
rect 10164 5441 10230 5479
rect 10264 5475 10298 5496
rect 10348 5530 10503 5555
rect 10621 5570 10626 5596
rect 10666 5570 10673 5606
rect 10382 5496 10503 5530
rect 10348 5475 10503 5496
rect 10537 5521 10587 5538
rect 10571 5487 10587 5521
rect 10537 5441 10587 5487
rect 10621 5536 10673 5570
rect 10655 5502 10673 5536
rect 10621 5475 10673 5502
rect 11112 5869 11192 5913
rect 11241 5909 11307 5947
rect 11241 5875 11257 5909
rect 11291 5875 11307 5909
rect 11341 5897 11543 5913
rect 11112 5835 11158 5869
rect 11341 5863 11509 5897
rect 11341 5841 11375 5863
rect 11509 5845 11543 5863
rect 11610 5892 11644 5913
rect 11678 5909 11744 5947
rect 11678 5875 11694 5909
rect 11728 5875 11744 5909
rect 11778 5892 11812 5913
rect 11112 5802 11192 5835
rect 11227 5807 11375 5841
rect 11610 5841 11644 5858
rect 11846 5900 11912 5947
rect 11846 5866 11862 5900
rect 11896 5866 11912 5900
rect 11966 5892 12000 5913
rect 11778 5841 11812 5858
rect 11112 5667 11178 5802
rect 11227 5765 11261 5807
rect 11212 5749 11261 5765
rect 11468 5777 11480 5811
rect 11514 5777 11567 5811
rect 11610 5807 11812 5841
rect 12034 5909 12100 5947
rect 12034 5875 12050 5909
rect 12084 5875 12100 5909
rect 12134 5892 12168 5913
rect 11966 5841 12000 5858
rect 12134 5841 12168 5858
rect 11966 5807 12168 5841
rect 12218 5892 12338 5913
rect 12252 5858 12338 5892
rect 12391 5905 12457 5947
rect 12904 5943 12933 5977
rect 12967 5943 13025 5977
rect 13059 5943 13117 5977
rect 13151 5943 13209 5977
rect 13243 5943 13301 5977
rect 13335 5943 13393 5977
rect 13427 5943 13485 5977
rect 13519 5943 13577 5977
rect 13611 5943 13669 5977
rect 13703 5943 13761 5977
rect 13795 5943 13853 5977
rect 13887 5943 13945 5977
rect 13979 5943 14037 5977
rect 14071 5943 14129 5977
rect 14163 5943 14221 5977
rect 14255 5943 14313 5977
rect 14347 5943 14376 5977
rect 12391 5871 12407 5905
rect 12441 5871 12457 5905
rect 12218 5837 12338 5858
rect 12491 5869 12543 5913
rect 12218 5811 12457 5837
rect 12218 5777 12220 5811
rect 12254 5803 12457 5811
rect 12254 5777 12266 5803
rect 11468 5773 11567 5777
rect 11246 5715 11261 5749
rect 11212 5699 11261 5715
rect 11295 5743 11311 5757
rect 11295 5709 11296 5743
rect 11345 5723 11383 5757
rect 11468 5739 11551 5773
rect 11585 5739 11601 5773
rect 11635 5739 11651 5773
rect 11685 5743 11710 5773
rect 11330 5709 11383 5723
rect 11635 5709 11664 5739
rect 11698 5709 11710 5743
rect 11769 5714 12002 5771
rect 12423 5765 12457 5803
rect 12525 5835 12543 5869
rect 12491 5798 12543 5835
rect 11112 5629 11192 5667
rect 11112 5595 11158 5629
rect 11112 5539 11192 5595
rect 11227 5577 11261 5699
rect 11349 5645 11388 5675
rect 11349 5611 11383 5645
rect 11422 5641 11433 5675
rect 11769 5661 11803 5714
rect 11417 5611 11433 5641
rect 11479 5645 11736 5661
rect 11513 5627 11736 5645
rect 11770 5627 11803 5661
rect 11848 5675 11920 5677
rect 11882 5661 11920 5675
rect 11848 5627 11853 5641
rect 11887 5627 11920 5661
rect 11513 5611 11529 5627
rect 11848 5611 11920 5627
rect 11968 5645 12002 5714
rect 12036 5743 12114 5758
rect 12312 5749 12378 5765
rect 12312 5743 12344 5749
rect 12070 5742 12114 5743
rect 12070 5709 12080 5742
rect 12036 5708 12080 5709
rect 12036 5692 12114 5708
rect 12152 5709 12176 5743
rect 12210 5709 12226 5743
rect 12346 5709 12378 5715
rect 12152 5645 12186 5709
rect 12344 5699 12378 5709
rect 12423 5749 12474 5765
rect 12423 5715 12440 5749
rect 12423 5699 12474 5715
rect 11968 5611 12186 5645
rect 12254 5641 12300 5675
rect 12220 5638 12300 5641
rect 12423 5639 12457 5699
rect 12508 5667 12543 5798
rect 11479 5608 11529 5611
rect 11227 5543 11360 5577
rect 11479 5574 11486 5608
rect 11520 5574 11529 5608
rect 12220 5604 12266 5638
rect 12220 5588 12300 5604
rect 11479 5573 11529 5574
rect 11112 5505 11158 5539
rect 11326 5539 11360 5543
rect 11610 5543 11812 5577
rect 11326 5521 11543 5539
rect 11112 5471 11192 5505
rect 11226 5475 11242 5509
rect 11276 5475 11292 5509
rect 8522 5383 8761 5409
rect 8522 5349 8524 5383
rect 8558 5375 8761 5383
rect 8558 5349 8570 5375
rect 7772 5345 7871 5349
rect 7550 5287 7565 5321
rect 7516 5271 7565 5287
rect 7599 5315 7615 5329
rect 7599 5281 7600 5315
rect 7649 5295 7687 5329
rect 7772 5311 7855 5345
rect 7889 5311 7905 5345
rect 7939 5311 7955 5345
rect 7989 5315 8014 5345
rect 7634 5281 7687 5295
rect 7939 5281 7968 5311
rect 8002 5281 8014 5315
rect 8073 5286 8306 5343
rect 8727 5337 8761 5375
rect 8829 5407 8847 5441
rect 9218 5407 9247 5441
rect 9281 5407 9339 5441
rect 9373 5407 9431 5441
rect 9465 5407 9523 5441
rect 9557 5407 9615 5441
rect 9649 5407 9707 5441
rect 9741 5407 9799 5441
rect 9833 5407 9891 5441
rect 9925 5407 9983 5441
rect 10017 5407 10075 5441
rect 10109 5407 10167 5441
rect 10201 5407 10259 5441
rect 10293 5407 10351 5441
rect 10385 5407 10443 5441
rect 10477 5407 10535 5441
rect 10569 5407 10627 5441
rect 10661 5407 10690 5441
rect 11226 5437 11292 5475
rect 11326 5487 11509 5521
rect 11326 5471 11543 5487
rect 11610 5526 11644 5543
rect 11778 5526 11812 5543
rect 11610 5471 11644 5492
rect 11678 5475 11694 5509
rect 11728 5475 11744 5509
rect 11678 5437 11744 5475
rect 11953 5543 12168 5577
rect 12339 5575 12457 5639
rect 12491 5626 12543 5667
rect 12525 5602 12543 5626
rect 12339 5551 12373 5575
rect 11953 5526 12000 5543
rect 11778 5471 11812 5492
rect 11846 5479 11862 5513
rect 11896 5479 11912 5513
rect 11846 5437 11912 5479
rect 11953 5492 11966 5526
rect 12134 5526 12168 5543
rect 11953 5471 12000 5492
rect 12034 5475 12050 5509
rect 12084 5475 12100 5509
rect 12034 5437 12100 5475
rect 12134 5471 12168 5492
rect 12218 5526 12373 5551
rect 12491 5568 12502 5592
rect 12538 5568 12543 5602
rect 12252 5492 12373 5526
rect 12218 5471 12373 5492
rect 12407 5517 12457 5534
rect 12441 5483 12457 5517
rect 12407 5437 12457 5483
rect 12491 5532 12543 5568
rect 12525 5498 12543 5532
rect 12491 5471 12543 5498
rect 12928 5865 13008 5909
rect 13057 5905 13123 5943
rect 13057 5871 13073 5905
rect 13107 5871 13123 5905
rect 13157 5893 13359 5909
rect 12928 5831 12974 5865
rect 13157 5859 13325 5893
rect 13157 5837 13191 5859
rect 13325 5841 13359 5859
rect 13426 5888 13460 5909
rect 13494 5905 13560 5943
rect 13494 5871 13510 5905
rect 13544 5871 13560 5905
rect 13594 5888 13628 5909
rect 12928 5798 13008 5831
rect 13043 5803 13191 5837
rect 13426 5837 13460 5854
rect 13662 5896 13728 5943
rect 13662 5862 13678 5896
rect 13712 5862 13728 5896
rect 13782 5888 13816 5909
rect 13594 5837 13628 5854
rect 12928 5663 12994 5798
rect 13043 5761 13077 5803
rect 13028 5745 13077 5761
rect 13284 5773 13296 5807
rect 13330 5773 13383 5807
rect 13426 5803 13628 5837
rect 13850 5905 13916 5943
rect 13850 5871 13866 5905
rect 13900 5871 13916 5905
rect 13950 5888 13984 5909
rect 13782 5837 13816 5854
rect 13950 5837 13984 5854
rect 13782 5803 13984 5837
rect 14034 5888 14154 5909
rect 14068 5854 14154 5888
rect 14207 5901 14273 5943
rect 14774 5939 14803 5973
rect 14837 5939 14895 5973
rect 14929 5939 14987 5973
rect 15021 5939 15079 5973
rect 15113 5939 15171 5973
rect 15205 5939 15263 5973
rect 15297 5939 15355 5973
rect 15389 5939 15447 5973
rect 15481 5939 15539 5973
rect 15573 5939 15631 5973
rect 15665 5939 15723 5973
rect 15757 5939 15815 5973
rect 15849 5939 15907 5973
rect 15941 5939 15999 5973
rect 16033 5939 16091 5973
rect 16125 5939 16183 5973
rect 16217 5939 16246 5973
rect 14207 5867 14223 5901
rect 14257 5867 14273 5901
rect 14034 5833 14154 5854
rect 14307 5865 14359 5909
rect 14034 5807 14273 5833
rect 14034 5773 14036 5807
rect 14070 5799 14273 5807
rect 14070 5773 14082 5799
rect 13284 5769 13383 5773
rect 13062 5711 13077 5745
rect 13028 5695 13077 5711
rect 13111 5739 13127 5753
rect 13111 5705 13112 5739
rect 13161 5719 13199 5753
rect 13284 5735 13367 5769
rect 13401 5735 13417 5769
rect 13451 5735 13467 5769
rect 13501 5739 13526 5769
rect 13146 5705 13199 5719
rect 13451 5705 13480 5735
rect 13514 5705 13526 5739
rect 13585 5710 13818 5767
rect 14239 5761 14273 5799
rect 14341 5831 14359 5865
rect 14307 5794 14359 5831
rect 12928 5625 13008 5663
rect 12928 5591 12974 5625
rect 12928 5535 13008 5591
rect 13043 5573 13077 5695
rect 13165 5641 13204 5671
rect 13165 5607 13199 5641
rect 13238 5637 13249 5671
rect 13585 5657 13619 5710
rect 13233 5607 13249 5637
rect 13295 5641 13552 5657
rect 13329 5623 13552 5641
rect 13586 5623 13619 5657
rect 13664 5671 13736 5673
rect 13698 5657 13736 5671
rect 13664 5623 13669 5637
rect 13703 5623 13736 5657
rect 13329 5607 13345 5623
rect 13664 5607 13736 5623
rect 13784 5641 13818 5710
rect 13852 5739 13930 5754
rect 14128 5745 14194 5761
rect 14128 5739 14160 5745
rect 13886 5738 13930 5739
rect 13886 5705 13896 5738
rect 13852 5704 13896 5705
rect 13852 5688 13930 5704
rect 13968 5705 13992 5739
rect 14026 5705 14042 5739
rect 14162 5705 14194 5711
rect 13968 5641 14002 5705
rect 14160 5695 14194 5705
rect 14239 5745 14290 5761
rect 14239 5711 14256 5745
rect 14239 5695 14290 5711
rect 13784 5607 14002 5641
rect 14070 5637 14116 5671
rect 14036 5634 14116 5637
rect 14239 5635 14273 5695
rect 14324 5663 14359 5794
rect 13295 5604 13345 5607
rect 13043 5539 13176 5573
rect 13295 5570 13302 5604
rect 13336 5570 13345 5604
rect 14036 5600 14082 5634
rect 14036 5584 14116 5600
rect 13295 5569 13345 5570
rect 12928 5501 12974 5535
rect 13142 5535 13176 5539
rect 13426 5539 13628 5573
rect 13142 5517 13359 5535
rect 12928 5467 13008 5501
rect 13042 5471 13058 5505
rect 13092 5471 13108 5505
rect 8795 5370 8847 5407
rect 11088 5403 11117 5437
rect 11151 5403 11209 5437
rect 11243 5403 11301 5437
rect 11335 5403 11393 5437
rect 11427 5403 11485 5437
rect 11519 5403 11577 5437
rect 11611 5403 11669 5437
rect 11703 5403 11761 5437
rect 11795 5403 11853 5437
rect 11887 5403 11945 5437
rect 11979 5403 12037 5437
rect 12071 5403 12129 5437
rect 12163 5403 12221 5437
rect 12255 5403 12313 5437
rect 12347 5403 12405 5437
rect 12439 5403 12497 5437
rect 12531 5403 12560 5437
rect 13042 5433 13108 5471
rect 13142 5483 13325 5517
rect 13142 5467 13359 5483
rect 13426 5522 13460 5539
rect 13594 5522 13628 5539
rect 13426 5467 13460 5488
rect 13494 5471 13510 5505
rect 13544 5471 13560 5505
rect 13494 5433 13560 5471
rect 13769 5539 13984 5573
rect 14155 5571 14273 5635
rect 14307 5622 14359 5663
rect 14341 5598 14359 5622
rect 14155 5547 14189 5571
rect 13769 5522 13816 5539
rect 13594 5467 13628 5488
rect 13662 5475 13678 5509
rect 13712 5475 13728 5509
rect 13662 5433 13728 5475
rect 13769 5488 13782 5522
rect 13950 5522 13984 5539
rect 13769 5467 13816 5488
rect 13850 5471 13866 5505
rect 13900 5471 13916 5505
rect 13850 5433 13916 5471
rect 13950 5467 13984 5488
rect 14034 5522 14189 5547
rect 14307 5562 14312 5588
rect 14352 5562 14359 5598
rect 14068 5488 14189 5522
rect 14034 5467 14189 5488
rect 14223 5513 14273 5530
rect 14257 5479 14273 5513
rect 14223 5433 14273 5479
rect 14307 5528 14359 5562
rect 14341 5494 14359 5528
rect 14307 5467 14359 5494
rect 14798 5861 14878 5905
rect 14927 5901 14993 5939
rect 14927 5867 14943 5901
rect 14977 5867 14993 5901
rect 15027 5889 15229 5905
rect 14798 5827 14844 5861
rect 15027 5855 15195 5889
rect 15027 5833 15061 5855
rect 15195 5837 15229 5855
rect 15296 5884 15330 5905
rect 15364 5901 15430 5939
rect 15364 5867 15380 5901
rect 15414 5867 15430 5901
rect 15464 5884 15498 5905
rect 14798 5794 14878 5827
rect 14913 5799 15061 5833
rect 15296 5833 15330 5850
rect 15532 5892 15598 5939
rect 15532 5858 15548 5892
rect 15582 5858 15598 5892
rect 15652 5884 15686 5905
rect 15464 5833 15498 5850
rect 14798 5659 14864 5794
rect 14913 5757 14947 5799
rect 14898 5741 14947 5757
rect 15154 5769 15166 5803
rect 15200 5769 15253 5803
rect 15296 5799 15498 5833
rect 15720 5901 15786 5939
rect 15720 5867 15736 5901
rect 15770 5867 15786 5901
rect 15820 5884 15854 5905
rect 15652 5833 15686 5850
rect 15820 5833 15854 5850
rect 15652 5799 15854 5833
rect 15904 5884 16024 5905
rect 15938 5850 16024 5884
rect 16077 5897 16143 5939
rect 16077 5863 16093 5897
rect 16127 5863 16143 5897
rect 15904 5829 16024 5850
rect 16177 5861 16229 5905
rect 15904 5803 16143 5829
rect 15904 5769 15906 5803
rect 15940 5795 16143 5803
rect 15940 5769 15952 5795
rect 15154 5765 15253 5769
rect 14932 5707 14947 5741
rect 14898 5691 14947 5707
rect 14981 5735 14997 5749
rect 14981 5701 14982 5735
rect 15031 5715 15069 5749
rect 15154 5731 15237 5765
rect 15271 5731 15287 5765
rect 15321 5731 15337 5765
rect 15371 5735 15396 5765
rect 15016 5701 15069 5715
rect 15321 5701 15350 5731
rect 15384 5701 15396 5735
rect 15455 5706 15688 5763
rect 16109 5757 16143 5795
rect 16211 5827 16229 5861
rect 16177 5790 16229 5827
rect 14798 5621 14878 5659
rect 14798 5587 14844 5621
rect 14798 5531 14878 5587
rect 14913 5569 14947 5691
rect 15035 5637 15074 5667
rect 15035 5603 15069 5637
rect 15108 5633 15119 5667
rect 15455 5653 15489 5706
rect 15103 5603 15119 5633
rect 15165 5637 15422 5653
rect 15199 5619 15422 5637
rect 15456 5619 15489 5653
rect 15534 5667 15606 5669
rect 15568 5653 15606 5667
rect 15534 5619 15539 5633
rect 15573 5619 15606 5653
rect 15199 5603 15215 5619
rect 15534 5603 15606 5619
rect 15654 5637 15688 5706
rect 15722 5735 15800 5750
rect 15998 5741 16064 5757
rect 15998 5735 16030 5741
rect 15756 5734 15800 5735
rect 15756 5701 15766 5734
rect 15722 5700 15766 5701
rect 15722 5684 15800 5700
rect 15838 5701 15862 5735
rect 15896 5701 15912 5735
rect 16032 5701 16064 5707
rect 15838 5637 15872 5701
rect 16030 5691 16064 5701
rect 16109 5741 16160 5757
rect 16109 5707 16126 5741
rect 16109 5691 16160 5707
rect 15654 5603 15872 5637
rect 15940 5633 15986 5667
rect 15906 5630 15986 5633
rect 16109 5631 16143 5691
rect 16194 5659 16229 5790
rect 15165 5600 15215 5603
rect 14913 5535 15046 5569
rect 15165 5566 15172 5600
rect 15206 5566 15215 5600
rect 15906 5596 15952 5630
rect 15906 5580 15986 5596
rect 15165 5565 15215 5566
rect 14798 5497 14844 5531
rect 15012 5531 15046 5535
rect 15296 5535 15498 5569
rect 15012 5513 15229 5531
rect 14798 5463 14878 5497
rect 14912 5467 14928 5501
rect 14962 5467 14978 5501
rect 12904 5399 12933 5433
rect 12967 5399 13025 5433
rect 13059 5399 13117 5433
rect 13151 5399 13209 5433
rect 13243 5399 13301 5433
rect 13335 5399 13393 5433
rect 13427 5399 13485 5433
rect 13519 5399 13577 5433
rect 13611 5399 13669 5433
rect 13703 5399 13761 5433
rect 13795 5399 13853 5433
rect 13887 5399 13945 5433
rect 13979 5399 14037 5433
rect 14071 5399 14129 5433
rect 14163 5399 14221 5433
rect 14255 5399 14313 5433
rect 14347 5399 14376 5433
rect 14912 5429 14978 5467
rect 15012 5479 15195 5513
rect 15012 5463 15229 5479
rect 15296 5518 15330 5535
rect 15464 5518 15498 5535
rect 15296 5463 15330 5484
rect 15364 5467 15380 5501
rect 15414 5467 15430 5501
rect 15364 5429 15430 5467
rect 15639 5535 15854 5569
rect 16025 5567 16143 5631
rect 16177 5618 16229 5659
rect 16211 5600 16229 5618
rect 16025 5543 16059 5567
rect 15639 5518 15686 5535
rect 15464 5463 15498 5484
rect 15532 5471 15548 5505
rect 15582 5471 15598 5505
rect 15532 5429 15598 5471
rect 15639 5484 15652 5518
rect 15820 5518 15854 5535
rect 15639 5463 15686 5484
rect 15720 5467 15736 5501
rect 15770 5467 15786 5501
rect 15720 5429 15786 5467
rect 15820 5463 15854 5484
rect 15904 5518 16059 5543
rect 16177 5564 16182 5584
rect 16216 5564 16229 5600
rect 15938 5484 16059 5518
rect 15904 5463 16059 5484
rect 16093 5509 16143 5526
rect 16127 5475 16143 5509
rect 16093 5429 16143 5475
rect 16177 5524 16229 5564
rect 16211 5490 16229 5524
rect 16177 5463 16229 5490
rect 14774 5395 14803 5429
rect 14837 5395 14895 5429
rect 14929 5395 14987 5429
rect 15021 5395 15079 5429
rect 15113 5395 15171 5429
rect 15205 5395 15263 5429
rect 15297 5395 15355 5429
rect 15389 5395 15447 5429
rect 15481 5395 15539 5429
rect 15573 5395 15631 5429
rect 15665 5395 15723 5429
rect 15757 5395 15815 5429
rect 15849 5395 15907 5429
rect 15941 5395 15999 5429
rect 16033 5395 16091 5429
rect 16125 5395 16183 5429
rect 16217 5395 16246 5429
rect 7416 5201 7496 5239
rect 7416 5167 7462 5201
rect 7416 5111 7496 5167
rect 7531 5149 7565 5271
rect 7653 5217 7692 5247
rect 7653 5183 7687 5217
rect 7726 5213 7737 5247
rect 8073 5233 8107 5286
rect 7721 5183 7737 5213
rect 7783 5217 8040 5233
rect 7817 5199 8040 5217
rect 8074 5199 8107 5233
rect 8152 5247 8224 5249
rect 8186 5233 8224 5247
rect 8152 5199 8157 5213
rect 8191 5199 8224 5233
rect 7817 5183 7833 5199
rect 8152 5183 8224 5199
rect 8272 5217 8306 5286
rect 8340 5315 8418 5330
rect 8616 5321 8682 5337
rect 8616 5315 8648 5321
rect 8374 5314 8418 5315
rect 8374 5281 8384 5314
rect 8340 5280 8384 5281
rect 8340 5264 8418 5280
rect 8456 5281 8480 5315
rect 8514 5281 8530 5315
rect 8650 5281 8682 5287
rect 8456 5217 8490 5281
rect 8648 5271 8682 5281
rect 8727 5321 8778 5337
rect 8727 5287 8744 5321
rect 8727 5271 8778 5287
rect 8272 5183 8490 5217
rect 8558 5213 8604 5247
rect 8524 5210 8604 5213
rect 8727 5211 8761 5271
rect 8812 5239 8847 5370
rect 7783 5180 7833 5183
rect 7531 5115 7664 5149
rect 7783 5146 7790 5180
rect 7824 5146 7833 5180
rect 8524 5176 8570 5210
rect 8524 5160 8604 5176
rect 7783 5145 7833 5146
rect 7416 5077 7462 5111
rect 7630 5111 7664 5115
rect 7914 5115 8116 5149
rect 7630 5093 7847 5111
rect 7416 5043 7496 5077
rect 7530 5047 7546 5081
rect 7580 5047 7596 5081
rect 5522 4979 5551 5013
rect 5585 4979 5643 5013
rect 5677 4979 5735 5013
rect 5769 4979 5827 5013
rect 5861 4979 5919 5013
rect 5953 4979 6011 5013
rect 6045 4979 6103 5013
rect 6137 4979 6195 5013
rect 6229 4979 6287 5013
rect 6321 4979 6379 5013
rect 6413 4979 6471 5013
rect 6505 4979 6563 5013
rect 6597 4979 6655 5013
rect 6689 4979 6747 5013
rect 6781 4979 6839 5013
rect 6873 4979 6931 5013
rect 6965 4979 6994 5013
rect 7530 5009 7596 5047
rect 7630 5059 7813 5093
rect 7630 5043 7847 5059
rect 7914 5098 7948 5115
rect 8082 5098 8116 5115
rect 7914 5043 7948 5064
rect 7982 5047 7998 5081
rect 8032 5047 8048 5081
rect 7982 5009 8048 5047
rect 8257 5115 8472 5149
rect 8643 5147 8761 5211
rect 8795 5198 8847 5239
rect 8829 5180 8847 5198
rect 8643 5123 8677 5147
rect 8257 5098 8304 5115
rect 8082 5043 8116 5064
rect 8150 5051 8166 5085
rect 8200 5051 8216 5085
rect 8150 5009 8216 5051
rect 8257 5064 8270 5098
rect 8438 5098 8472 5115
rect 8257 5043 8304 5064
rect 8338 5047 8354 5081
rect 8388 5047 8404 5081
rect 8338 5009 8404 5047
rect 8438 5043 8472 5064
rect 8522 5098 8677 5123
rect 8795 5144 8800 5164
rect 8834 5144 8847 5180
rect 8556 5064 8677 5098
rect 8522 5043 8677 5064
rect 8711 5089 8761 5106
rect 8745 5055 8761 5089
rect 8711 5009 8761 5055
rect 8795 5104 8847 5144
rect 8829 5070 8847 5104
rect 9246 5077 9275 5111
rect 9309 5077 9367 5111
rect 9401 5077 9459 5111
rect 9493 5077 9551 5111
rect 9585 5077 9643 5111
rect 9677 5077 9735 5111
rect 9769 5077 9827 5111
rect 9861 5077 9919 5111
rect 9953 5077 10011 5111
rect 10045 5077 10103 5111
rect 10137 5077 10195 5111
rect 10229 5077 10287 5111
rect 10321 5077 10379 5111
rect 10413 5077 10471 5111
rect 10505 5077 10563 5111
rect 10597 5077 10655 5111
rect 10689 5077 10718 5111
rect 8795 5043 8847 5070
rect 7392 4975 7421 5009
rect 7455 4975 7513 5009
rect 7547 4975 7605 5009
rect 7639 4975 7697 5009
rect 7731 4975 7789 5009
rect 7823 4975 7881 5009
rect 7915 4975 7973 5009
rect 8007 4975 8065 5009
rect 8099 4975 8157 5009
rect 8191 4975 8249 5009
rect 8283 4975 8341 5009
rect 8375 4975 8433 5009
rect 8467 4975 8525 5009
rect 8559 4975 8617 5009
rect 8651 4975 8709 5009
rect 8743 4975 8801 5009
rect 8835 4975 8864 5009
rect 9270 4999 9350 5043
rect 9399 5039 9465 5077
rect 9399 5005 9415 5039
rect 9449 5005 9465 5039
rect 9499 5027 9701 5043
rect 9270 4965 9316 4999
rect 9499 4993 9667 5027
rect 9499 4971 9533 4993
rect 9667 4975 9701 4993
rect 9768 5022 9802 5043
rect 9836 5039 9902 5077
rect 9836 5005 9852 5039
rect 9886 5005 9902 5039
rect 9936 5022 9970 5043
rect 9270 4932 9350 4965
rect 9385 4937 9533 4971
rect 9768 4971 9802 4988
rect 10004 5030 10070 5077
rect 10004 4996 10020 5030
rect 10054 4996 10070 5030
rect 10124 5022 10158 5043
rect 9936 4971 9970 4988
rect 9270 4797 9336 4932
rect 9385 4895 9419 4937
rect 9370 4879 9419 4895
rect 9626 4907 9638 4941
rect 9672 4907 9725 4941
rect 9768 4937 9970 4971
rect 10192 5039 10258 5077
rect 10192 5005 10208 5039
rect 10242 5005 10258 5039
rect 10292 5022 10326 5043
rect 10124 4971 10158 4988
rect 10292 4971 10326 4988
rect 10124 4937 10326 4971
rect 10376 5022 10496 5043
rect 10410 4988 10496 5022
rect 10549 5035 10615 5077
rect 11116 5073 11145 5107
rect 11179 5073 11237 5107
rect 11271 5073 11329 5107
rect 11363 5073 11421 5107
rect 11455 5073 11513 5107
rect 11547 5073 11605 5107
rect 11639 5073 11697 5107
rect 11731 5073 11789 5107
rect 11823 5073 11881 5107
rect 11915 5073 11973 5107
rect 12007 5073 12065 5107
rect 12099 5073 12157 5107
rect 12191 5073 12249 5107
rect 12283 5073 12341 5107
rect 12375 5073 12433 5107
rect 12467 5073 12525 5107
rect 12559 5073 12588 5107
rect 10549 5001 10565 5035
rect 10599 5001 10615 5035
rect 10376 4967 10496 4988
rect 10649 4999 10701 5043
rect 10376 4941 10615 4967
rect 10376 4907 10378 4941
rect 10412 4933 10615 4941
rect 10412 4907 10424 4933
rect 9626 4903 9725 4907
rect 9404 4845 9419 4879
rect 9370 4829 9419 4845
rect 9453 4873 9469 4887
rect 9453 4839 9454 4873
rect 9503 4853 9541 4887
rect 9626 4869 9709 4903
rect 9743 4869 9759 4903
rect 9793 4869 9809 4903
rect 9843 4873 9868 4903
rect 9488 4839 9541 4853
rect 9793 4839 9822 4869
rect 9856 4839 9868 4873
rect 9927 4844 10160 4901
rect 10581 4895 10615 4933
rect 10683 4965 10701 4999
rect 10649 4928 10701 4965
rect 9270 4759 9350 4797
rect 9270 4725 9316 4759
rect 9270 4669 9350 4725
rect 9385 4707 9419 4829
rect 9507 4775 9546 4805
rect 9507 4741 9541 4775
rect 9580 4771 9591 4805
rect 9927 4791 9961 4844
rect 9575 4741 9591 4771
rect 9637 4775 9894 4791
rect 9671 4757 9894 4775
rect 9928 4757 9961 4791
rect 10006 4805 10078 4807
rect 10040 4791 10078 4805
rect 10006 4757 10011 4771
rect 10045 4757 10078 4791
rect 9671 4741 9687 4757
rect 10006 4741 10078 4757
rect 10126 4775 10160 4844
rect 10194 4873 10272 4888
rect 10470 4879 10536 4895
rect 10470 4873 10502 4879
rect 10228 4872 10272 4873
rect 10228 4839 10238 4872
rect 10194 4838 10238 4839
rect 10194 4822 10272 4838
rect 10310 4839 10334 4873
rect 10368 4839 10384 4873
rect 10504 4839 10536 4845
rect 10310 4775 10344 4839
rect 10502 4829 10536 4839
rect 10581 4879 10632 4895
rect 10581 4845 10598 4879
rect 10581 4829 10632 4845
rect 10126 4741 10344 4775
rect 10412 4771 10458 4805
rect 10378 4768 10458 4771
rect 10581 4769 10615 4829
rect 10666 4797 10701 4928
rect 9637 4740 9687 4741
rect 9385 4673 9518 4707
rect 9637 4706 9646 4740
rect 9680 4706 9687 4740
rect 10378 4734 10424 4768
rect 10378 4718 10458 4734
rect 9637 4703 9687 4706
rect 9270 4635 9316 4669
rect 9484 4669 9518 4673
rect 9768 4673 9970 4707
rect 9484 4651 9701 4669
rect 9270 4601 9350 4635
rect 9384 4605 9400 4639
rect 9434 4605 9450 4639
rect 9384 4567 9450 4605
rect 9484 4617 9667 4651
rect 9484 4601 9701 4617
rect 9768 4656 9802 4673
rect 9936 4656 9970 4673
rect 9768 4601 9802 4622
rect 9836 4605 9852 4639
rect 9886 4605 9902 4639
rect 9836 4567 9902 4605
rect 10111 4673 10326 4707
rect 10497 4705 10615 4769
rect 10649 4756 10701 4797
rect 10683 4732 10701 4756
rect 10497 4681 10531 4705
rect 10111 4656 10158 4673
rect 9936 4601 9970 4622
rect 10004 4609 10020 4643
rect 10054 4609 10070 4643
rect 10004 4567 10070 4609
rect 10111 4622 10124 4656
rect 10292 4656 10326 4673
rect 10111 4601 10158 4622
rect 10192 4605 10208 4639
rect 10242 4605 10258 4639
rect 10192 4567 10258 4605
rect 10292 4601 10326 4622
rect 10376 4656 10531 4681
rect 10649 4696 10654 4722
rect 10694 4696 10701 4732
rect 10410 4622 10531 4656
rect 10376 4601 10531 4622
rect 10565 4647 10615 4664
rect 10599 4613 10615 4647
rect 10565 4567 10615 4613
rect 10649 4662 10701 4696
rect 10683 4628 10701 4662
rect 10649 4601 10701 4628
rect 11140 4995 11220 5039
rect 11269 5035 11335 5073
rect 11269 5001 11285 5035
rect 11319 5001 11335 5035
rect 11369 5023 11571 5039
rect 11140 4961 11186 4995
rect 11369 4989 11537 5023
rect 11369 4967 11403 4989
rect 11537 4971 11571 4989
rect 11638 5018 11672 5039
rect 11706 5035 11772 5073
rect 11706 5001 11722 5035
rect 11756 5001 11772 5035
rect 11806 5018 11840 5039
rect 11140 4928 11220 4961
rect 11255 4933 11403 4967
rect 11638 4967 11672 4984
rect 11874 5026 11940 5073
rect 11874 4992 11890 5026
rect 11924 4992 11940 5026
rect 11994 5018 12028 5039
rect 11806 4967 11840 4984
rect 11140 4793 11206 4928
rect 11255 4891 11289 4933
rect 11240 4875 11289 4891
rect 11496 4903 11508 4937
rect 11542 4903 11595 4937
rect 11638 4933 11840 4967
rect 12062 5035 12128 5073
rect 12062 5001 12078 5035
rect 12112 5001 12128 5035
rect 12162 5018 12196 5039
rect 11994 4967 12028 4984
rect 12162 4967 12196 4984
rect 11994 4933 12196 4967
rect 12246 5018 12366 5039
rect 12280 4984 12366 5018
rect 12419 5031 12485 5073
rect 12932 5069 12961 5103
rect 12995 5069 13053 5103
rect 13087 5069 13145 5103
rect 13179 5069 13237 5103
rect 13271 5069 13329 5103
rect 13363 5069 13421 5103
rect 13455 5069 13513 5103
rect 13547 5069 13605 5103
rect 13639 5069 13697 5103
rect 13731 5069 13789 5103
rect 13823 5069 13881 5103
rect 13915 5069 13973 5103
rect 14007 5069 14065 5103
rect 14099 5069 14157 5103
rect 14191 5069 14249 5103
rect 14283 5069 14341 5103
rect 14375 5069 14404 5103
rect 12419 4997 12435 5031
rect 12469 4997 12485 5031
rect 12246 4963 12366 4984
rect 12519 4995 12571 5039
rect 12246 4937 12485 4963
rect 12246 4903 12248 4937
rect 12282 4929 12485 4937
rect 12282 4903 12294 4929
rect 11496 4899 11595 4903
rect 11274 4841 11289 4875
rect 11240 4825 11289 4841
rect 11323 4869 11339 4883
rect 11323 4835 11324 4869
rect 11373 4849 11411 4883
rect 11496 4865 11579 4899
rect 11613 4865 11629 4899
rect 11663 4865 11679 4899
rect 11713 4869 11738 4899
rect 11358 4835 11411 4849
rect 11663 4835 11692 4865
rect 11726 4835 11738 4869
rect 11797 4840 12030 4897
rect 12451 4891 12485 4929
rect 12553 4961 12571 4995
rect 12519 4924 12571 4961
rect 11140 4755 11220 4793
rect 11140 4721 11186 4755
rect 11140 4665 11220 4721
rect 11255 4703 11289 4825
rect 11377 4771 11416 4801
rect 11377 4737 11411 4771
rect 11450 4767 11461 4801
rect 11797 4787 11831 4840
rect 11445 4737 11461 4767
rect 11507 4771 11764 4787
rect 11541 4753 11764 4771
rect 11798 4753 11831 4787
rect 11876 4801 11948 4803
rect 11910 4787 11948 4801
rect 11876 4753 11881 4767
rect 11915 4753 11948 4787
rect 11541 4737 11557 4753
rect 11876 4737 11948 4753
rect 11996 4771 12030 4840
rect 12064 4869 12142 4884
rect 12340 4875 12406 4891
rect 12340 4869 12372 4875
rect 12098 4868 12142 4869
rect 12098 4835 12108 4868
rect 12064 4834 12108 4835
rect 12064 4818 12142 4834
rect 12180 4835 12204 4869
rect 12238 4835 12254 4869
rect 12374 4835 12406 4841
rect 12180 4771 12214 4835
rect 12372 4825 12406 4835
rect 12451 4875 12502 4891
rect 12451 4841 12468 4875
rect 12451 4825 12502 4841
rect 11996 4737 12214 4771
rect 12282 4767 12328 4801
rect 12248 4764 12328 4767
rect 12451 4765 12485 4825
rect 12536 4793 12571 4924
rect 11507 4734 11557 4737
rect 11255 4669 11388 4703
rect 11507 4700 11514 4734
rect 11548 4700 11557 4734
rect 12248 4730 12294 4764
rect 12248 4714 12328 4730
rect 11507 4699 11557 4700
rect 11140 4631 11186 4665
rect 11354 4665 11388 4669
rect 11638 4669 11840 4703
rect 11354 4647 11571 4665
rect 11140 4597 11220 4631
rect 11254 4601 11270 4635
rect 11304 4601 11320 4635
rect 9246 4533 9275 4567
rect 9309 4533 9367 4567
rect 9401 4533 9459 4567
rect 9493 4533 9551 4567
rect 9585 4533 9643 4567
rect 9677 4533 9735 4567
rect 9769 4533 9827 4567
rect 9861 4533 9919 4567
rect 9953 4533 10011 4567
rect 10045 4533 10103 4567
rect 10137 4533 10195 4567
rect 10229 4533 10287 4567
rect 10321 4533 10379 4567
rect 10413 4533 10471 4567
rect 10505 4533 10563 4567
rect 10597 4533 10655 4567
rect 10689 4533 10718 4567
rect 11254 4563 11320 4601
rect 11354 4613 11537 4647
rect 11354 4597 11571 4613
rect 11638 4652 11672 4669
rect 11806 4652 11840 4669
rect 11638 4597 11672 4618
rect 11706 4601 11722 4635
rect 11756 4601 11772 4635
rect 11706 4563 11772 4601
rect 11981 4669 12196 4703
rect 12367 4701 12485 4765
rect 12519 4752 12571 4793
rect 12553 4718 12571 4752
rect 12367 4677 12401 4701
rect 11981 4652 12028 4669
rect 11806 4597 11840 4618
rect 11874 4605 11890 4639
rect 11924 4605 11940 4639
rect 11874 4563 11940 4605
rect 11981 4618 11994 4652
rect 12162 4652 12196 4669
rect 11981 4597 12028 4618
rect 12062 4601 12078 4635
rect 12112 4601 12128 4635
rect 12062 4563 12128 4601
rect 12162 4597 12196 4618
rect 12246 4652 12401 4677
rect 12519 4684 12530 4718
rect 12564 4684 12571 4718
rect 12280 4618 12401 4652
rect 12246 4597 12401 4618
rect 12435 4643 12485 4660
rect 12469 4609 12485 4643
rect 12435 4563 12485 4609
rect 12519 4658 12571 4684
rect 12553 4624 12571 4658
rect 12519 4597 12571 4624
rect 12956 4991 13036 5035
rect 13085 5031 13151 5069
rect 13085 4997 13101 5031
rect 13135 4997 13151 5031
rect 13185 5019 13387 5035
rect 12956 4957 13002 4991
rect 13185 4985 13353 5019
rect 13185 4963 13219 4985
rect 13353 4967 13387 4985
rect 13454 5014 13488 5035
rect 13522 5031 13588 5069
rect 13522 4997 13538 5031
rect 13572 4997 13588 5031
rect 13622 5014 13656 5035
rect 12956 4924 13036 4957
rect 13071 4929 13219 4963
rect 13454 4963 13488 4980
rect 13690 5022 13756 5069
rect 13690 4988 13706 5022
rect 13740 4988 13756 5022
rect 13810 5014 13844 5035
rect 13622 4963 13656 4980
rect 12956 4789 13022 4924
rect 13071 4887 13105 4929
rect 13056 4871 13105 4887
rect 13312 4899 13324 4933
rect 13358 4899 13411 4933
rect 13454 4929 13656 4963
rect 13878 5031 13944 5069
rect 13878 4997 13894 5031
rect 13928 4997 13944 5031
rect 13978 5014 14012 5035
rect 13810 4963 13844 4980
rect 13978 4963 14012 4980
rect 13810 4929 14012 4963
rect 14062 5014 14182 5035
rect 14096 4980 14182 5014
rect 14235 5027 14301 5069
rect 14802 5065 14831 5099
rect 14865 5065 14923 5099
rect 14957 5065 15015 5099
rect 15049 5065 15107 5099
rect 15141 5065 15199 5099
rect 15233 5065 15291 5099
rect 15325 5065 15383 5099
rect 15417 5065 15475 5099
rect 15509 5065 15567 5099
rect 15601 5065 15659 5099
rect 15693 5065 15751 5099
rect 15785 5065 15843 5099
rect 15877 5065 15935 5099
rect 15969 5065 16027 5099
rect 16061 5065 16119 5099
rect 16153 5065 16211 5099
rect 16245 5065 16274 5099
rect 14235 4993 14251 5027
rect 14285 4993 14301 5027
rect 14062 4959 14182 4980
rect 14335 4991 14387 5035
rect 14062 4933 14301 4959
rect 14062 4899 14064 4933
rect 14098 4925 14301 4933
rect 14098 4899 14110 4925
rect 13312 4895 13411 4899
rect 13090 4837 13105 4871
rect 13056 4821 13105 4837
rect 13139 4865 13155 4879
rect 13139 4831 13140 4865
rect 13189 4845 13227 4879
rect 13312 4861 13395 4895
rect 13429 4861 13445 4895
rect 13479 4861 13495 4895
rect 13529 4865 13554 4895
rect 13174 4831 13227 4845
rect 13479 4831 13508 4861
rect 13542 4831 13554 4865
rect 13613 4836 13846 4893
rect 14267 4887 14301 4925
rect 14369 4957 14387 4991
rect 14335 4920 14387 4957
rect 12956 4751 13036 4789
rect 12956 4717 13002 4751
rect 12956 4661 13036 4717
rect 13071 4699 13105 4821
rect 13193 4767 13232 4797
rect 13193 4733 13227 4767
rect 13266 4763 13277 4797
rect 13613 4783 13647 4836
rect 13261 4733 13277 4763
rect 13323 4767 13580 4783
rect 13357 4749 13580 4767
rect 13614 4749 13647 4783
rect 13692 4797 13764 4799
rect 13726 4783 13764 4797
rect 13692 4749 13697 4763
rect 13731 4749 13764 4783
rect 13357 4733 13373 4749
rect 13692 4733 13764 4749
rect 13812 4767 13846 4836
rect 13880 4865 13958 4880
rect 14156 4871 14222 4887
rect 14156 4865 14188 4871
rect 13914 4864 13958 4865
rect 13914 4831 13924 4864
rect 13880 4830 13924 4831
rect 13880 4814 13958 4830
rect 13996 4831 14020 4865
rect 14054 4831 14070 4865
rect 14190 4831 14222 4837
rect 13996 4767 14030 4831
rect 14188 4821 14222 4831
rect 14267 4871 14318 4887
rect 14267 4837 14284 4871
rect 14267 4821 14318 4837
rect 13812 4733 14030 4767
rect 14098 4763 14144 4797
rect 14064 4760 14144 4763
rect 14267 4761 14301 4821
rect 14352 4789 14387 4920
rect 13323 4730 13373 4733
rect 13071 4665 13204 4699
rect 13323 4696 13330 4730
rect 13364 4696 13373 4730
rect 14064 4726 14110 4760
rect 14064 4710 14144 4726
rect 13323 4695 13373 4696
rect 12956 4627 13002 4661
rect 13170 4661 13204 4665
rect 13454 4665 13656 4699
rect 13170 4643 13387 4661
rect 12956 4593 13036 4627
rect 13070 4597 13086 4631
rect 13120 4597 13136 4631
rect 11116 4529 11145 4563
rect 11179 4529 11237 4563
rect 11271 4529 11329 4563
rect 11363 4529 11421 4563
rect 11455 4529 11513 4563
rect 11547 4529 11605 4563
rect 11639 4529 11697 4563
rect 11731 4529 11789 4563
rect 11823 4529 11881 4563
rect 11915 4529 11973 4563
rect 12007 4529 12065 4563
rect 12099 4529 12157 4563
rect 12191 4529 12249 4563
rect 12283 4529 12341 4563
rect 12375 4529 12433 4563
rect 12467 4529 12525 4563
rect 12559 4529 12588 4563
rect 13070 4559 13136 4597
rect 13170 4609 13353 4643
rect 13170 4593 13387 4609
rect 13454 4648 13488 4665
rect 13622 4648 13656 4665
rect 13454 4593 13488 4614
rect 13522 4597 13538 4631
rect 13572 4597 13588 4631
rect 13522 4559 13588 4597
rect 13797 4665 14012 4699
rect 14183 4697 14301 4761
rect 14335 4748 14387 4789
rect 14369 4724 14387 4748
rect 14183 4673 14217 4697
rect 13797 4648 13844 4665
rect 13622 4593 13656 4614
rect 13690 4601 13706 4635
rect 13740 4601 13756 4635
rect 13690 4559 13756 4601
rect 13797 4614 13810 4648
rect 13978 4648 14012 4665
rect 13797 4593 13844 4614
rect 13878 4597 13894 4631
rect 13928 4597 13944 4631
rect 13878 4559 13944 4597
rect 13978 4593 14012 4614
rect 14062 4648 14217 4673
rect 14335 4688 14340 4714
rect 14380 4688 14387 4724
rect 14096 4614 14217 4648
rect 14062 4593 14217 4614
rect 14251 4639 14301 4656
rect 14285 4605 14301 4639
rect 14251 4559 14301 4605
rect 14335 4654 14387 4688
rect 14369 4620 14387 4654
rect 14335 4593 14387 4620
rect 14826 4987 14906 5031
rect 14955 5027 15021 5065
rect 14955 4993 14971 5027
rect 15005 4993 15021 5027
rect 15055 5015 15257 5031
rect 14826 4953 14872 4987
rect 15055 4981 15223 5015
rect 15055 4959 15089 4981
rect 15223 4963 15257 4981
rect 15324 5010 15358 5031
rect 15392 5027 15458 5065
rect 15392 4993 15408 5027
rect 15442 4993 15458 5027
rect 15492 5010 15526 5031
rect 14826 4920 14906 4953
rect 14941 4925 15089 4959
rect 15324 4959 15358 4976
rect 15560 5018 15626 5065
rect 15560 4984 15576 5018
rect 15610 4984 15626 5018
rect 15680 5010 15714 5031
rect 15492 4959 15526 4976
rect 14826 4785 14892 4920
rect 14941 4883 14975 4925
rect 14926 4867 14975 4883
rect 15182 4895 15194 4929
rect 15228 4895 15281 4929
rect 15324 4925 15526 4959
rect 15748 5027 15814 5065
rect 15748 4993 15764 5027
rect 15798 4993 15814 5027
rect 15848 5010 15882 5031
rect 15680 4959 15714 4976
rect 15848 4959 15882 4976
rect 15680 4925 15882 4959
rect 15932 5010 16052 5031
rect 15966 4976 16052 5010
rect 16105 5023 16171 5065
rect 16105 4989 16121 5023
rect 16155 4989 16171 5023
rect 15932 4955 16052 4976
rect 16205 4987 16257 5031
rect 15932 4929 16171 4955
rect 15932 4895 15934 4929
rect 15968 4921 16171 4929
rect 15968 4895 15980 4921
rect 15182 4891 15281 4895
rect 14960 4833 14975 4867
rect 14926 4817 14975 4833
rect 15009 4861 15025 4875
rect 15009 4827 15010 4861
rect 15059 4841 15097 4875
rect 15182 4857 15265 4891
rect 15299 4857 15315 4891
rect 15349 4857 15365 4891
rect 15399 4861 15424 4891
rect 15044 4827 15097 4841
rect 15349 4827 15378 4857
rect 15412 4827 15424 4861
rect 15483 4832 15716 4889
rect 16137 4883 16171 4921
rect 16239 4953 16257 4987
rect 16205 4916 16257 4953
rect 14826 4747 14906 4785
rect 14826 4713 14872 4747
rect 14826 4657 14906 4713
rect 14941 4695 14975 4817
rect 15063 4763 15102 4793
rect 15063 4729 15097 4763
rect 15136 4759 15147 4793
rect 15483 4779 15517 4832
rect 15131 4729 15147 4759
rect 15193 4763 15450 4779
rect 15227 4745 15450 4763
rect 15484 4745 15517 4779
rect 15562 4793 15634 4795
rect 15596 4779 15634 4793
rect 15562 4745 15567 4759
rect 15601 4745 15634 4779
rect 15227 4729 15243 4745
rect 15562 4729 15634 4745
rect 15682 4763 15716 4832
rect 15750 4861 15828 4876
rect 16026 4867 16092 4883
rect 16026 4861 16058 4867
rect 15784 4860 15828 4861
rect 15784 4827 15794 4860
rect 15750 4826 15794 4827
rect 15750 4810 15828 4826
rect 15866 4827 15890 4861
rect 15924 4827 15940 4861
rect 16060 4827 16092 4833
rect 15866 4763 15900 4827
rect 16058 4817 16092 4827
rect 16137 4867 16188 4883
rect 16137 4833 16154 4867
rect 16137 4817 16188 4833
rect 15682 4729 15900 4763
rect 15968 4759 16014 4793
rect 15934 4756 16014 4759
rect 16137 4757 16171 4817
rect 16222 4785 16257 4916
rect 15193 4726 15243 4729
rect 14941 4661 15074 4695
rect 15193 4692 15200 4726
rect 15234 4692 15243 4726
rect 15934 4722 15980 4756
rect 15934 4706 16014 4722
rect 15193 4691 15243 4692
rect 14826 4623 14872 4657
rect 15040 4657 15074 4661
rect 15324 4661 15526 4695
rect 15040 4639 15257 4657
rect 14826 4589 14906 4623
rect 14940 4593 14956 4627
rect 14990 4593 15006 4627
rect 12932 4525 12961 4559
rect 12995 4525 13053 4559
rect 13087 4525 13145 4559
rect 13179 4525 13237 4559
rect 13271 4525 13329 4559
rect 13363 4525 13421 4559
rect 13455 4525 13513 4559
rect 13547 4525 13605 4559
rect 13639 4525 13697 4559
rect 13731 4525 13789 4559
rect 13823 4525 13881 4559
rect 13915 4525 13973 4559
rect 14007 4525 14065 4559
rect 14099 4525 14157 4559
rect 14191 4525 14249 4559
rect 14283 4525 14341 4559
rect 14375 4525 14404 4559
rect 14940 4555 15006 4593
rect 15040 4605 15223 4639
rect 15040 4589 15257 4605
rect 15324 4644 15358 4661
rect 15492 4644 15526 4661
rect 15324 4589 15358 4610
rect 15392 4593 15408 4627
rect 15442 4593 15458 4627
rect 15392 4555 15458 4593
rect 15667 4661 15882 4695
rect 16053 4693 16171 4757
rect 16205 4744 16257 4785
rect 16239 4726 16257 4744
rect 16053 4669 16087 4693
rect 15667 4644 15714 4661
rect 15492 4589 15526 4610
rect 15560 4597 15576 4631
rect 15610 4597 15626 4631
rect 15560 4555 15626 4597
rect 15667 4610 15680 4644
rect 15848 4644 15882 4661
rect 15667 4589 15714 4610
rect 15748 4593 15764 4627
rect 15798 4593 15814 4627
rect 15748 4555 15814 4593
rect 15848 4589 15882 4610
rect 15932 4644 16087 4669
rect 16205 4690 16210 4710
rect 16244 4690 16257 4726
rect 15966 4610 16087 4644
rect 15932 4589 16087 4610
rect 16121 4635 16171 4652
rect 16155 4601 16171 4635
rect 16121 4555 16171 4601
rect 16205 4650 16257 4690
rect 16239 4616 16257 4650
rect 16205 4589 16257 4616
rect 14802 4521 14831 4555
rect 14865 4521 14923 4555
rect 14957 4521 15015 4555
rect 15049 4521 15107 4555
rect 15141 4521 15199 4555
rect 15233 4521 15291 4555
rect 15325 4521 15383 4555
rect 15417 4521 15475 4555
rect 15509 4521 15567 4555
rect 15601 4521 15659 4555
rect 15693 4521 15751 4555
rect 15785 4521 15843 4555
rect 15877 4521 15935 4555
rect 15969 4521 16027 4555
rect 16061 4521 16119 4555
rect 16153 4521 16211 4555
rect 16245 4521 16274 4555
rect 1806 2271 1835 2305
rect 1869 2271 1927 2305
rect 1961 2271 2019 2305
rect 2053 2271 2111 2305
rect 2145 2271 2203 2305
rect 2237 2271 2295 2305
rect 2329 2271 2387 2305
rect 2421 2271 2479 2305
rect 2513 2271 2571 2305
rect 2605 2271 2663 2305
rect 2697 2271 2755 2305
rect 2789 2271 2847 2305
rect 2881 2271 2939 2305
rect 2973 2271 3031 2305
rect 3065 2271 3123 2305
rect 3157 2271 3215 2305
rect 3249 2271 3278 2305
rect 1830 2193 1910 2237
rect 1959 2233 2025 2271
rect 1959 2199 1975 2233
rect 2009 2199 2025 2233
rect 2059 2221 2261 2237
rect 1830 2159 1876 2193
rect 2059 2187 2227 2221
rect 2059 2165 2093 2187
rect 2227 2169 2261 2187
rect 2328 2216 2362 2237
rect 2396 2233 2462 2271
rect 2396 2199 2412 2233
rect 2446 2199 2462 2233
rect 2496 2216 2530 2237
rect 1830 2126 1910 2159
rect 1945 2131 2093 2165
rect 2328 2165 2362 2182
rect 2564 2224 2630 2271
rect 2564 2190 2580 2224
rect 2614 2190 2630 2224
rect 2684 2216 2718 2237
rect 2496 2165 2530 2182
rect 1830 1991 1896 2126
rect 1945 2089 1979 2131
rect 1930 2073 1979 2089
rect 2186 2101 2198 2135
rect 2232 2101 2285 2135
rect 2328 2131 2530 2165
rect 2752 2233 2818 2271
rect 2752 2199 2768 2233
rect 2802 2199 2818 2233
rect 2852 2216 2886 2237
rect 2684 2165 2718 2182
rect 2852 2165 2886 2182
rect 2684 2131 2886 2165
rect 2936 2216 3056 2237
rect 2970 2182 3056 2216
rect 3109 2229 3175 2271
rect 3676 2267 3705 2301
rect 3739 2267 3797 2301
rect 3831 2267 3889 2301
rect 3923 2267 3981 2301
rect 4015 2267 4073 2301
rect 4107 2267 4165 2301
rect 4199 2267 4257 2301
rect 4291 2267 4349 2301
rect 4383 2267 4441 2301
rect 4475 2267 4533 2301
rect 4567 2267 4625 2301
rect 4659 2267 4717 2301
rect 4751 2267 4809 2301
rect 4843 2267 4901 2301
rect 4935 2267 4993 2301
rect 5027 2267 5085 2301
rect 5119 2267 5148 2301
rect 3109 2195 3125 2229
rect 3159 2195 3175 2229
rect 2936 2161 3056 2182
rect 3209 2193 3261 2237
rect 2936 2135 3175 2161
rect 2936 2101 2938 2135
rect 2972 2127 3175 2135
rect 2972 2101 2984 2127
rect 2186 2097 2285 2101
rect 1964 2039 1979 2073
rect 1930 2023 1979 2039
rect 2013 2067 2029 2081
rect 2013 2033 2014 2067
rect 2063 2047 2101 2081
rect 2186 2063 2269 2097
rect 2303 2063 2319 2097
rect 2353 2063 2369 2097
rect 2403 2067 2428 2097
rect 2048 2033 2101 2047
rect 2353 2033 2382 2063
rect 2416 2033 2428 2067
rect 2487 2038 2720 2095
rect 3141 2089 3175 2127
rect 3243 2159 3261 2193
rect 3209 2122 3261 2159
rect 1830 1953 1910 1991
rect 1830 1919 1876 1953
rect 1830 1863 1910 1919
rect 1945 1901 1979 2023
rect 2067 1969 2106 1999
rect 2067 1935 2101 1969
rect 2140 1965 2151 1999
rect 2487 1985 2521 2038
rect 2135 1935 2151 1965
rect 2197 1969 2454 1985
rect 2231 1951 2454 1969
rect 2488 1951 2521 1985
rect 2566 1999 2638 2001
rect 2600 1985 2638 1999
rect 2566 1951 2571 1965
rect 2605 1951 2638 1985
rect 2231 1935 2247 1951
rect 2566 1935 2638 1951
rect 2686 1969 2720 2038
rect 2754 2067 2832 2082
rect 3030 2073 3096 2089
rect 3030 2067 3062 2073
rect 2788 2066 2832 2067
rect 2788 2033 2798 2066
rect 2754 2032 2798 2033
rect 2754 2016 2832 2032
rect 2870 2033 2894 2067
rect 2928 2033 2944 2067
rect 3064 2033 3096 2039
rect 2870 1969 2904 2033
rect 3062 2023 3096 2033
rect 3141 2073 3192 2089
rect 3141 2039 3158 2073
rect 3141 2023 3192 2039
rect 2686 1935 2904 1969
rect 2972 1965 3018 1999
rect 2938 1962 3018 1965
rect 3141 1963 3175 2023
rect 3226 1991 3261 2122
rect 2197 1934 2247 1935
rect 1945 1867 2078 1901
rect 2197 1900 2206 1934
rect 2240 1900 2247 1934
rect 2938 1928 2984 1962
rect 2938 1912 3018 1928
rect 2197 1897 2247 1900
rect 1830 1829 1876 1863
rect 2044 1863 2078 1867
rect 2328 1867 2530 1901
rect 2044 1845 2261 1863
rect 1830 1795 1910 1829
rect 1944 1799 1960 1833
rect 1994 1799 2010 1833
rect 1944 1761 2010 1799
rect 2044 1811 2227 1845
rect 2044 1795 2261 1811
rect 2328 1850 2362 1867
rect 2496 1850 2530 1867
rect 2328 1795 2362 1816
rect 2396 1799 2412 1833
rect 2446 1799 2462 1833
rect 2396 1761 2462 1799
rect 2671 1867 2886 1901
rect 3057 1899 3175 1963
rect 3209 1950 3261 1991
rect 3243 1926 3261 1950
rect 3057 1875 3091 1899
rect 2671 1850 2718 1867
rect 2496 1795 2530 1816
rect 2564 1803 2580 1837
rect 2614 1803 2630 1837
rect 2564 1761 2630 1803
rect 2671 1816 2684 1850
rect 2852 1850 2886 1867
rect 2671 1795 2718 1816
rect 2752 1799 2768 1833
rect 2802 1799 2818 1833
rect 2752 1761 2818 1799
rect 2852 1795 2886 1816
rect 2936 1850 3091 1875
rect 3209 1890 3214 1916
rect 3254 1890 3261 1926
rect 2970 1816 3091 1850
rect 2936 1795 3091 1816
rect 3125 1841 3175 1858
rect 3159 1807 3175 1841
rect 3125 1761 3175 1807
rect 3209 1856 3261 1890
rect 3243 1822 3261 1856
rect 3209 1795 3261 1822
rect 3700 2189 3780 2233
rect 3829 2229 3895 2267
rect 3829 2195 3845 2229
rect 3879 2195 3895 2229
rect 3929 2217 4131 2233
rect 3700 2155 3746 2189
rect 3929 2183 4097 2217
rect 3929 2161 3963 2183
rect 4097 2165 4131 2183
rect 4198 2212 4232 2233
rect 4266 2229 4332 2267
rect 4266 2195 4282 2229
rect 4316 2195 4332 2229
rect 4366 2212 4400 2233
rect 3700 2122 3780 2155
rect 3815 2127 3963 2161
rect 4198 2161 4232 2178
rect 4434 2220 4500 2267
rect 4434 2186 4450 2220
rect 4484 2186 4500 2220
rect 4554 2212 4588 2233
rect 4366 2161 4400 2178
rect 3700 1987 3766 2122
rect 3815 2085 3849 2127
rect 3800 2069 3849 2085
rect 4056 2097 4068 2131
rect 4102 2097 4155 2131
rect 4198 2127 4400 2161
rect 4622 2229 4688 2267
rect 4622 2195 4638 2229
rect 4672 2195 4688 2229
rect 4722 2212 4756 2233
rect 4554 2161 4588 2178
rect 4722 2161 4756 2178
rect 4554 2127 4756 2161
rect 4806 2212 4926 2233
rect 4840 2178 4926 2212
rect 4979 2225 5045 2267
rect 5492 2263 5521 2297
rect 5555 2263 5613 2297
rect 5647 2263 5705 2297
rect 5739 2263 5797 2297
rect 5831 2263 5889 2297
rect 5923 2263 5981 2297
rect 6015 2263 6073 2297
rect 6107 2263 6165 2297
rect 6199 2263 6257 2297
rect 6291 2263 6349 2297
rect 6383 2263 6441 2297
rect 6475 2263 6533 2297
rect 6567 2263 6625 2297
rect 6659 2263 6717 2297
rect 6751 2263 6809 2297
rect 6843 2263 6901 2297
rect 6935 2263 6964 2297
rect 4979 2191 4995 2225
rect 5029 2191 5045 2225
rect 4806 2157 4926 2178
rect 5079 2189 5131 2233
rect 4806 2131 5045 2157
rect 4806 2097 4808 2131
rect 4842 2123 5045 2131
rect 4842 2097 4854 2123
rect 4056 2093 4155 2097
rect 3834 2035 3849 2069
rect 3800 2019 3849 2035
rect 3883 2063 3899 2077
rect 3883 2029 3884 2063
rect 3933 2043 3971 2077
rect 4056 2059 4139 2093
rect 4173 2059 4189 2093
rect 4223 2059 4239 2093
rect 4273 2063 4298 2093
rect 3918 2029 3971 2043
rect 4223 2029 4252 2059
rect 4286 2029 4298 2063
rect 4357 2034 4590 2091
rect 5011 2085 5045 2123
rect 5113 2155 5131 2189
rect 5079 2118 5131 2155
rect 3700 1949 3780 1987
rect 3700 1915 3746 1949
rect 3700 1859 3780 1915
rect 3815 1897 3849 2019
rect 3937 1965 3976 1995
rect 3937 1931 3971 1965
rect 4010 1961 4021 1995
rect 4357 1981 4391 2034
rect 4005 1931 4021 1961
rect 4067 1965 4324 1981
rect 4101 1947 4324 1965
rect 4358 1947 4391 1981
rect 4436 1995 4508 1997
rect 4470 1981 4508 1995
rect 4436 1947 4441 1961
rect 4475 1947 4508 1981
rect 4101 1931 4117 1947
rect 4436 1931 4508 1947
rect 4556 1965 4590 2034
rect 4624 2063 4702 2078
rect 4900 2069 4966 2085
rect 4900 2063 4932 2069
rect 4658 2062 4702 2063
rect 4658 2029 4668 2062
rect 4624 2028 4668 2029
rect 4624 2012 4702 2028
rect 4740 2029 4764 2063
rect 4798 2029 4814 2063
rect 4934 2029 4966 2035
rect 4740 1965 4774 2029
rect 4932 2019 4966 2029
rect 5011 2069 5062 2085
rect 5011 2035 5028 2069
rect 5011 2019 5062 2035
rect 4556 1931 4774 1965
rect 4842 1961 4888 1995
rect 4808 1958 4888 1961
rect 5011 1959 5045 2019
rect 5096 1987 5131 2118
rect 4067 1928 4117 1931
rect 3815 1863 3948 1897
rect 4067 1894 4074 1928
rect 4108 1894 4117 1928
rect 4808 1924 4854 1958
rect 4808 1908 4888 1924
rect 4067 1893 4117 1894
rect 3700 1825 3746 1859
rect 3914 1859 3948 1863
rect 4198 1863 4400 1897
rect 3914 1841 4131 1859
rect 3700 1791 3780 1825
rect 3814 1795 3830 1829
rect 3864 1795 3880 1829
rect 1806 1727 1835 1761
rect 1869 1727 1927 1761
rect 1961 1727 2019 1761
rect 2053 1727 2111 1761
rect 2145 1727 2203 1761
rect 2237 1727 2295 1761
rect 2329 1727 2387 1761
rect 2421 1727 2479 1761
rect 2513 1727 2571 1761
rect 2605 1727 2663 1761
rect 2697 1727 2755 1761
rect 2789 1727 2847 1761
rect 2881 1727 2939 1761
rect 2973 1727 3031 1761
rect 3065 1727 3123 1761
rect 3157 1727 3215 1761
rect 3249 1727 3278 1761
rect 3814 1757 3880 1795
rect 3914 1807 4097 1841
rect 3914 1791 4131 1807
rect 4198 1846 4232 1863
rect 4366 1846 4400 1863
rect 4198 1791 4232 1812
rect 4266 1795 4282 1829
rect 4316 1795 4332 1829
rect 4266 1757 4332 1795
rect 4541 1863 4756 1897
rect 4927 1895 5045 1959
rect 5079 1946 5131 1987
rect 5113 1922 5131 1946
rect 4927 1871 4961 1895
rect 4541 1846 4588 1863
rect 4366 1791 4400 1812
rect 4434 1799 4450 1833
rect 4484 1799 4500 1833
rect 4434 1757 4500 1799
rect 4541 1812 4554 1846
rect 4722 1846 4756 1863
rect 4541 1791 4588 1812
rect 4622 1795 4638 1829
rect 4672 1795 4688 1829
rect 4622 1757 4688 1795
rect 4722 1791 4756 1812
rect 4806 1846 4961 1871
rect 5079 1886 5090 1912
rect 5124 1886 5131 1922
rect 4840 1812 4961 1846
rect 4806 1791 4961 1812
rect 4995 1837 5045 1854
rect 5029 1803 5045 1837
rect 4995 1757 5045 1803
rect 5079 1852 5131 1886
rect 5113 1818 5131 1852
rect 5079 1791 5131 1818
rect 5516 2185 5596 2229
rect 5645 2225 5711 2263
rect 5645 2191 5661 2225
rect 5695 2191 5711 2225
rect 5745 2213 5947 2229
rect 5516 2151 5562 2185
rect 5745 2179 5913 2213
rect 5745 2157 5779 2179
rect 5913 2161 5947 2179
rect 6014 2208 6048 2229
rect 6082 2225 6148 2263
rect 6082 2191 6098 2225
rect 6132 2191 6148 2225
rect 6182 2208 6216 2229
rect 5516 2118 5596 2151
rect 5631 2123 5779 2157
rect 6014 2157 6048 2174
rect 6250 2216 6316 2263
rect 6250 2182 6266 2216
rect 6300 2182 6316 2216
rect 6370 2208 6404 2229
rect 6182 2157 6216 2174
rect 5516 1983 5582 2118
rect 5631 2081 5665 2123
rect 5616 2065 5665 2081
rect 5872 2093 5884 2127
rect 5918 2093 5971 2127
rect 6014 2123 6216 2157
rect 6438 2225 6504 2263
rect 6438 2191 6454 2225
rect 6488 2191 6504 2225
rect 6538 2208 6572 2229
rect 6370 2157 6404 2174
rect 6538 2157 6572 2174
rect 6370 2123 6572 2157
rect 6622 2208 6742 2229
rect 6656 2174 6742 2208
rect 6795 2221 6861 2263
rect 7362 2259 7391 2293
rect 7425 2259 7483 2293
rect 7517 2259 7575 2293
rect 7609 2259 7667 2293
rect 7701 2259 7759 2293
rect 7793 2259 7851 2293
rect 7885 2259 7943 2293
rect 7977 2259 8035 2293
rect 8069 2259 8127 2293
rect 8161 2259 8219 2293
rect 8253 2259 8311 2293
rect 8345 2259 8403 2293
rect 8437 2259 8495 2293
rect 8529 2259 8587 2293
rect 8621 2259 8679 2293
rect 8713 2259 8771 2293
rect 8805 2259 8834 2293
rect 6795 2187 6811 2221
rect 6845 2187 6861 2221
rect 6622 2153 6742 2174
rect 6895 2185 6947 2229
rect 6622 2127 6861 2153
rect 6622 2093 6624 2127
rect 6658 2119 6861 2127
rect 6658 2093 6670 2119
rect 5872 2089 5971 2093
rect 5650 2031 5665 2065
rect 5616 2015 5665 2031
rect 5699 2059 5715 2073
rect 5699 2025 5700 2059
rect 5749 2039 5787 2073
rect 5872 2055 5955 2089
rect 5989 2055 6005 2089
rect 6039 2055 6055 2089
rect 6089 2059 6114 2089
rect 5734 2025 5787 2039
rect 6039 2025 6068 2055
rect 6102 2025 6114 2059
rect 6173 2030 6406 2087
rect 6827 2081 6861 2119
rect 6929 2151 6947 2185
rect 6895 2114 6947 2151
rect 5516 1945 5596 1983
rect 5516 1911 5562 1945
rect 5516 1855 5596 1911
rect 5631 1893 5665 2015
rect 5753 1961 5792 1991
rect 5753 1927 5787 1961
rect 5826 1957 5837 1991
rect 6173 1977 6207 2030
rect 5821 1927 5837 1957
rect 5883 1961 6140 1977
rect 5917 1943 6140 1961
rect 6174 1943 6207 1977
rect 6252 1991 6324 1993
rect 6286 1977 6324 1991
rect 6252 1943 6257 1957
rect 6291 1943 6324 1977
rect 5917 1927 5933 1943
rect 6252 1927 6324 1943
rect 6372 1961 6406 2030
rect 6440 2059 6518 2074
rect 6716 2065 6782 2081
rect 6716 2059 6748 2065
rect 6474 2058 6518 2059
rect 6474 2025 6484 2058
rect 6440 2024 6484 2025
rect 6440 2008 6518 2024
rect 6556 2025 6580 2059
rect 6614 2025 6630 2059
rect 6750 2025 6782 2031
rect 6556 1961 6590 2025
rect 6748 2015 6782 2025
rect 6827 2065 6878 2081
rect 6827 2031 6844 2065
rect 6827 2015 6878 2031
rect 6372 1927 6590 1961
rect 6658 1957 6704 1991
rect 6624 1954 6704 1957
rect 6827 1955 6861 2015
rect 6912 1983 6947 2114
rect 5883 1924 5933 1927
rect 5631 1859 5764 1893
rect 5883 1890 5890 1924
rect 5924 1890 5933 1924
rect 6624 1920 6670 1954
rect 6624 1904 6704 1920
rect 5883 1889 5933 1890
rect 5516 1821 5562 1855
rect 5730 1855 5764 1859
rect 6014 1859 6216 1893
rect 5730 1837 5947 1855
rect 5516 1787 5596 1821
rect 5630 1791 5646 1825
rect 5680 1791 5696 1825
rect 3676 1723 3705 1757
rect 3739 1723 3797 1757
rect 3831 1723 3889 1757
rect 3923 1723 3981 1757
rect 4015 1723 4073 1757
rect 4107 1723 4165 1757
rect 4199 1723 4257 1757
rect 4291 1723 4349 1757
rect 4383 1723 4441 1757
rect 4475 1723 4533 1757
rect 4567 1723 4625 1757
rect 4659 1723 4717 1757
rect 4751 1723 4809 1757
rect 4843 1723 4901 1757
rect 4935 1723 4993 1757
rect 5027 1723 5085 1757
rect 5119 1723 5148 1757
rect 5630 1753 5696 1791
rect 5730 1803 5913 1837
rect 5730 1787 5947 1803
rect 6014 1842 6048 1859
rect 6182 1842 6216 1859
rect 6014 1787 6048 1808
rect 6082 1791 6098 1825
rect 6132 1791 6148 1825
rect 6082 1753 6148 1791
rect 6357 1859 6572 1893
rect 6743 1891 6861 1955
rect 6895 1942 6947 1983
rect 6929 1918 6947 1942
rect 6743 1867 6777 1891
rect 6357 1842 6404 1859
rect 6182 1787 6216 1808
rect 6250 1795 6266 1829
rect 6300 1795 6316 1829
rect 6250 1753 6316 1795
rect 6357 1808 6370 1842
rect 6538 1842 6572 1859
rect 6357 1787 6404 1808
rect 6438 1791 6454 1825
rect 6488 1791 6504 1825
rect 6438 1753 6504 1791
rect 6538 1787 6572 1808
rect 6622 1842 6777 1867
rect 6895 1882 6900 1908
rect 6940 1882 6947 1918
rect 6656 1808 6777 1842
rect 6622 1787 6777 1808
rect 6811 1833 6861 1850
rect 6845 1799 6861 1833
rect 6811 1753 6861 1799
rect 6895 1848 6947 1882
rect 6929 1814 6947 1848
rect 6895 1787 6947 1814
rect 7386 2181 7466 2225
rect 7515 2221 7581 2259
rect 7515 2187 7531 2221
rect 7565 2187 7581 2221
rect 7615 2209 7817 2225
rect 7386 2147 7432 2181
rect 7615 2175 7783 2209
rect 7615 2153 7649 2175
rect 7783 2157 7817 2175
rect 7884 2204 7918 2225
rect 7952 2221 8018 2259
rect 7952 2187 7968 2221
rect 8002 2187 8018 2221
rect 8052 2204 8086 2225
rect 7386 2114 7466 2147
rect 7501 2119 7649 2153
rect 7884 2153 7918 2170
rect 8120 2212 8186 2259
rect 8120 2178 8136 2212
rect 8170 2178 8186 2212
rect 8240 2204 8274 2225
rect 8052 2153 8086 2170
rect 7386 1979 7452 2114
rect 7501 2077 7535 2119
rect 7486 2061 7535 2077
rect 7742 2089 7754 2123
rect 7788 2089 7841 2123
rect 7884 2119 8086 2153
rect 8308 2221 8374 2259
rect 8308 2187 8324 2221
rect 8358 2187 8374 2221
rect 8408 2204 8442 2225
rect 8240 2153 8274 2170
rect 8408 2153 8442 2170
rect 8240 2119 8442 2153
rect 8492 2204 8612 2225
rect 8526 2170 8612 2204
rect 8665 2217 8731 2259
rect 9176 2257 9205 2291
rect 9239 2257 9297 2291
rect 9331 2257 9389 2291
rect 9423 2257 9481 2291
rect 9515 2257 9573 2291
rect 9607 2257 9665 2291
rect 9699 2257 9757 2291
rect 9791 2257 9849 2291
rect 9883 2257 9941 2291
rect 9975 2257 10033 2291
rect 10067 2257 10125 2291
rect 10159 2257 10217 2291
rect 10251 2257 10309 2291
rect 10343 2257 10401 2291
rect 10435 2257 10493 2291
rect 10527 2257 10585 2291
rect 10619 2257 10648 2291
rect 8665 2183 8681 2217
rect 8715 2183 8731 2217
rect 8492 2149 8612 2170
rect 8765 2181 8817 2225
rect 8492 2123 8731 2149
rect 8492 2089 8494 2123
rect 8528 2115 8731 2123
rect 8528 2089 8540 2115
rect 7742 2085 7841 2089
rect 7520 2027 7535 2061
rect 7486 2011 7535 2027
rect 7569 2055 7585 2069
rect 7569 2021 7570 2055
rect 7619 2035 7657 2069
rect 7742 2051 7825 2085
rect 7859 2051 7875 2085
rect 7909 2051 7925 2085
rect 7959 2055 7984 2085
rect 7604 2021 7657 2035
rect 7909 2021 7938 2051
rect 7972 2021 7984 2055
rect 8043 2026 8276 2083
rect 8697 2077 8731 2115
rect 8799 2147 8817 2181
rect 8765 2110 8817 2147
rect 7386 1941 7466 1979
rect 7386 1907 7432 1941
rect 7386 1851 7466 1907
rect 7501 1889 7535 2011
rect 7623 1957 7662 1987
rect 7623 1923 7657 1957
rect 7696 1953 7707 1987
rect 8043 1973 8077 2026
rect 7691 1923 7707 1953
rect 7753 1957 8010 1973
rect 7787 1939 8010 1957
rect 8044 1939 8077 1973
rect 8122 1987 8194 1989
rect 8156 1973 8194 1987
rect 8122 1939 8127 1953
rect 8161 1939 8194 1973
rect 7787 1923 7803 1939
rect 8122 1923 8194 1939
rect 8242 1957 8276 2026
rect 8310 2055 8388 2070
rect 8586 2061 8652 2077
rect 8586 2055 8618 2061
rect 8344 2054 8388 2055
rect 8344 2021 8354 2054
rect 8310 2020 8354 2021
rect 8310 2004 8388 2020
rect 8426 2021 8450 2055
rect 8484 2021 8500 2055
rect 8620 2021 8652 2027
rect 8426 1957 8460 2021
rect 8618 2011 8652 2021
rect 8697 2061 8748 2077
rect 8697 2027 8714 2061
rect 8697 2011 8748 2027
rect 8242 1923 8460 1957
rect 8528 1953 8574 1987
rect 8494 1950 8574 1953
rect 8697 1951 8731 2011
rect 8782 1979 8817 2110
rect 7753 1920 7803 1923
rect 7501 1855 7634 1889
rect 7753 1886 7760 1920
rect 7794 1886 7803 1920
rect 8494 1916 8540 1950
rect 8494 1900 8574 1916
rect 7753 1885 7803 1886
rect 7386 1817 7432 1851
rect 7600 1851 7634 1855
rect 7884 1855 8086 1889
rect 7600 1833 7817 1851
rect 7386 1783 7466 1817
rect 7500 1787 7516 1821
rect 7550 1787 7566 1821
rect 5492 1719 5521 1753
rect 5555 1719 5613 1753
rect 5647 1719 5705 1753
rect 5739 1719 5797 1753
rect 5831 1719 5889 1753
rect 5923 1719 5981 1753
rect 6015 1719 6073 1753
rect 6107 1719 6165 1753
rect 6199 1719 6257 1753
rect 6291 1719 6349 1753
rect 6383 1719 6441 1753
rect 6475 1719 6533 1753
rect 6567 1719 6625 1753
rect 6659 1719 6717 1753
rect 6751 1719 6809 1753
rect 6843 1719 6901 1753
rect 6935 1719 6964 1753
rect 7500 1749 7566 1787
rect 7600 1799 7783 1833
rect 7600 1783 7817 1799
rect 7884 1838 7918 1855
rect 8052 1838 8086 1855
rect 7884 1783 7918 1804
rect 7952 1787 7968 1821
rect 8002 1787 8018 1821
rect 7952 1749 8018 1787
rect 8227 1855 8442 1889
rect 8613 1887 8731 1951
rect 8765 1938 8817 1979
rect 8799 1920 8817 1938
rect 8613 1863 8647 1887
rect 8227 1838 8274 1855
rect 8052 1783 8086 1804
rect 8120 1791 8136 1825
rect 8170 1791 8186 1825
rect 8120 1749 8186 1791
rect 8227 1804 8240 1838
rect 8408 1838 8442 1855
rect 8227 1783 8274 1804
rect 8308 1787 8324 1821
rect 8358 1787 8374 1821
rect 8308 1749 8374 1787
rect 8408 1783 8442 1804
rect 8492 1838 8647 1863
rect 8765 1884 8770 1904
rect 8804 1884 8817 1920
rect 8526 1804 8647 1838
rect 8492 1783 8647 1804
rect 8681 1829 8731 1846
rect 8715 1795 8731 1829
rect 8681 1749 8731 1795
rect 8765 1844 8817 1884
rect 8799 1810 8817 1844
rect 8765 1783 8817 1810
rect 9200 2179 9280 2223
rect 9329 2219 9395 2257
rect 9329 2185 9345 2219
rect 9379 2185 9395 2219
rect 9429 2207 9631 2223
rect 9200 2145 9246 2179
rect 9429 2173 9597 2207
rect 9429 2151 9463 2173
rect 9597 2155 9631 2173
rect 9698 2202 9732 2223
rect 9766 2219 9832 2257
rect 9766 2185 9782 2219
rect 9816 2185 9832 2219
rect 9866 2202 9900 2223
rect 9200 2112 9280 2145
rect 9315 2117 9463 2151
rect 9698 2151 9732 2168
rect 9934 2210 10000 2257
rect 9934 2176 9950 2210
rect 9984 2176 10000 2210
rect 10054 2202 10088 2223
rect 9866 2151 9900 2168
rect 9200 1977 9266 2112
rect 9315 2075 9349 2117
rect 9300 2059 9349 2075
rect 9556 2087 9568 2121
rect 9602 2087 9655 2121
rect 9698 2117 9900 2151
rect 10122 2219 10188 2257
rect 10122 2185 10138 2219
rect 10172 2185 10188 2219
rect 10222 2202 10256 2223
rect 10054 2151 10088 2168
rect 10222 2151 10256 2168
rect 10054 2117 10256 2151
rect 10306 2202 10426 2223
rect 10340 2168 10426 2202
rect 10479 2215 10545 2257
rect 11046 2253 11075 2287
rect 11109 2253 11167 2287
rect 11201 2253 11259 2287
rect 11293 2253 11351 2287
rect 11385 2253 11443 2287
rect 11477 2253 11535 2287
rect 11569 2253 11627 2287
rect 11661 2253 11719 2287
rect 11753 2253 11811 2287
rect 11845 2253 11903 2287
rect 11937 2253 11995 2287
rect 12029 2253 12087 2287
rect 12121 2253 12179 2287
rect 12213 2253 12271 2287
rect 12305 2253 12363 2287
rect 12397 2253 12455 2287
rect 12489 2253 12518 2287
rect 10479 2181 10495 2215
rect 10529 2181 10545 2215
rect 10306 2147 10426 2168
rect 10579 2179 10631 2223
rect 10306 2121 10545 2147
rect 10306 2087 10308 2121
rect 10342 2113 10545 2121
rect 10342 2087 10354 2113
rect 9556 2083 9655 2087
rect 9334 2025 9349 2059
rect 9300 2009 9349 2025
rect 9383 2053 9399 2067
rect 9383 2019 9384 2053
rect 9433 2033 9471 2067
rect 9556 2049 9639 2083
rect 9673 2049 9689 2083
rect 9723 2049 9739 2083
rect 9773 2053 9798 2083
rect 9418 2019 9471 2033
rect 9723 2019 9752 2049
rect 9786 2019 9798 2053
rect 9857 2024 10090 2081
rect 10511 2075 10545 2113
rect 10613 2145 10631 2179
rect 10579 2108 10631 2145
rect 9200 1939 9280 1977
rect 9200 1905 9246 1939
rect 9200 1849 9280 1905
rect 9315 1887 9349 2009
rect 9437 1955 9476 1985
rect 9437 1921 9471 1955
rect 9510 1951 9521 1985
rect 9857 1971 9891 2024
rect 9505 1921 9521 1951
rect 9567 1955 9824 1971
rect 9601 1937 9824 1955
rect 9858 1937 9891 1971
rect 9936 1985 10008 1987
rect 9970 1971 10008 1985
rect 9936 1937 9941 1951
rect 9975 1937 10008 1971
rect 9601 1921 9617 1937
rect 9936 1921 10008 1937
rect 10056 1955 10090 2024
rect 10124 2053 10202 2068
rect 10400 2059 10466 2075
rect 10400 2053 10432 2059
rect 10158 2052 10202 2053
rect 10158 2019 10168 2052
rect 10124 2018 10168 2019
rect 10124 2002 10202 2018
rect 10240 2019 10264 2053
rect 10298 2019 10314 2053
rect 10434 2019 10466 2025
rect 10240 1955 10274 2019
rect 10432 2009 10466 2019
rect 10511 2059 10562 2075
rect 10511 2025 10528 2059
rect 10511 2009 10562 2025
rect 10056 1921 10274 1955
rect 10342 1951 10388 1985
rect 10308 1948 10388 1951
rect 10511 1949 10545 2009
rect 10596 1977 10631 2108
rect 9567 1918 9617 1921
rect 9315 1853 9448 1887
rect 9567 1884 9574 1918
rect 9610 1884 9617 1918
rect 10308 1914 10354 1948
rect 10308 1898 10388 1914
rect 9567 1883 9617 1884
rect 9200 1815 9246 1849
rect 9414 1849 9448 1853
rect 9698 1853 9900 1887
rect 9414 1831 9631 1849
rect 9200 1781 9280 1815
rect 9314 1785 9330 1819
rect 9364 1785 9380 1819
rect 7362 1715 7391 1749
rect 7425 1715 7483 1749
rect 7517 1715 7575 1749
rect 7609 1715 7667 1749
rect 7701 1715 7759 1749
rect 7793 1715 7851 1749
rect 7885 1715 7943 1749
rect 7977 1715 8035 1749
rect 8069 1715 8127 1749
rect 8161 1715 8219 1749
rect 8253 1715 8311 1749
rect 8345 1715 8403 1749
rect 8437 1715 8495 1749
rect 8529 1715 8587 1749
rect 8621 1715 8679 1749
rect 8713 1715 8771 1749
rect 8805 1715 8834 1749
rect 9314 1747 9380 1785
rect 9414 1797 9597 1831
rect 9414 1781 9631 1797
rect 9698 1836 9732 1853
rect 9866 1836 9900 1853
rect 9698 1781 9732 1802
rect 9766 1785 9782 1819
rect 9816 1785 9832 1819
rect 9766 1747 9832 1785
rect 10041 1853 10256 1887
rect 10427 1885 10545 1949
rect 10579 1936 10631 1977
rect 10613 1912 10631 1936
rect 10427 1861 10461 1885
rect 10041 1836 10088 1853
rect 9866 1781 9900 1802
rect 9934 1789 9950 1823
rect 9984 1789 10000 1823
rect 9934 1747 10000 1789
rect 10041 1802 10054 1836
rect 10222 1836 10256 1853
rect 10041 1781 10088 1802
rect 10122 1785 10138 1819
rect 10172 1785 10188 1819
rect 10122 1747 10188 1785
rect 10222 1781 10256 1802
rect 10306 1836 10461 1861
rect 10579 1876 10584 1902
rect 10624 1876 10631 1912
rect 10340 1802 10461 1836
rect 10306 1781 10461 1802
rect 10495 1827 10545 1844
rect 10529 1793 10545 1827
rect 10495 1747 10545 1793
rect 10579 1842 10631 1876
rect 10613 1808 10631 1842
rect 10579 1781 10631 1808
rect 11070 2175 11150 2219
rect 11199 2215 11265 2253
rect 11199 2181 11215 2215
rect 11249 2181 11265 2215
rect 11299 2203 11501 2219
rect 11070 2141 11116 2175
rect 11299 2169 11467 2203
rect 11299 2147 11333 2169
rect 11467 2151 11501 2169
rect 11568 2198 11602 2219
rect 11636 2215 11702 2253
rect 11636 2181 11652 2215
rect 11686 2181 11702 2215
rect 11736 2198 11770 2219
rect 11070 2108 11150 2141
rect 11185 2113 11333 2147
rect 11568 2147 11602 2164
rect 11804 2206 11870 2253
rect 11804 2172 11820 2206
rect 11854 2172 11870 2206
rect 11924 2198 11958 2219
rect 11736 2147 11770 2164
rect 11070 1973 11136 2108
rect 11185 2071 11219 2113
rect 11170 2055 11219 2071
rect 11426 2083 11438 2117
rect 11472 2083 11525 2117
rect 11568 2113 11770 2147
rect 11992 2215 12058 2253
rect 11992 2181 12008 2215
rect 12042 2181 12058 2215
rect 12092 2198 12126 2219
rect 11924 2147 11958 2164
rect 12092 2147 12126 2164
rect 11924 2113 12126 2147
rect 12176 2198 12296 2219
rect 12210 2164 12296 2198
rect 12349 2211 12415 2253
rect 12862 2249 12891 2283
rect 12925 2249 12983 2283
rect 13017 2249 13075 2283
rect 13109 2249 13167 2283
rect 13201 2249 13259 2283
rect 13293 2249 13351 2283
rect 13385 2249 13443 2283
rect 13477 2249 13535 2283
rect 13569 2249 13627 2283
rect 13661 2249 13719 2283
rect 13753 2249 13811 2283
rect 13845 2249 13903 2283
rect 13937 2249 13995 2283
rect 14029 2249 14087 2283
rect 14121 2249 14179 2283
rect 14213 2249 14271 2283
rect 14305 2249 14334 2283
rect 12349 2177 12365 2211
rect 12399 2177 12415 2211
rect 12176 2143 12296 2164
rect 12449 2175 12501 2219
rect 12176 2117 12415 2143
rect 12176 2083 12178 2117
rect 12212 2109 12415 2117
rect 12212 2083 12224 2109
rect 11426 2079 11525 2083
rect 11204 2021 11219 2055
rect 11170 2005 11219 2021
rect 11253 2049 11269 2063
rect 11253 2015 11254 2049
rect 11303 2029 11341 2063
rect 11426 2045 11509 2079
rect 11543 2045 11559 2079
rect 11593 2045 11609 2079
rect 11643 2049 11668 2079
rect 11288 2015 11341 2029
rect 11593 2015 11622 2045
rect 11656 2015 11668 2049
rect 11727 2020 11960 2077
rect 12381 2071 12415 2109
rect 12483 2141 12501 2175
rect 12449 2104 12501 2141
rect 11070 1935 11150 1973
rect 11070 1901 11116 1935
rect 11070 1845 11150 1901
rect 11185 1883 11219 2005
rect 11307 1951 11346 1981
rect 11307 1917 11341 1951
rect 11380 1947 11391 1981
rect 11727 1967 11761 2020
rect 11375 1917 11391 1947
rect 11437 1951 11694 1967
rect 11471 1933 11694 1951
rect 11728 1933 11761 1967
rect 11806 1981 11878 1983
rect 11840 1967 11878 1981
rect 11806 1933 11811 1947
rect 11845 1933 11878 1967
rect 11471 1917 11487 1933
rect 11806 1917 11878 1933
rect 11926 1951 11960 2020
rect 11994 2049 12072 2064
rect 12270 2055 12336 2071
rect 12270 2049 12302 2055
rect 12028 2048 12072 2049
rect 12028 2015 12038 2048
rect 11994 2014 12038 2015
rect 11994 1998 12072 2014
rect 12110 2015 12134 2049
rect 12168 2015 12184 2049
rect 12304 2015 12336 2021
rect 12110 1951 12144 2015
rect 12302 2005 12336 2015
rect 12381 2055 12432 2071
rect 12381 2021 12398 2055
rect 12381 2005 12432 2021
rect 11926 1917 12144 1951
rect 12212 1947 12258 1981
rect 12178 1944 12258 1947
rect 12381 1945 12415 2005
rect 12466 1973 12501 2104
rect 11437 1914 11487 1917
rect 11185 1849 11318 1883
rect 11437 1880 11444 1914
rect 11478 1880 11487 1914
rect 12178 1910 12224 1944
rect 12178 1894 12258 1910
rect 11437 1879 11487 1880
rect 11070 1811 11116 1845
rect 11284 1845 11318 1849
rect 11568 1849 11770 1883
rect 11284 1827 11501 1845
rect 11070 1777 11150 1811
rect 11184 1781 11200 1815
rect 11234 1781 11250 1815
rect 9176 1713 9205 1747
rect 9239 1713 9297 1747
rect 9331 1713 9389 1747
rect 9423 1713 9481 1747
rect 9515 1713 9573 1747
rect 9607 1713 9665 1747
rect 9699 1713 9757 1747
rect 9791 1713 9849 1747
rect 9883 1713 9941 1747
rect 9975 1713 10033 1747
rect 10067 1713 10125 1747
rect 10159 1713 10217 1747
rect 10251 1713 10309 1747
rect 10343 1713 10401 1747
rect 10435 1713 10493 1747
rect 10527 1713 10585 1747
rect 10619 1713 10648 1747
rect 11184 1743 11250 1781
rect 11284 1793 11467 1827
rect 11284 1777 11501 1793
rect 11568 1832 11602 1849
rect 11736 1832 11770 1849
rect 11568 1777 11602 1798
rect 11636 1781 11652 1815
rect 11686 1781 11702 1815
rect 11636 1743 11702 1781
rect 11911 1849 12126 1883
rect 12297 1881 12415 1945
rect 12449 1932 12501 1973
rect 12483 1912 12501 1932
rect 12297 1857 12331 1881
rect 11911 1832 11958 1849
rect 11736 1777 11770 1798
rect 11804 1785 11820 1819
rect 11854 1785 11870 1819
rect 11804 1743 11870 1785
rect 11911 1798 11924 1832
rect 12092 1832 12126 1849
rect 11911 1777 11958 1798
rect 11992 1781 12008 1815
rect 12042 1781 12058 1815
rect 11992 1743 12058 1781
rect 12092 1777 12126 1798
rect 12176 1832 12331 1857
rect 12449 1878 12454 1898
rect 12488 1878 12501 1912
rect 12210 1798 12331 1832
rect 12176 1777 12331 1798
rect 12365 1823 12415 1840
rect 12399 1789 12415 1823
rect 12365 1743 12415 1789
rect 12449 1838 12501 1878
rect 12483 1804 12501 1838
rect 12449 1777 12501 1804
rect 12886 2171 12966 2215
rect 13015 2211 13081 2249
rect 13015 2177 13031 2211
rect 13065 2177 13081 2211
rect 13115 2199 13317 2215
rect 12886 2137 12932 2171
rect 13115 2165 13283 2199
rect 13115 2143 13149 2165
rect 13283 2147 13317 2165
rect 13384 2194 13418 2215
rect 13452 2211 13518 2249
rect 13452 2177 13468 2211
rect 13502 2177 13518 2211
rect 13552 2194 13586 2215
rect 12886 2104 12966 2137
rect 13001 2109 13149 2143
rect 13384 2143 13418 2160
rect 13620 2202 13686 2249
rect 13620 2168 13636 2202
rect 13670 2168 13686 2202
rect 13740 2194 13774 2215
rect 13552 2143 13586 2160
rect 12886 1969 12952 2104
rect 13001 2067 13035 2109
rect 12986 2051 13035 2067
rect 13242 2079 13254 2113
rect 13288 2079 13341 2113
rect 13384 2109 13586 2143
rect 13808 2211 13874 2249
rect 13808 2177 13824 2211
rect 13858 2177 13874 2211
rect 13908 2194 13942 2215
rect 13740 2143 13774 2160
rect 13908 2143 13942 2160
rect 13740 2109 13942 2143
rect 13992 2194 14112 2215
rect 14026 2160 14112 2194
rect 14165 2207 14231 2249
rect 14732 2245 14761 2279
rect 14795 2245 14853 2279
rect 14887 2245 14945 2279
rect 14979 2245 15037 2279
rect 15071 2245 15129 2279
rect 15163 2245 15221 2279
rect 15255 2245 15313 2279
rect 15347 2245 15405 2279
rect 15439 2245 15497 2279
rect 15531 2245 15589 2279
rect 15623 2245 15681 2279
rect 15715 2245 15773 2279
rect 15807 2245 15865 2279
rect 15899 2245 15957 2279
rect 15991 2245 16049 2279
rect 16083 2245 16141 2279
rect 16175 2245 16204 2279
rect 14165 2173 14181 2207
rect 14215 2173 14231 2207
rect 13992 2139 14112 2160
rect 14265 2171 14317 2215
rect 13992 2113 14231 2139
rect 13992 2079 13994 2113
rect 14028 2105 14231 2113
rect 14028 2079 14040 2105
rect 13242 2075 13341 2079
rect 13020 2017 13035 2051
rect 12986 2001 13035 2017
rect 13069 2045 13085 2059
rect 13069 2011 13070 2045
rect 13119 2025 13157 2059
rect 13242 2041 13325 2075
rect 13359 2041 13375 2075
rect 13409 2041 13425 2075
rect 13459 2045 13484 2075
rect 13104 2011 13157 2025
rect 13409 2011 13438 2041
rect 13472 2011 13484 2045
rect 13543 2016 13776 2073
rect 14197 2067 14231 2105
rect 14299 2137 14317 2171
rect 14265 2100 14317 2137
rect 12886 1931 12966 1969
rect 12886 1897 12932 1931
rect 12886 1841 12966 1897
rect 13001 1879 13035 2001
rect 13123 1947 13162 1977
rect 13123 1913 13157 1947
rect 13196 1943 13207 1977
rect 13543 1963 13577 2016
rect 13191 1913 13207 1943
rect 13253 1947 13510 1963
rect 13287 1929 13510 1947
rect 13544 1929 13577 1963
rect 13622 1977 13694 1979
rect 13656 1963 13694 1977
rect 13622 1929 13627 1943
rect 13661 1929 13694 1963
rect 13287 1913 13303 1929
rect 13622 1913 13694 1929
rect 13742 1947 13776 2016
rect 13810 2045 13888 2060
rect 14086 2051 14152 2067
rect 14086 2045 14118 2051
rect 13844 2044 13888 2045
rect 13844 2011 13854 2044
rect 13810 2010 13854 2011
rect 13810 1994 13888 2010
rect 13926 2011 13950 2045
rect 13984 2011 14000 2045
rect 14120 2011 14152 2017
rect 13926 1947 13960 2011
rect 14118 2001 14152 2011
rect 14197 2051 14248 2067
rect 14197 2017 14214 2051
rect 14197 2001 14248 2017
rect 13742 1913 13960 1947
rect 14028 1943 14074 1977
rect 13994 1940 14074 1943
rect 14197 1941 14231 2001
rect 14282 1969 14317 2100
rect 13253 1910 13303 1913
rect 13001 1845 13134 1879
rect 13253 1876 13260 1910
rect 13294 1876 13303 1910
rect 13994 1906 14040 1940
rect 13994 1890 14074 1906
rect 13253 1875 13303 1876
rect 12886 1807 12932 1841
rect 13100 1841 13134 1845
rect 13384 1845 13586 1879
rect 13100 1823 13317 1841
rect 12886 1773 12966 1807
rect 13000 1777 13016 1811
rect 13050 1777 13066 1811
rect 11046 1709 11075 1743
rect 11109 1709 11167 1743
rect 11201 1709 11259 1743
rect 11293 1709 11351 1743
rect 11385 1709 11443 1743
rect 11477 1709 11535 1743
rect 11569 1709 11627 1743
rect 11661 1709 11719 1743
rect 11753 1709 11811 1743
rect 11845 1709 11903 1743
rect 11937 1709 11995 1743
rect 12029 1709 12087 1743
rect 12121 1709 12179 1743
rect 12213 1709 12271 1743
rect 12305 1709 12363 1743
rect 12397 1709 12455 1743
rect 12489 1709 12518 1743
rect 13000 1739 13066 1777
rect 13100 1789 13283 1823
rect 13100 1773 13317 1789
rect 13384 1828 13418 1845
rect 13552 1828 13586 1845
rect 13384 1773 13418 1794
rect 13452 1777 13468 1811
rect 13502 1777 13518 1811
rect 13452 1739 13518 1777
rect 13727 1845 13942 1879
rect 14113 1877 14231 1941
rect 14265 1928 14317 1969
rect 14299 1904 14317 1928
rect 14113 1853 14147 1877
rect 13727 1828 13774 1845
rect 13552 1773 13586 1794
rect 13620 1781 13636 1815
rect 13670 1781 13686 1815
rect 13620 1739 13686 1781
rect 13727 1794 13740 1828
rect 13908 1828 13942 1845
rect 13727 1773 13774 1794
rect 13808 1777 13824 1811
rect 13858 1777 13874 1811
rect 13808 1739 13874 1777
rect 13908 1773 13942 1794
rect 13992 1828 14147 1853
rect 14265 1868 14270 1894
rect 14310 1868 14317 1904
rect 14026 1794 14147 1828
rect 13992 1773 14147 1794
rect 14181 1819 14231 1836
rect 14215 1785 14231 1819
rect 14181 1739 14231 1785
rect 14265 1834 14317 1868
rect 14299 1800 14317 1834
rect 14265 1773 14317 1800
rect 14756 2167 14836 2211
rect 14885 2207 14951 2245
rect 14885 2173 14901 2207
rect 14935 2173 14951 2207
rect 14985 2195 15187 2211
rect 14756 2133 14802 2167
rect 14985 2161 15153 2195
rect 14985 2139 15019 2161
rect 15153 2143 15187 2161
rect 15254 2190 15288 2211
rect 15322 2207 15388 2245
rect 15322 2173 15338 2207
rect 15372 2173 15388 2207
rect 15422 2190 15456 2211
rect 14756 2100 14836 2133
rect 14871 2105 15019 2139
rect 15254 2139 15288 2156
rect 15490 2198 15556 2245
rect 15490 2164 15506 2198
rect 15540 2164 15556 2198
rect 15610 2190 15644 2211
rect 15422 2139 15456 2156
rect 14756 1965 14822 2100
rect 14871 2063 14905 2105
rect 14856 2047 14905 2063
rect 15112 2075 15124 2109
rect 15158 2075 15211 2109
rect 15254 2105 15456 2139
rect 15678 2207 15744 2245
rect 15678 2173 15694 2207
rect 15728 2173 15744 2207
rect 15778 2190 15812 2211
rect 15610 2139 15644 2156
rect 15778 2139 15812 2156
rect 15610 2105 15812 2139
rect 15862 2190 15982 2211
rect 15896 2156 15982 2190
rect 16035 2203 16101 2245
rect 16035 2169 16051 2203
rect 16085 2169 16101 2203
rect 15862 2135 15982 2156
rect 16135 2167 16187 2211
rect 15862 2109 16101 2135
rect 15862 2075 15864 2109
rect 15898 2101 16101 2109
rect 15898 2075 15910 2101
rect 15112 2071 15211 2075
rect 14890 2013 14905 2047
rect 14856 1997 14905 2013
rect 14939 2041 14955 2055
rect 14939 2007 14940 2041
rect 14989 2021 15027 2055
rect 15112 2037 15195 2071
rect 15229 2037 15245 2071
rect 15279 2037 15295 2071
rect 15329 2041 15354 2071
rect 14974 2007 15027 2021
rect 15279 2007 15308 2037
rect 15342 2007 15354 2041
rect 15413 2012 15646 2069
rect 16067 2063 16101 2101
rect 16169 2133 16187 2167
rect 16135 2096 16187 2133
rect 14756 1927 14836 1965
rect 14756 1893 14802 1927
rect 14756 1837 14836 1893
rect 14871 1875 14905 1997
rect 14993 1943 15032 1973
rect 14993 1909 15027 1943
rect 15066 1939 15077 1973
rect 15413 1959 15447 2012
rect 15061 1909 15077 1939
rect 15123 1943 15380 1959
rect 15157 1925 15380 1943
rect 15414 1925 15447 1959
rect 15492 1973 15564 1975
rect 15526 1959 15564 1973
rect 15492 1925 15497 1939
rect 15531 1925 15564 1959
rect 15157 1909 15173 1925
rect 15492 1909 15564 1925
rect 15612 1943 15646 2012
rect 15680 2041 15758 2056
rect 15956 2047 16022 2063
rect 15956 2041 15988 2047
rect 15714 2040 15758 2041
rect 15714 2007 15724 2040
rect 15680 2006 15724 2007
rect 15680 1990 15758 2006
rect 15796 2007 15820 2041
rect 15854 2007 15870 2041
rect 15990 2007 16022 2013
rect 15796 1943 15830 2007
rect 15988 1997 16022 2007
rect 16067 2047 16118 2063
rect 16067 2013 16084 2047
rect 16067 1997 16118 2013
rect 15612 1909 15830 1943
rect 15898 1939 15944 1973
rect 15864 1936 15944 1939
rect 16067 1937 16101 1997
rect 16152 1965 16187 2096
rect 15123 1906 15173 1909
rect 14871 1841 15004 1875
rect 15123 1872 15130 1906
rect 15164 1872 15173 1906
rect 15864 1902 15910 1936
rect 15864 1886 15944 1902
rect 15123 1871 15173 1872
rect 14756 1803 14802 1837
rect 14970 1837 15004 1841
rect 15254 1841 15456 1875
rect 14970 1819 15187 1837
rect 14756 1769 14836 1803
rect 14870 1773 14886 1807
rect 14920 1773 14936 1807
rect 12862 1705 12891 1739
rect 12925 1705 12983 1739
rect 13017 1705 13075 1739
rect 13109 1705 13167 1739
rect 13201 1705 13259 1739
rect 13293 1705 13351 1739
rect 13385 1705 13443 1739
rect 13477 1705 13535 1739
rect 13569 1705 13627 1739
rect 13661 1705 13719 1739
rect 13753 1705 13811 1739
rect 13845 1705 13903 1739
rect 13937 1705 13995 1739
rect 14029 1705 14087 1739
rect 14121 1705 14179 1739
rect 14213 1705 14271 1739
rect 14305 1705 14334 1739
rect 14870 1735 14936 1773
rect 14970 1785 15153 1819
rect 14970 1769 15187 1785
rect 15254 1824 15288 1841
rect 15422 1824 15456 1841
rect 15254 1769 15288 1790
rect 15322 1773 15338 1807
rect 15372 1773 15388 1807
rect 15322 1735 15388 1773
rect 15597 1841 15812 1875
rect 15983 1873 16101 1937
rect 16135 1924 16187 1965
rect 16169 1918 16187 1924
rect 16135 1884 16150 1890
rect 16186 1884 16187 1918
rect 15983 1849 16017 1873
rect 15597 1824 15644 1841
rect 15422 1769 15456 1790
rect 15490 1777 15506 1811
rect 15540 1777 15556 1811
rect 15490 1735 15556 1777
rect 15597 1790 15610 1824
rect 15778 1824 15812 1841
rect 15597 1769 15644 1790
rect 15678 1773 15694 1807
rect 15728 1773 15744 1807
rect 15678 1735 15744 1773
rect 15778 1769 15812 1790
rect 15862 1824 16017 1849
rect 15896 1790 16017 1824
rect 15862 1769 16017 1790
rect 16051 1815 16101 1832
rect 16085 1781 16101 1815
rect 16051 1735 16101 1781
rect 16135 1830 16187 1884
rect 16169 1796 16187 1830
rect 16135 1769 16187 1796
rect 14732 1701 14761 1735
rect 14795 1701 14853 1735
rect 14887 1701 14945 1735
rect 14979 1701 15037 1735
rect 15071 1701 15129 1735
rect 15163 1701 15221 1735
rect 15255 1701 15313 1735
rect 15347 1701 15405 1735
rect 15439 1701 15497 1735
rect 15531 1701 15589 1735
rect 15623 1701 15681 1735
rect 15715 1701 15773 1735
rect 15807 1701 15865 1735
rect 15899 1701 15957 1735
rect 15991 1701 16049 1735
rect 16083 1701 16141 1735
rect 16175 1701 16204 1735
<< viali >>
rect 9496 17532 9532 17568
rect 9596 17536 9632 17572
rect 9459 16553 9493 16587
rect 9551 16553 9585 16587
rect 9643 16553 9677 16587
rect 9735 16553 9769 16587
rect 9827 16553 9861 16587
rect 9919 16553 9953 16587
rect 10011 16553 10045 16587
rect 10006 16367 10040 16374
rect 10006 16336 10031 16367
rect 10031 16336 10040 16367
rect 16416 16366 16452 16400
rect 16502 16354 16540 16388
rect 17184 16358 17222 16392
rect 17278 16350 17312 16384
rect 18048 16362 18082 16396
rect 18150 16358 18186 16392
rect 18672 16356 18708 16390
rect 18758 16344 18796 16378
rect 19440 16348 19478 16382
rect 19534 16340 19568 16374
rect 20304 16352 20338 16386
rect 20406 16348 20442 16382
rect 21436 16350 21472 16384
rect 21522 16338 21560 16372
rect 22204 16342 22242 16376
rect 22298 16334 22332 16368
rect 23068 16346 23102 16380
rect 23170 16342 23206 16376
rect 9516 16275 9550 16276
rect 9516 16242 9549 16275
rect 9549 16242 9550 16275
rect 9636 16275 9670 16278
rect 9636 16244 9666 16275
rect 9666 16244 9670 16275
rect 9459 16009 9493 16043
rect 9551 16009 9585 16043
rect 9643 16009 9677 16043
rect 9735 16009 9769 16043
rect 9827 16009 9861 16043
rect 9919 16009 9953 16043
rect 10011 16009 10045 16043
rect 9557 15809 9591 15843
rect 9649 15809 9683 15843
rect 9741 15809 9775 15843
rect 9833 15809 9867 15843
rect 9925 15809 9959 15843
rect 11599 15699 11633 15733
rect 11691 15699 11725 15733
rect 11783 15699 11817 15733
rect 11875 15699 11909 15733
rect 11967 15699 12001 15733
rect 12059 15699 12093 15733
rect 12151 15699 12185 15733
rect 9550 15514 9592 15554
rect 9740 15531 9782 15544
rect 9740 15504 9743 15531
rect 9743 15504 9777 15531
rect 9777 15504 9782 15531
rect 9932 15440 9968 15474
rect 11594 15348 11630 15384
rect 9557 15265 9591 15299
rect 9649 15265 9683 15299
rect 9741 15265 9775 15299
rect 9833 15265 9867 15299
rect 9925 15265 9959 15299
rect 11766 15387 11781 15418
rect 11781 15387 11800 15418
rect 11766 15382 11800 15387
rect 11864 15260 11898 15294
rect 11960 15328 11994 15364
rect 12152 15382 12186 15416
rect 10741 15199 10775 15233
rect 10833 15199 10867 15233
rect 10925 15199 10959 15233
rect 11017 15199 11051 15233
rect 11109 15199 11143 15233
rect 9469 14989 9503 15023
rect 9561 14989 9595 15023
rect 9653 14989 9687 15023
rect 9745 14989 9779 15023
rect 9837 14989 9871 15023
rect 9929 14989 9963 15023
rect 10021 14989 10055 15023
rect 11599 15155 11633 15189
rect 11691 15155 11725 15189
rect 11783 15155 11817 15189
rect 11875 15155 11909 15189
rect 11967 15155 12001 15189
rect 12059 15155 12093 15189
rect 12151 15155 12185 15189
rect 11106 15123 11113 15132
rect 11113 15123 11146 15132
rect 11106 15096 11146 15123
rect 10018 14905 10041 14914
rect 10041 14905 10052 14914
rect 10018 14880 10052 14905
rect 10786 14921 10820 14922
rect 10786 14888 10820 14921
rect 10926 14921 10962 14922
rect 10926 14888 10927 14921
rect 10927 14888 10961 14921
rect 10961 14888 10962 14921
rect 9526 14711 9560 14712
rect 9526 14678 9559 14711
rect 9559 14678 9560 14711
rect 9646 14711 9680 14714
rect 9646 14680 9676 14711
rect 9676 14680 9680 14711
rect 10741 14655 10775 14689
rect 10833 14655 10867 14689
rect 10925 14655 10959 14689
rect 11017 14655 11051 14689
rect 11109 14655 11143 14689
rect 24150 14616 24186 14650
rect 23530 14546 23568 14580
rect 23672 14528 23708 14562
rect 24556 14554 24592 14588
rect 25364 14562 25400 14598
rect 24456 14518 24492 14552
rect 24712 14528 24746 14562
rect 9469 14445 9503 14479
rect 9561 14445 9595 14479
rect 9653 14445 9687 14479
rect 9745 14445 9779 14479
rect 9837 14445 9871 14479
rect 9929 14445 9963 14479
rect 10021 14445 10055 14479
rect 9567 14245 9601 14279
rect 9659 14245 9693 14279
rect 9751 14245 9785 14279
rect 9843 14245 9877 14279
rect 9935 14245 9969 14279
rect 10815 14233 10849 14267
rect 10907 14233 10941 14267
rect 10999 14233 11033 14267
rect 11091 14233 11125 14267
rect 11183 14233 11217 14267
rect 11275 14233 11309 14267
rect 11367 14233 11401 14267
rect 8130 14032 8172 14072
rect 9560 13950 9602 13990
rect 7674 13914 7714 13948
rect 9750 13967 9792 13980
rect 9750 13940 9753 13967
rect 9753 13940 9787 13967
rect 9787 13940 9792 13967
rect 9940 13834 9976 13868
rect 12633 14217 12667 14251
rect 12725 14217 12759 14251
rect 12817 14217 12851 14251
rect 12909 14217 12943 14251
rect 13001 14217 13035 14251
rect 13093 14217 13127 14251
rect 12778 14116 12814 14150
rect 10812 13955 10846 13960
rect 10812 13926 10817 13955
rect 10817 13926 10846 13955
rect 10982 13830 11016 13864
rect 11080 13870 11114 13904
rect 11174 13921 11199 13954
rect 11199 13921 11210 13954
rect 11174 13916 11210 13921
rect 13092 14042 13119 14056
rect 13119 14042 13134 14056
rect 12636 13905 12639 13932
rect 12639 13905 12673 13932
rect 12673 13905 12676 13932
rect 12636 13898 12676 13905
rect 11356 13833 11361 13836
rect 11361 13833 11394 13836
rect 11785 13859 11819 13893
rect 11877 13859 11911 13893
rect 11969 13859 12003 13893
rect 12061 13859 12095 13893
rect 12153 13859 12187 13893
rect 11356 13799 11394 13833
rect 11356 13798 11361 13799
rect 11361 13798 11394 13799
rect 13092 14016 13134 14042
rect 12762 13939 12812 13944
rect 12762 13905 12765 13939
rect 12765 13905 12799 13939
rect 12799 13905 12812 13939
rect 12762 13902 12812 13905
rect 12934 13939 12972 13940
rect 12934 13905 12941 13939
rect 12941 13905 12972 13939
rect 12934 13904 12972 13905
rect 9567 13701 9601 13735
rect 9659 13701 9693 13735
rect 9751 13701 9785 13735
rect 9843 13701 9877 13735
rect 9935 13701 9969 13735
rect 10815 13689 10849 13723
rect 10907 13689 10941 13723
rect 10999 13689 11033 13723
rect 11091 13689 11125 13723
rect 11183 13689 11217 13723
rect 11275 13689 11309 13723
rect 11367 13689 11401 13723
rect 12124 13715 12135 13748
rect 12135 13715 12158 13748
rect 12124 13714 12158 13715
rect 11796 13504 11830 13538
rect 11974 13581 12008 13588
rect 11974 13554 11992 13581
rect 11992 13554 12008 13581
rect 12633 13673 12667 13707
rect 12725 13673 12759 13707
rect 12817 13673 12851 13707
rect 12909 13673 12943 13707
rect 13001 13673 13035 13707
rect 13093 13673 13127 13707
rect 10939 13391 10973 13425
rect 11031 13391 11065 13425
rect 11123 13391 11157 13425
rect 11215 13391 11249 13425
rect 11307 13391 11341 13425
rect 9461 13321 9495 13355
rect 9553 13321 9587 13355
rect 9645 13321 9679 13355
rect 9737 13321 9771 13355
rect 9829 13321 9863 13355
rect 9921 13321 9955 13355
rect 10013 13321 10047 13355
rect 11108 13306 11117 13318
rect 11117 13306 11144 13318
rect 11108 13282 11144 13306
rect 11785 13315 11819 13349
rect 11877 13315 11911 13349
rect 11969 13315 12003 13349
rect 12061 13315 12095 13349
rect 12153 13315 12187 13349
rect 10010 13203 10044 13204
rect 10010 13170 10033 13203
rect 10033 13170 10044 13203
rect 11304 13233 11335 13262
rect 11335 13233 11342 13262
rect 11304 13224 11342 13233
rect 9518 13043 9552 13044
rect 9518 13010 9551 13043
rect 9551 13010 9552 13043
rect 9638 13043 9672 13046
rect 9638 13012 9668 13043
rect 9668 13012 9672 13043
rect 10956 13033 10979 13044
rect 10979 13033 10990 13044
rect 10956 13010 10990 13033
rect 11158 13016 11194 13050
rect 10939 12847 10973 12881
rect 11031 12847 11065 12881
rect 11123 12847 11157 12881
rect 11215 12847 11249 12881
rect 11307 12847 11341 12881
rect 9461 12777 9495 12811
rect 9553 12777 9587 12811
rect 9645 12777 9679 12811
rect 9737 12777 9771 12811
rect 9829 12777 9863 12811
rect 9921 12777 9955 12811
rect 10013 12777 10047 12811
rect 9559 12577 9593 12611
rect 9651 12577 9685 12611
rect 9743 12577 9777 12611
rect 9835 12577 9869 12611
rect 9927 12577 9961 12611
rect 9552 12282 9594 12322
rect 10935 12371 10969 12405
rect 11027 12371 11061 12405
rect 11119 12371 11153 12405
rect 11211 12371 11245 12405
rect 11303 12371 11337 12405
rect 9932 12320 9968 12354
rect 9742 12299 9784 12312
rect 9742 12272 9745 12299
rect 9745 12272 9779 12299
rect 9779 12272 9784 12299
rect 11308 12146 11342 12180
rect 9559 12033 9593 12067
rect 9651 12033 9685 12067
rect 9743 12033 9777 12067
rect 9835 12033 9869 12067
rect 9927 12033 9961 12067
rect 10980 12093 11016 12096
rect 10980 12062 11014 12093
rect 11014 12062 11016 12093
rect 11120 12093 11156 12094
rect 11120 12060 11121 12093
rect 11121 12060 11155 12093
rect 11155 12060 11156 12093
rect 10935 11827 10969 11861
rect 11027 11827 11061 11861
rect 11119 11827 11153 11861
rect 11211 11827 11245 11861
rect 11303 11827 11337 11861
rect 9471 11757 9505 11791
rect 9563 11757 9597 11791
rect 9655 11757 9689 11791
rect 9747 11757 9781 11791
rect 9839 11757 9873 11791
rect 9931 11757 9965 11791
rect 10023 11757 10057 11791
rect 10010 11639 10046 11640
rect 10010 11606 10043 11639
rect 10043 11606 10046 11639
rect 9528 11479 9562 11480
rect 9528 11446 9561 11479
rect 9561 11446 9562 11479
rect 9648 11479 9682 11482
rect 9648 11448 9678 11479
rect 9678 11448 9682 11479
rect 9471 11213 9505 11247
rect 9563 11213 9597 11247
rect 9655 11213 9689 11247
rect 9747 11213 9781 11247
rect 9839 11213 9873 11247
rect 9931 11213 9965 11247
rect 10023 11213 10057 11247
rect 9569 11013 9603 11047
rect 9661 11013 9695 11047
rect 9753 11013 9787 11047
rect 9845 11013 9879 11047
rect 9937 11013 9971 11047
rect 4982 10694 5016 10730
rect 9562 10718 9604 10758
rect 9752 10735 9794 10748
rect 9752 10708 9755 10735
rect 9755 10708 9789 10735
rect 9789 10708 9794 10735
rect 9944 10678 9978 10714
rect 9569 10469 9603 10503
rect 9661 10469 9695 10503
rect 9753 10469 9787 10503
rect 9845 10469 9879 10503
rect 9937 10469 9971 10503
rect 6141 6583 6175 6617
rect 6233 6583 6267 6617
rect 6325 6583 6359 6617
rect 6178 6348 6212 6382
rect 6274 6351 6308 6384
rect 6274 6350 6308 6351
rect 6141 6039 6175 6073
rect 6233 6039 6267 6073
rect 6325 6039 6359 6073
rect 9247 5951 9281 5985
rect 9339 5951 9373 5985
rect 9431 5951 9465 5985
rect 9523 5951 9557 5985
rect 9615 5951 9649 5985
rect 9707 5951 9741 5985
rect 9799 5951 9833 5985
rect 9891 5951 9925 5985
rect 9983 5951 10017 5985
rect 10075 5951 10109 5985
rect 10167 5951 10201 5985
rect 10259 5951 10293 5985
rect 10351 5951 10385 5985
rect 10443 5951 10477 5985
rect 10535 5951 10569 5985
rect 10627 5951 10661 5985
rect 9610 5781 9644 5815
rect 11117 5947 11151 5981
rect 11209 5947 11243 5981
rect 11301 5947 11335 5981
rect 11393 5947 11427 5981
rect 11485 5947 11519 5981
rect 11577 5947 11611 5981
rect 11669 5947 11703 5981
rect 11761 5947 11795 5981
rect 11853 5947 11887 5981
rect 11945 5947 11979 5981
rect 12037 5947 12071 5981
rect 12129 5947 12163 5981
rect 12221 5947 12255 5981
rect 12313 5947 12347 5981
rect 12405 5947 12439 5981
rect 12497 5947 12531 5981
rect 10350 5781 10384 5815
rect 9426 5727 9441 5747
rect 9441 5727 9460 5747
rect 9794 5743 9815 5747
rect 9815 5743 9828 5747
rect 9426 5713 9460 5727
rect 9794 5713 9828 5743
rect 1865 5531 1899 5565
rect 1957 5531 1991 5565
rect 2049 5531 2083 5565
rect 2141 5531 2175 5565
rect 2233 5531 2267 5565
rect 2325 5531 2359 5565
rect 2417 5531 2451 5565
rect 2509 5531 2543 5565
rect 2601 5531 2635 5565
rect 2693 5531 2727 5565
rect 2785 5531 2819 5565
rect 2877 5531 2911 5565
rect 2969 5531 3003 5565
rect 3061 5531 3095 5565
rect 3153 5531 3187 5565
rect 3245 5531 3279 5565
rect 2228 5361 2262 5395
rect 3735 5527 3769 5561
rect 3827 5527 3861 5561
rect 3919 5527 3953 5561
rect 4011 5527 4045 5561
rect 4103 5527 4137 5561
rect 4195 5527 4229 5561
rect 4287 5527 4321 5561
rect 4379 5527 4413 5561
rect 4471 5527 4505 5561
rect 4563 5527 4597 5561
rect 4655 5527 4689 5561
rect 4747 5527 4781 5561
rect 4839 5527 4873 5561
rect 4931 5527 4965 5561
rect 5023 5527 5057 5561
rect 5115 5527 5149 5561
rect 2968 5361 3002 5395
rect 2044 5307 2059 5327
rect 2059 5307 2078 5327
rect 2412 5323 2433 5327
rect 2433 5323 2446 5327
rect 2044 5293 2078 5307
rect 2412 5293 2446 5323
rect 2136 5229 2170 5259
rect 2136 5225 2165 5229
rect 2165 5225 2170 5229
rect 2596 5245 2630 5259
rect 2596 5225 2601 5245
rect 2601 5225 2630 5245
rect 2784 5293 2818 5327
rect 3060 5299 3092 5327
rect 3092 5299 3094 5327
rect 3060 5293 3094 5299
rect 2968 5225 3002 5259
rect 2236 5160 2270 5194
rect 3244 5176 3273 5186
rect 3273 5176 3284 5186
rect 3244 5150 3284 5176
rect 4098 5357 4132 5391
rect 5551 5523 5585 5557
rect 5643 5523 5677 5557
rect 5735 5523 5769 5557
rect 5827 5523 5861 5557
rect 5919 5523 5953 5557
rect 6011 5523 6045 5557
rect 6103 5523 6137 5557
rect 6195 5523 6229 5557
rect 6287 5523 6321 5557
rect 6379 5523 6413 5557
rect 6471 5523 6505 5557
rect 6563 5523 6597 5557
rect 6655 5523 6689 5557
rect 6747 5523 6781 5557
rect 6839 5523 6873 5557
rect 6931 5523 6965 5557
rect 4838 5357 4872 5391
rect 3914 5303 3929 5323
rect 3929 5303 3948 5323
rect 4282 5319 4303 5323
rect 4303 5319 4316 5323
rect 3914 5289 3948 5303
rect 4282 5289 4316 5319
rect 4006 5225 4040 5255
rect 4006 5221 4035 5225
rect 4035 5221 4040 5225
rect 4466 5241 4500 5255
rect 4466 5221 4471 5241
rect 4471 5221 4500 5241
rect 4654 5289 4688 5323
rect 4930 5295 4962 5323
rect 4962 5295 4964 5323
rect 4930 5289 4964 5295
rect 4838 5221 4872 5255
rect 4104 5154 4138 5188
rect 1865 4987 1899 5021
rect 1957 4987 1991 5021
rect 2049 4987 2083 5021
rect 2141 4987 2175 5021
rect 2233 4987 2267 5021
rect 2325 4987 2359 5021
rect 2417 4987 2451 5021
rect 2509 4987 2543 5021
rect 2601 4987 2635 5021
rect 2693 4987 2727 5021
rect 2785 4987 2819 5021
rect 2877 4987 2911 5021
rect 2969 4987 3003 5021
rect 3061 4987 3095 5021
rect 3153 4987 3187 5021
rect 3245 4987 3279 5021
rect 5120 5172 5143 5182
rect 5143 5172 5156 5182
rect 5120 5144 5156 5172
rect 5914 5353 5948 5387
rect 7421 5519 7455 5553
rect 7513 5519 7547 5553
rect 7605 5519 7639 5553
rect 7697 5519 7731 5553
rect 7789 5519 7823 5553
rect 7881 5519 7915 5553
rect 7973 5519 8007 5553
rect 8065 5519 8099 5553
rect 8157 5519 8191 5553
rect 8249 5519 8283 5553
rect 8341 5519 8375 5553
rect 8433 5519 8467 5553
rect 8525 5519 8559 5553
rect 8617 5519 8651 5553
rect 8709 5519 8743 5553
rect 8801 5519 8835 5553
rect 9518 5649 9552 5679
rect 9518 5645 9547 5649
rect 9547 5645 9552 5649
rect 9978 5665 10012 5679
rect 9978 5645 9983 5665
rect 9983 5645 10012 5665
rect 10166 5713 10200 5747
rect 10442 5719 10474 5747
rect 10474 5719 10476 5747
rect 10442 5713 10476 5719
rect 10350 5645 10384 5679
rect 9618 5580 9652 5614
rect 6654 5353 6688 5387
rect 5730 5299 5745 5319
rect 5745 5299 5764 5319
rect 6098 5315 6119 5319
rect 6119 5315 6132 5319
rect 5730 5285 5764 5299
rect 6098 5285 6132 5315
rect 5822 5221 5856 5251
rect 5822 5217 5851 5221
rect 5851 5217 5856 5221
rect 6282 5237 6316 5251
rect 6282 5217 6287 5237
rect 6287 5217 6316 5237
rect 6470 5285 6504 5319
rect 6746 5291 6778 5319
rect 6778 5291 6780 5319
rect 6746 5285 6780 5291
rect 6654 5217 6688 5251
rect 5920 5150 5954 5184
rect 3735 4983 3769 5017
rect 3827 4983 3861 5017
rect 3919 4983 3953 5017
rect 4011 4983 4045 5017
rect 4103 4983 4137 5017
rect 4195 4983 4229 5017
rect 4287 4983 4321 5017
rect 4379 4983 4413 5017
rect 4471 4983 4505 5017
rect 4563 4983 4597 5017
rect 4655 4983 4689 5017
rect 4747 4983 4781 5017
rect 4839 4983 4873 5017
rect 4931 4983 4965 5017
rect 5023 4983 5057 5017
rect 5115 4983 5149 5017
rect 6930 5168 6959 5178
rect 6959 5168 6970 5178
rect 6930 5142 6970 5168
rect 7784 5349 7818 5383
rect 10626 5596 10655 5606
rect 10655 5596 10666 5606
rect 10626 5570 10666 5596
rect 11480 5777 11514 5811
rect 12933 5943 12967 5977
rect 13025 5943 13059 5977
rect 13117 5943 13151 5977
rect 13209 5943 13243 5977
rect 13301 5943 13335 5977
rect 13393 5943 13427 5977
rect 13485 5943 13519 5977
rect 13577 5943 13611 5977
rect 13669 5943 13703 5977
rect 13761 5943 13795 5977
rect 13853 5943 13887 5977
rect 13945 5943 13979 5977
rect 14037 5943 14071 5977
rect 14129 5943 14163 5977
rect 14221 5943 14255 5977
rect 14313 5943 14347 5977
rect 12220 5777 12254 5811
rect 11296 5723 11311 5743
rect 11311 5723 11330 5743
rect 11664 5739 11685 5743
rect 11685 5739 11698 5743
rect 11296 5709 11330 5723
rect 11664 5709 11698 5739
rect 11388 5645 11422 5675
rect 11388 5641 11417 5645
rect 11417 5641 11422 5645
rect 11848 5661 11882 5675
rect 11848 5641 11853 5661
rect 11853 5641 11882 5661
rect 12036 5709 12070 5743
rect 12312 5715 12344 5743
rect 12344 5715 12346 5743
rect 12312 5709 12346 5715
rect 12220 5641 12254 5675
rect 11486 5574 11520 5608
rect 8524 5349 8558 5383
rect 7600 5295 7615 5315
rect 7615 5295 7634 5315
rect 7968 5311 7989 5315
rect 7989 5311 8002 5315
rect 7600 5281 7634 5295
rect 7968 5281 8002 5311
rect 9247 5407 9281 5441
rect 9339 5407 9373 5441
rect 9431 5407 9465 5441
rect 9523 5407 9557 5441
rect 9615 5407 9649 5441
rect 9707 5407 9741 5441
rect 9799 5407 9833 5441
rect 9891 5407 9925 5441
rect 9983 5407 10017 5441
rect 10075 5407 10109 5441
rect 10167 5407 10201 5441
rect 10259 5407 10293 5441
rect 10351 5407 10385 5441
rect 10443 5407 10477 5441
rect 10535 5407 10569 5441
rect 10627 5407 10661 5441
rect 12502 5592 12525 5602
rect 12525 5592 12538 5602
rect 12502 5568 12538 5592
rect 13296 5773 13330 5807
rect 14803 5939 14837 5973
rect 14895 5939 14929 5973
rect 14987 5939 15021 5973
rect 15079 5939 15113 5973
rect 15171 5939 15205 5973
rect 15263 5939 15297 5973
rect 15355 5939 15389 5973
rect 15447 5939 15481 5973
rect 15539 5939 15573 5973
rect 15631 5939 15665 5973
rect 15723 5939 15757 5973
rect 15815 5939 15849 5973
rect 15907 5939 15941 5973
rect 15999 5939 16033 5973
rect 16091 5939 16125 5973
rect 16183 5939 16217 5973
rect 14036 5773 14070 5807
rect 13112 5719 13127 5739
rect 13127 5719 13146 5739
rect 13480 5735 13501 5739
rect 13501 5735 13514 5739
rect 13112 5705 13146 5719
rect 13480 5705 13514 5735
rect 13204 5641 13238 5671
rect 13204 5637 13233 5641
rect 13233 5637 13238 5641
rect 13664 5657 13698 5671
rect 13664 5637 13669 5657
rect 13669 5637 13698 5657
rect 13852 5705 13886 5739
rect 14128 5711 14160 5739
rect 14160 5711 14162 5739
rect 14128 5705 14162 5711
rect 14036 5637 14070 5671
rect 13302 5570 13336 5604
rect 11117 5403 11151 5437
rect 11209 5403 11243 5437
rect 11301 5403 11335 5437
rect 11393 5403 11427 5437
rect 11485 5403 11519 5437
rect 11577 5403 11611 5437
rect 11669 5403 11703 5437
rect 11761 5403 11795 5437
rect 11853 5403 11887 5437
rect 11945 5403 11979 5437
rect 12037 5403 12071 5437
rect 12129 5403 12163 5437
rect 12221 5403 12255 5437
rect 12313 5403 12347 5437
rect 12405 5403 12439 5437
rect 12497 5403 12531 5437
rect 14312 5588 14341 5598
rect 14341 5588 14352 5598
rect 14312 5562 14352 5588
rect 15166 5769 15200 5803
rect 15906 5769 15940 5803
rect 14982 5715 14997 5735
rect 14997 5715 15016 5735
rect 15350 5731 15371 5735
rect 15371 5731 15384 5735
rect 14982 5701 15016 5715
rect 15350 5701 15384 5731
rect 15074 5637 15108 5667
rect 15074 5633 15103 5637
rect 15103 5633 15108 5637
rect 15534 5653 15568 5667
rect 15534 5633 15539 5653
rect 15539 5633 15568 5653
rect 15722 5701 15756 5735
rect 15998 5707 16030 5735
rect 16030 5707 16032 5735
rect 15998 5701 16032 5707
rect 15906 5633 15940 5667
rect 15172 5566 15206 5600
rect 12933 5399 12967 5433
rect 13025 5399 13059 5433
rect 13117 5399 13151 5433
rect 13209 5399 13243 5433
rect 13301 5399 13335 5433
rect 13393 5399 13427 5433
rect 13485 5399 13519 5433
rect 13577 5399 13611 5433
rect 13669 5399 13703 5433
rect 13761 5399 13795 5433
rect 13853 5399 13887 5433
rect 13945 5399 13979 5433
rect 14037 5399 14071 5433
rect 14129 5399 14163 5433
rect 14221 5399 14255 5433
rect 14313 5399 14347 5433
rect 16182 5584 16211 5600
rect 16211 5584 16216 5600
rect 16182 5564 16216 5584
rect 14803 5395 14837 5429
rect 14895 5395 14929 5429
rect 14987 5395 15021 5429
rect 15079 5395 15113 5429
rect 15171 5395 15205 5429
rect 15263 5395 15297 5429
rect 15355 5395 15389 5429
rect 15447 5395 15481 5429
rect 15539 5395 15573 5429
rect 15631 5395 15665 5429
rect 15723 5395 15757 5429
rect 15815 5395 15849 5429
rect 15907 5395 15941 5429
rect 15999 5395 16033 5429
rect 16091 5395 16125 5429
rect 16183 5395 16217 5429
rect 7692 5217 7726 5247
rect 7692 5213 7721 5217
rect 7721 5213 7726 5217
rect 8152 5233 8186 5247
rect 8152 5213 8157 5233
rect 8157 5213 8186 5233
rect 8340 5281 8374 5315
rect 8616 5287 8648 5315
rect 8648 5287 8650 5315
rect 8616 5281 8650 5287
rect 8524 5213 8558 5247
rect 7790 5146 7824 5180
rect 5551 4979 5585 5013
rect 5643 4979 5677 5013
rect 5735 4979 5769 5013
rect 5827 4979 5861 5013
rect 5919 4979 5953 5013
rect 6011 4979 6045 5013
rect 6103 4979 6137 5013
rect 6195 4979 6229 5013
rect 6287 4979 6321 5013
rect 6379 4979 6413 5013
rect 6471 4979 6505 5013
rect 6563 4979 6597 5013
rect 6655 4979 6689 5013
rect 6747 4979 6781 5013
rect 6839 4979 6873 5013
rect 6931 4979 6965 5013
rect 17108 5188 17142 5222
rect 8800 5164 8829 5180
rect 8829 5164 8834 5180
rect 8800 5144 8834 5164
rect 17190 5160 17224 5194
rect 9275 5077 9309 5111
rect 9367 5077 9401 5111
rect 9459 5077 9493 5111
rect 9551 5077 9585 5111
rect 9643 5077 9677 5111
rect 9735 5077 9769 5111
rect 9827 5077 9861 5111
rect 9919 5077 9953 5111
rect 10011 5077 10045 5111
rect 10103 5077 10137 5111
rect 10195 5077 10229 5111
rect 10287 5077 10321 5111
rect 10379 5077 10413 5111
rect 10471 5077 10505 5111
rect 10563 5077 10597 5111
rect 10655 5077 10689 5111
rect 7421 4975 7455 5009
rect 7513 4975 7547 5009
rect 7605 4975 7639 5009
rect 7697 4975 7731 5009
rect 7789 4975 7823 5009
rect 7881 4975 7915 5009
rect 7973 4975 8007 5009
rect 8065 4975 8099 5009
rect 8157 4975 8191 5009
rect 8249 4975 8283 5009
rect 8341 4975 8375 5009
rect 8433 4975 8467 5009
rect 8525 4975 8559 5009
rect 8617 4975 8651 5009
rect 8709 4975 8743 5009
rect 8801 4975 8835 5009
rect 9638 4907 9672 4941
rect 11145 5073 11179 5107
rect 11237 5073 11271 5107
rect 11329 5073 11363 5107
rect 11421 5073 11455 5107
rect 11513 5073 11547 5107
rect 11605 5073 11639 5107
rect 11697 5073 11731 5107
rect 11789 5073 11823 5107
rect 11881 5073 11915 5107
rect 11973 5073 12007 5107
rect 12065 5073 12099 5107
rect 12157 5073 12191 5107
rect 12249 5073 12283 5107
rect 12341 5073 12375 5107
rect 12433 5073 12467 5107
rect 12525 5073 12559 5107
rect 10378 4907 10412 4941
rect 9454 4853 9469 4873
rect 9469 4853 9488 4873
rect 9822 4869 9843 4873
rect 9843 4869 9856 4873
rect 9454 4839 9488 4853
rect 9822 4839 9856 4869
rect 9546 4775 9580 4805
rect 9546 4771 9575 4775
rect 9575 4771 9580 4775
rect 10006 4791 10040 4805
rect 10006 4771 10011 4791
rect 10011 4771 10040 4791
rect 10194 4839 10228 4873
rect 10470 4845 10502 4873
rect 10502 4845 10504 4873
rect 10470 4839 10504 4845
rect 10378 4771 10412 4805
rect 9646 4706 9680 4740
rect 10654 4722 10683 4732
rect 10683 4722 10694 4732
rect 10654 4696 10694 4722
rect 11508 4903 11542 4937
rect 12961 5069 12995 5103
rect 13053 5069 13087 5103
rect 13145 5069 13179 5103
rect 13237 5069 13271 5103
rect 13329 5069 13363 5103
rect 13421 5069 13455 5103
rect 13513 5069 13547 5103
rect 13605 5069 13639 5103
rect 13697 5069 13731 5103
rect 13789 5069 13823 5103
rect 13881 5069 13915 5103
rect 13973 5069 14007 5103
rect 14065 5069 14099 5103
rect 14157 5069 14191 5103
rect 14249 5069 14283 5103
rect 14341 5069 14375 5103
rect 12248 4903 12282 4937
rect 11324 4849 11339 4869
rect 11339 4849 11358 4869
rect 11692 4865 11713 4869
rect 11713 4865 11726 4869
rect 11324 4835 11358 4849
rect 11692 4835 11726 4865
rect 11416 4771 11450 4801
rect 11416 4767 11445 4771
rect 11445 4767 11450 4771
rect 11876 4787 11910 4801
rect 11876 4767 11881 4787
rect 11881 4767 11910 4787
rect 12064 4835 12098 4869
rect 12340 4841 12372 4869
rect 12372 4841 12374 4869
rect 12340 4835 12374 4841
rect 12248 4767 12282 4801
rect 11514 4700 11548 4734
rect 9275 4533 9309 4567
rect 9367 4533 9401 4567
rect 9459 4533 9493 4567
rect 9551 4533 9585 4567
rect 9643 4533 9677 4567
rect 9735 4533 9769 4567
rect 9827 4533 9861 4567
rect 9919 4533 9953 4567
rect 10011 4533 10045 4567
rect 10103 4533 10137 4567
rect 10195 4533 10229 4567
rect 10287 4533 10321 4567
rect 10379 4533 10413 4567
rect 10471 4533 10505 4567
rect 10563 4533 10597 4567
rect 10655 4533 10689 4567
rect 12530 4684 12564 4718
rect 13324 4899 13358 4933
rect 14831 5065 14865 5099
rect 14923 5065 14957 5099
rect 15015 5065 15049 5099
rect 15107 5065 15141 5099
rect 15199 5065 15233 5099
rect 15291 5065 15325 5099
rect 15383 5065 15417 5099
rect 15475 5065 15509 5099
rect 15567 5065 15601 5099
rect 15659 5065 15693 5099
rect 15751 5065 15785 5099
rect 15843 5065 15877 5099
rect 15935 5065 15969 5099
rect 16027 5065 16061 5099
rect 16119 5065 16153 5099
rect 16211 5065 16245 5099
rect 16932 5070 16970 5108
rect 14064 4899 14098 4933
rect 13140 4845 13155 4865
rect 13155 4845 13174 4865
rect 13508 4861 13529 4865
rect 13529 4861 13542 4865
rect 13140 4831 13174 4845
rect 13508 4831 13542 4861
rect 13232 4767 13266 4797
rect 13232 4763 13261 4767
rect 13261 4763 13266 4767
rect 13692 4783 13726 4797
rect 13692 4763 13697 4783
rect 13697 4763 13726 4783
rect 13880 4831 13914 4865
rect 14156 4837 14188 4865
rect 14188 4837 14190 4865
rect 14156 4831 14190 4837
rect 14064 4763 14098 4797
rect 13330 4696 13364 4730
rect 11145 4529 11179 4563
rect 11237 4529 11271 4563
rect 11329 4529 11363 4563
rect 11421 4529 11455 4563
rect 11513 4529 11547 4563
rect 11605 4529 11639 4563
rect 11697 4529 11731 4563
rect 11789 4529 11823 4563
rect 11881 4529 11915 4563
rect 11973 4529 12007 4563
rect 12065 4529 12099 4563
rect 12157 4529 12191 4563
rect 12249 4529 12283 4563
rect 12341 4529 12375 4563
rect 12433 4529 12467 4563
rect 12525 4529 12559 4563
rect 14340 4714 14369 4724
rect 14369 4714 14380 4724
rect 14340 4688 14380 4714
rect 15194 4895 15228 4929
rect 17564 5004 17602 5042
rect 15934 4895 15968 4929
rect 15010 4841 15025 4861
rect 15025 4841 15044 4861
rect 15378 4857 15399 4861
rect 15399 4857 15412 4861
rect 15010 4827 15044 4841
rect 15378 4827 15412 4857
rect 15102 4763 15136 4793
rect 15102 4759 15131 4763
rect 15131 4759 15136 4763
rect 15562 4779 15596 4793
rect 15562 4759 15567 4779
rect 15567 4759 15596 4779
rect 15750 4827 15784 4861
rect 16026 4833 16058 4861
rect 16058 4833 16060 4861
rect 16026 4827 16060 4833
rect 15934 4759 15968 4793
rect 15200 4692 15234 4726
rect 12961 4525 12995 4559
rect 13053 4525 13087 4559
rect 13145 4525 13179 4559
rect 13237 4525 13271 4559
rect 13329 4525 13363 4559
rect 13421 4525 13455 4559
rect 13513 4525 13547 4559
rect 13605 4525 13639 4559
rect 13697 4525 13731 4559
rect 13789 4525 13823 4559
rect 13881 4525 13915 4559
rect 13973 4525 14007 4559
rect 14065 4525 14099 4559
rect 14157 4525 14191 4559
rect 14249 4525 14283 4559
rect 14341 4525 14375 4559
rect 16210 4710 16239 4726
rect 16239 4710 16244 4726
rect 16210 4690 16244 4710
rect 14831 4521 14865 4555
rect 14923 4521 14957 4555
rect 15015 4521 15049 4555
rect 15107 4521 15141 4555
rect 15199 4521 15233 4555
rect 15291 4521 15325 4555
rect 15383 4521 15417 4555
rect 15475 4521 15509 4555
rect 15567 4521 15601 4555
rect 15659 4521 15693 4555
rect 15751 4521 15785 4555
rect 15843 4521 15877 4555
rect 15935 4521 15969 4555
rect 16027 4521 16061 4555
rect 16119 4521 16153 4555
rect 16211 4521 16245 4555
rect 6148 3088 6182 3122
rect 6244 3090 6278 3124
rect 1835 2271 1869 2305
rect 1927 2271 1961 2305
rect 2019 2271 2053 2305
rect 2111 2271 2145 2305
rect 2203 2271 2237 2305
rect 2295 2271 2329 2305
rect 2387 2271 2421 2305
rect 2479 2271 2513 2305
rect 2571 2271 2605 2305
rect 2663 2271 2697 2305
rect 2755 2271 2789 2305
rect 2847 2271 2881 2305
rect 2939 2271 2973 2305
rect 3031 2271 3065 2305
rect 3123 2271 3157 2305
rect 3215 2271 3249 2305
rect 2198 2101 2232 2135
rect 3705 2267 3739 2301
rect 3797 2267 3831 2301
rect 3889 2267 3923 2301
rect 3981 2267 4015 2301
rect 4073 2267 4107 2301
rect 4165 2267 4199 2301
rect 4257 2267 4291 2301
rect 4349 2267 4383 2301
rect 4441 2267 4475 2301
rect 4533 2267 4567 2301
rect 4625 2267 4659 2301
rect 4717 2267 4751 2301
rect 4809 2267 4843 2301
rect 4901 2267 4935 2301
rect 4993 2267 5027 2301
rect 5085 2267 5119 2301
rect 2938 2101 2972 2135
rect 2014 2047 2029 2067
rect 2029 2047 2048 2067
rect 2382 2063 2403 2067
rect 2403 2063 2416 2067
rect 2014 2033 2048 2047
rect 2382 2033 2416 2063
rect 2106 1969 2140 1999
rect 2106 1965 2135 1969
rect 2135 1965 2140 1969
rect 2566 1985 2600 1999
rect 2566 1965 2571 1985
rect 2571 1965 2600 1985
rect 2754 2033 2788 2067
rect 3030 2039 3062 2067
rect 3062 2039 3064 2067
rect 3030 2033 3064 2039
rect 2938 1965 2972 1999
rect 2206 1900 2240 1934
rect 3214 1916 3243 1926
rect 3243 1916 3254 1926
rect 3214 1890 3254 1916
rect 4068 2097 4102 2131
rect 5521 2263 5555 2297
rect 5613 2263 5647 2297
rect 5705 2263 5739 2297
rect 5797 2263 5831 2297
rect 5889 2263 5923 2297
rect 5981 2263 6015 2297
rect 6073 2263 6107 2297
rect 6165 2263 6199 2297
rect 6257 2263 6291 2297
rect 6349 2263 6383 2297
rect 6441 2263 6475 2297
rect 6533 2263 6567 2297
rect 6625 2263 6659 2297
rect 6717 2263 6751 2297
rect 6809 2263 6843 2297
rect 6901 2263 6935 2297
rect 4808 2097 4842 2131
rect 3884 2043 3899 2063
rect 3899 2043 3918 2063
rect 4252 2059 4273 2063
rect 4273 2059 4286 2063
rect 3884 2029 3918 2043
rect 4252 2029 4286 2059
rect 3976 1965 4010 1995
rect 3976 1961 4005 1965
rect 4005 1961 4010 1965
rect 4436 1981 4470 1995
rect 4436 1961 4441 1981
rect 4441 1961 4470 1981
rect 4624 2029 4658 2063
rect 4900 2035 4932 2063
rect 4932 2035 4934 2063
rect 4900 2029 4934 2035
rect 4808 1961 4842 1995
rect 4074 1894 4108 1928
rect 1835 1727 1869 1761
rect 1927 1727 1961 1761
rect 2019 1727 2053 1761
rect 2111 1727 2145 1761
rect 2203 1727 2237 1761
rect 2295 1727 2329 1761
rect 2387 1727 2421 1761
rect 2479 1727 2513 1761
rect 2571 1727 2605 1761
rect 2663 1727 2697 1761
rect 2755 1727 2789 1761
rect 2847 1727 2881 1761
rect 2939 1727 2973 1761
rect 3031 1727 3065 1761
rect 3123 1727 3157 1761
rect 3215 1727 3249 1761
rect 5090 1912 5113 1922
rect 5113 1912 5124 1922
rect 5090 1886 5124 1912
rect 5884 2093 5918 2127
rect 7391 2259 7425 2293
rect 7483 2259 7517 2293
rect 7575 2259 7609 2293
rect 7667 2259 7701 2293
rect 7759 2259 7793 2293
rect 7851 2259 7885 2293
rect 7943 2259 7977 2293
rect 8035 2259 8069 2293
rect 8127 2259 8161 2293
rect 8219 2259 8253 2293
rect 8311 2259 8345 2293
rect 8403 2259 8437 2293
rect 8495 2259 8529 2293
rect 8587 2259 8621 2293
rect 8679 2259 8713 2293
rect 8771 2259 8805 2293
rect 6624 2093 6658 2127
rect 5700 2039 5715 2059
rect 5715 2039 5734 2059
rect 6068 2055 6089 2059
rect 6089 2055 6102 2059
rect 5700 2025 5734 2039
rect 6068 2025 6102 2055
rect 5792 1961 5826 1991
rect 5792 1957 5821 1961
rect 5821 1957 5826 1961
rect 6252 1977 6286 1991
rect 6252 1957 6257 1977
rect 6257 1957 6286 1977
rect 6440 2025 6474 2059
rect 6716 2031 6748 2059
rect 6748 2031 6750 2059
rect 6716 2025 6750 2031
rect 6624 1957 6658 1991
rect 5890 1890 5924 1924
rect 3705 1723 3739 1757
rect 3797 1723 3831 1757
rect 3889 1723 3923 1757
rect 3981 1723 4015 1757
rect 4073 1723 4107 1757
rect 4165 1723 4199 1757
rect 4257 1723 4291 1757
rect 4349 1723 4383 1757
rect 4441 1723 4475 1757
rect 4533 1723 4567 1757
rect 4625 1723 4659 1757
rect 4717 1723 4751 1757
rect 4809 1723 4843 1757
rect 4901 1723 4935 1757
rect 4993 1723 5027 1757
rect 5085 1723 5119 1757
rect 6900 1908 6929 1918
rect 6929 1908 6940 1918
rect 6900 1882 6940 1908
rect 7754 2089 7788 2123
rect 9205 2257 9239 2291
rect 9297 2257 9331 2291
rect 9389 2257 9423 2291
rect 9481 2257 9515 2291
rect 9573 2257 9607 2291
rect 9665 2257 9699 2291
rect 9757 2257 9791 2291
rect 9849 2257 9883 2291
rect 9941 2257 9975 2291
rect 10033 2257 10067 2291
rect 10125 2257 10159 2291
rect 10217 2257 10251 2291
rect 10309 2257 10343 2291
rect 10401 2257 10435 2291
rect 10493 2257 10527 2291
rect 10585 2257 10619 2291
rect 8494 2089 8528 2123
rect 7570 2035 7585 2055
rect 7585 2035 7604 2055
rect 7938 2051 7959 2055
rect 7959 2051 7972 2055
rect 7570 2021 7604 2035
rect 7938 2021 7972 2051
rect 7662 1957 7696 1987
rect 7662 1953 7691 1957
rect 7691 1953 7696 1957
rect 8122 1973 8156 1987
rect 8122 1953 8127 1973
rect 8127 1953 8156 1973
rect 8310 2021 8344 2055
rect 8586 2027 8618 2055
rect 8618 2027 8620 2055
rect 8586 2021 8620 2027
rect 8494 1953 8528 1987
rect 7760 1886 7794 1920
rect 5521 1719 5555 1753
rect 5613 1719 5647 1753
rect 5705 1719 5739 1753
rect 5797 1719 5831 1753
rect 5889 1719 5923 1753
rect 5981 1719 6015 1753
rect 6073 1719 6107 1753
rect 6165 1719 6199 1753
rect 6257 1719 6291 1753
rect 6349 1719 6383 1753
rect 6441 1719 6475 1753
rect 6533 1719 6567 1753
rect 6625 1719 6659 1753
rect 6717 1719 6751 1753
rect 6809 1719 6843 1753
rect 6901 1719 6935 1753
rect 8770 1904 8799 1920
rect 8799 1904 8804 1920
rect 8770 1884 8804 1904
rect 9568 2087 9602 2121
rect 11075 2253 11109 2287
rect 11167 2253 11201 2287
rect 11259 2253 11293 2287
rect 11351 2253 11385 2287
rect 11443 2253 11477 2287
rect 11535 2253 11569 2287
rect 11627 2253 11661 2287
rect 11719 2253 11753 2287
rect 11811 2253 11845 2287
rect 11903 2253 11937 2287
rect 11995 2253 12029 2287
rect 12087 2253 12121 2287
rect 12179 2253 12213 2287
rect 12271 2253 12305 2287
rect 12363 2253 12397 2287
rect 12455 2253 12489 2287
rect 10308 2087 10342 2121
rect 9384 2033 9399 2053
rect 9399 2033 9418 2053
rect 9752 2049 9773 2053
rect 9773 2049 9786 2053
rect 9384 2019 9418 2033
rect 9752 2019 9786 2049
rect 9476 1955 9510 1985
rect 9476 1951 9505 1955
rect 9505 1951 9510 1955
rect 9936 1971 9970 1985
rect 9936 1951 9941 1971
rect 9941 1951 9970 1971
rect 10124 2019 10158 2053
rect 10400 2025 10432 2053
rect 10432 2025 10434 2053
rect 10400 2019 10434 2025
rect 10308 1951 10342 1985
rect 9574 1884 9610 1918
rect 7391 1715 7425 1749
rect 7483 1715 7517 1749
rect 7575 1715 7609 1749
rect 7667 1715 7701 1749
rect 7759 1715 7793 1749
rect 7851 1715 7885 1749
rect 7943 1715 7977 1749
rect 8035 1715 8069 1749
rect 8127 1715 8161 1749
rect 8219 1715 8253 1749
rect 8311 1715 8345 1749
rect 8403 1715 8437 1749
rect 8495 1715 8529 1749
rect 8587 1715 8621 1749
rect 8679 1715 8713 1749
rect 8771 1715 8805 1749
rect 10584 1902 10613 1912
rect 10613 1902 10624 1912
rect 10584 1876 10624 1902
rect 11438 2083 11472 2117
rect 12891 2249 12925 2283
rect 12983 2249 13017 2283
rect 13075 2249 13109 2283
rect 13167 2249 13201 2283
rect 13259 2249 13293 2283
rect 13351 2249 13385 2283
rect 13443 2249 13477 2283
rect 13535 2249 13569 2283
rect 13627 2249 13661 2283
rect 13719 2249 13753 2283
rect 13811 2249 13845 2283
rect 13903 2249 13937 2283
rect 13995 2249 14029 2283
rect 14087 2249 14121 2283
rect 14179 2249 14213 2283
rect 14271 2249 14305 2283
rect 12178 2083 12212 2117
rect 11254 2029 11269 2049
rect 11269 2029 11288 2049
rect 11622 2045 11643 2049
rect 11643 2045 11656 2049
rect 11254 2015 11288 2029
rect 11622 2015 11656 2045
rect 11346 1951 11380 1981
rect 11346 1947 11375 1951
rect 11375 1947 11380 1951
rect 11806 1967 11840 1981
rect 11806 1947 11811 1967
rect 11811 1947 11840 1967
rect 11994 2015 12028 2049
rect 12270 2021 12302 2049
rect 12302 2021 12304 2049
rect 12270 2015 12304 2021
rect 12178 1947 12212 1981
rect 11444 1880 11478 1914
rect 9205 1713 9239 1747
rect 9297 1713 9331 1747
rect 9389 1713 9423 1747
rect 9481 1713 9515 1747
rect 9573 1713 9607 1747
rect 9665 1713 9699 1747
rect 9757 1713 9791 1747
rect 9849 1713 9883 1747
rect 9941 1713 9975 1747
rect 10033 1713 10067 1747
rect 10125 1713 10159 1747
rect 10217 1713 10251 1747
rect 10309 1713 10343 1747
rect 10401 1713 10435 1747
rect 10493 1713 10527 1747
rect 10585 1713 10619 1747
rect 12454 1898 12483 1912
rect 12483 1898 12488 1912
rect 12454 1878 12488 1898
rect 13254 2079 13288 2113
rect 14761 2245 14795 2279
rect 14853 2245 14887 2279
rect 14945 2245 14979 2279
rect 15037 2245 15071 2279
rect 15129 2245 15163 2279
rect 15221 2245 15255 2279
rect 15313 2245 15347 2279
rect 15405 2245 15439 2279
rect 15497 2245 15531 2279
rect 15589 2245 15623 2279
rect 15681 2245 15715 2279
rect 15773 2245 15807 2279
rect 15865 2245 15899 2279
rect 15957 2245 15991 2279
rect 16049 2245 16083 2279
rect 16141 2245 16175 2279
rect 13994 2079 14028 2113
rect 13070 2025 13085 2045
rect 13085 2025 13104 2045
rect 13438 2041 13459 2045
rect 13459 2041 13472 2045
rect 13070 2011 13104 2025
rect 13438 2011 13472 2041
rect 13162 1947 13196 1977
rect 13162 1943 13191 1947
rect 13191 1943 13196 1947
rect 13622 1963 13656 1977
rect 13622 1943 13627 1963
rect 13627 1943 13656 1963
rect 13810 2011 13844 2045
rect 14086 2017 14118 2045
rect 14118 2017 14120 2045
rect 14086 2011 14120 2017
rect 13994 1943 14028 1977
rect 13260 1876 13294 1910
rect 11075 1709 11109 1743
rect 11167 1709 11201 1743
rect 11259 1709 11293 1743
rect 11351 1709 11385 1743
rect 11443 1709 11477 1743
rect 11535 1709 11569 1743
rect 11627 1709 11661 1743
rect 11719 1709 11753 1743
rect 11811 1709 11845 1743
rect 11903 1709 11937 1743
rect 11995 1709 12029 1743
rect 12087 1709 12121 1743
rect 12179 1709 12213 1743
rect 12271 1709 12305 1743
rect 12363 1709 12397 1743
rect 12455 1709 12489 1743
rect 14270 1894 14299 1904
rect 14299 1894 14310 1904
rect 14270 1868 14310 1894
rect 15124 2075 15158 2109
rect 15864 2075 15898 2109
rect 14940 2021 14955 2041
rect 14955 2021 14974 2041
rect 15308 2037 15329 2041
rect 15329 2037 15342 2041
rect 14940 2007 14974 2021
rect 15308 2007 15342 2037
rect 15032 1943 15066 1973
rect 15032 1939 15061 1943
rect 15061 1939 15066 1943
rect 15492 1959 15526 1973
rect 15492 1939 15497 1959
rect 15497 1939 15526 1959
rect 15680 2007 15714 2041
rect 15956 2013 15988 2041
rect 15988 2013 15990 2041
rect 15956 2007 15990 2013
rect 15864 1939 15898 1973
rect 15130 1872 15164 1906
rect 12891 1705 12925 1739
rect 12983 1705 13017 1739
rect 13075 1705 13109 1739
rect 13167 1705 13201 1739
rect 13259 1705 13293 1739
rect 13351 1705 13385 1739
rect 13443 1705 13477 1739
rect 13535 1705 13569 1739
rect 13627 1705 13661 1739
rect 13719 1705 13753 1739
rect 13811 1705 13845 1739
rect 13903 1705 13937 1739
rect 13995 1705 14029 1739
rect 14087 1705 14121 1739
rect 14179 1705 14213 1739
rect 14271 1705 14305 1739
rect 16150 1890 16169 1918
rect 16169 1890 16186 1918
rect 16150 1884 16186 1890
rect 14761 1701 14795 1735
rect 14853 1701 14887 1735
rect 14945 1701 14979 1735
rect 15037 1701 15071 1735
rect 15129 1701 15163 1735
rect 15221 1701 15255 1735
rect 15313 1701 15347 1735
rect 15405 1701 15439 1735
rect 15497 1701 15531 1735
rect 15589 1701 15623 1735
rect 15681 1701 15715 1735
rect 15773 1701 15807 1735
rect 15865 1701 15899 1735
rect 15957 1701 15991 1735
rect 16049 1701 16083 1735
rect 16141 1701 16175 1735
<< metal1 >>
rect 6603 17576 9539 17587
rect 6603 17504 6646 17576
rect 6722 17568 9539 17576
rect 6722 17532 9496 17568
rect 9532 17532 9539 17568
rect 6722 17504 9539 17532
rect 6603 17497 9539 17504
rect 9573 17572 13733 17587
rect 9573 17536 9596 17572
rect 9632 17536 13733 17572
rect 9573 17497 13733 17536
rect 9045 17054 11482 17055
rect 9036 17042 11482 17054
rect 9036 16986 11414 17042
rect 11474 16986 11482 17042
rect 9036 16977 11482 16986
rect 9036 16700 9124 16977
rect 6578 15408 6682 15424
rect 6578 15356 6608 15408
rect 6660 15356 6682 15408
rect 6578 15342 6682 15356
rect 9036 14096 9126 16700
rect 9430 16608 10074 16618
rect 9430 16587 9552 16608
rect 9604 16587 10074 16608
rect 9430 16553 9459 16587
rect 9493 16553 9551 16587
rect 9604 16554 9643 16587
rect 9585 16553 9643 16554
rect 9677 16553 9735 16587
rect 9769 16553 9827 16587
rect 9861 16553 9919 16587
rect 9953 16553 10011 16587
rect 10045 16553 10074 16587
rect 9430 16522 10074 16553
rect 9508 16276 9568 16522
rect 10908 16390 11110 16422
rect 10908 16388 10968 16390
rect 9994 16374 10968 16388
rect 9994 16336 10006 16374
rect 10040 16336 10968 16374
rect 9994 16324 10968 16336
rect 11038 16388 11110 16390
rect 11038 16324 11221 16388
rect 9994 16322 11221 16324
rect 10908 16296 11110 16322
rect 9508 16242 9516 16276
rect 9550 16242 9568 16276
rect 9508 16222 9568 16242
rect 9598 16278 9708 16292
rect 9598 16244 9636 16278
rect 9670 16244 9708 16278
rect 9598 16236 9708 16244
rect 9632 16074 9663 16236
rect 9430 16058 10074 16074
rect 9430 16043 9938 16058
rect 9996 16043 10074 16058
rect 9430 16009 9459 16043
rect 9493 16009 9551 16043
rect 9585 16009 9643 16043
rect 9677 16009 9735 16043
rect 9769 16009 9827 16043
rect 9861 16009 9919 16043
rect 9996 16009 10011 16043
rect 10045 16009 10074 16043
rect 9430 16004 9938 16009
rect 9996 16004 10074 16009
rect 9430 15978 10074 16004
rect 9528 15858 9988 15874
rect 9528 15843 9708 15858
rect 9770 15843 9988 15858
rect 9528 15809 9557 15843
rect 9591 15809 9649 15843
rect 9683 15809 9708 15843
rect 9775 15809 9833 15843
rect 9867 15809 9925 15843
rect 9959 15809 9988 15843
rect 9528 15798 9708 15809
rect 9770 15798 9988 15809
rect 9528 15778 9988 15798
rect 9536 15554 9612 15570
rect 9738 15554 9792 15778
rect 11155 15617 11221 16322
rect 11570 15752 12214 15764
rect 11570 15733 11674 15752
rect 11742 15733 12214 15752
rect 11570 15699 11599 15733
rect 11633 15699 11674 15733
rect 11742 15699 11783 15733
rect 11817 15699 11875 15733
rect 11909 15699 11967 15733
rect 12001 15699 12059 15733
rect 12093 15699 12151 15733
rect 12185 15699 12214 15733
rect 11570 15690 11674 15699
rect 11742 15690 12214 15699
rect 11570 15668 12214 15690
rect 9536 15514 9550 15554
rect 9592 15514 9612 15554
rect 9536 15498 9612 15514
rect 9728 15544 9796 15554
rect 11155 15551 12009 15617
rect 11753 15548 11819 15551
rect 9728 15504 9740 15544
rect 9782 15504 9796 15544
rect 9546 15330 9600 15498
rect 9728 15492 9796 15504
rect 9920 15486 10006 15494
rect 9920 15474 9938 15486
rect 9920 15440 9932 15474
rect 9920 15432 9938 15440
rect 9992 15432 10006 15486
rect 9920 15420 10006 15432
rect 10156 15442 11818 15500
rect 10156 15436 11819 15442
rect 9728 15330 9796 15332
rect 9528 15316 9988 15330
rect 9528 15299 9860 15316
rect 9928 15299 9988 15316
rect 9528 15265 9557 15299
rect 9591 15265 9649 15299
rect 9683 15265 9741 15299
rect 9775 15265 9833 15299
rect 9959 15265 9988 15299
rect 9528 15254 9860 15265
rect 9928 15254 9988 15265
rect 9528 15234 9988 15254
rect 9440 15036 10084 15054
rect 9440 15023 9544 15036
rect 9610 15023 10084 15036
rect 9440 14989 9469 15023
rect 9503 14989 9544 15023
rect 9610 14989 9653 15023
rect 9687 14989 9745 15023
rect 9779 14989 9837 15023
rect 9871 14989 9929 15023
rect 9963 14989 10021 15023
rect 10055 14989 10084 15023
rect 9440 14970 9544 14989
rect 9610 14970 10084 14989
rect 9440 14958 10084 14970
rect 9518 14712 9578 14958
rect 10156 14926 10220 15436
rect 11753 15418 11819 15436
rect 11540 15392 11644 15408
rect 11540 15340 11570 15392
rect 11622 15384 11644 15392
rect 11630 15348 11644 15384
rect 11753 15382 11766 15418
rect 11800 15382 11819 15418
rect 11753 15374 11819 15382
rect 11622 15340 11644 15348
rect 11540 15326 11644 15340
rect 11943 15364 12009 15551
rect 12140 15424 12196 15428
rect 12140 15416 12362 15424
rect 12140 15382 12152 15416
rect 12186 15382 12362 15416
rect 12140 15374 12362 15382
rect 12140 15370 12196 15374
rect 11943 15328 11960 15364
rect 11994 15328 12009 15364
rect 11852 15298 11910 15314
rect 11310 15294 11910 15298
rect 10712 15248 11172 15264
rect 11310 15260 11864 15294
rect 11898 15260 11910 15294
rect 11310 15254 11910 15260
rect 10712 15233 11092 15248
rect 10712 15199 10741 15233
rect 10775 15199 10833 15233
rect 10867 15199 10925 15233
rect 10959 15199 11017 15233
rect 11051 15199 11092 15233
rect 10712 15186 11092 15199
rect 11160 15186 11172 15248
rect 10712 15168 11172 15186
rect 11312 15140 11392 15254
rect 11852 15248 11910 15254
rect 11943 15250 12009 15328
rect 11066 15132 11392 15140
rect 10002 14914 10220 14926
rect 10002 14880 10018 14914
rect 10052 14880 10220 14914
rect 10002 14862 10220 14880
rect 10252 15064 10982 15116
rect 11066 15096 11106 15132
rect 11146 15096 11392 15132
rect 11570 15202 12214 15220
rect 11570 15189 12076 15202
rect 12144 15189 12214 15202
rect 11570 15155 11599 15189
rect 11633 15155 11691 15189
rect 11725 15155 11783 15189
rect 11817 15155 11875 15189
rect 11909 15155 11967 15189
rect 12001 15155 12059 15189
rect 12144 15155 12151 15189
rect 12185 15155 12214 15189
rect 11570 15140 12076 15155
rect 12144 15140 12214 15155
rect 11570 15124 12214 15140
rect 11066 15082 11392 15096
rect 9518 14678 9526 14712
rect 9560 14678 9578 14712
rect 9518 14658 9578 14678
rect 9608 14714 9718 14728
rect 9608 14680 9646 14714
rect 9680 14680 9718 14714
rect 9608 14672 9718 14680
rect 9642 14510 9673 14672
rect 9440 14492 10084 14510
rect 9440 14479 9974 14492
rect 10040 14479 10084 14492
rect 9440 14445 9469 14479
rect 9503 14445 9561 14479
rect 9595 14445 9653 14479
rect 9687 14445 9745 14479
rect 9779 14445 9837 14479
rect 9871 14445 9929 14479
rect 9963 14445 9974 14479
rect 10055 14445 10084 14479
rect 9440 14426 9974 14445
rect 10040 14426 10084 14445
rect 9440 14414 10084 14426
rect 9538 14298 9998 14310
rect 9538 14279 9644 14298
rect 9716 14279 9998 14298
rect 9538 14245 9567 14279
rect 9601 14245 9644 14279
rect 9716 14245 9751 14279
rect 9785 14245 9843 14279
rect 9877 14245 9935 14279
rect 9969 14245 9998 14279
rect 9538 14228 9644 14245
rect 9716 14228 9998 14245
rect 9538 14214 9998 14228
rect 8118 14072 9126 14096
rect 8118 14032 8130 14072
rect 8172 14032 9126 14072
rect 8118 14018 9126 14032
rect 9546 13990 9622 14008
rect 9750 13990 9796 14214
rect 7636 13948 7724 13974
rect 7636 13936 7674 13948
rect 7636 13882 7652 13936
rect 7714 13914 7724 13948
rect 9546 13950 9560 13990
rect 9602 13950 9622 13990
rect 9546 13934 9622 13950
rect 9738 13980 9806 13990
rect 9738 13940 9750 13980
rect 9792 13940 9806 13980
rect 7704 13882 7724 13914
rect 7636 13856 7724 13882
rect 9554 13766 9608 13934
rect 9738 13928 9806 13940
rect 9928 13884 10100 13898
rect 9928 13868 9992 13884
rect 9928 13834 9940 13868
rect 9976 13834 9992 13868
rect 9928 13822 9992 13834
rect 10052 13822 10100 13884
rect 9928 13804 10100 13822
rect 9538 13754 9998 13766
rect 9538 13735 9846 13754
rect 9918 13735 9998 13754
rect 9538 13701 9567 13735
rect 9601 13701 9659 13735
rect 9693 13701 9751 13735
rect 9785 13701 9843 13735
rect 9918 13701 9935 13735
rect 9969 13701 9998 13735
rect 9538 13684 9846 13701
rect 9918 13684 9998 13701
rect 9538 13670 9998 13684
rect 9432 13368 10076 13386
rect 9432 13355 9538 13368
rect 9610 13355 10076 13368
rect 9432 13321 9461 13355
rect 9495 13321 9538 13355
rect 9610 13321 9645 13355
rect 9679 13321 9737 13355
rect 9771 13321 9829 13355
rect 9863 13321 9921 13355
rect 9955 13321 10013 13355
rect 10047 13321 10076 13355
rect 9432 13302 9538 13321
rect 9610 13302 10076 13321
rect 9432 13290 10076 13302
rect 10252 13350 10304 15064
rect 10930 14940 10982 15064
rect 10732 14935 10868 14936
rect 10524 14922 10868 14935
rect 10524 14888 10786 14922
rect 10820 14888 10868 14922
rect 10524 14862 10868 14888
rect 10902 14922 10982 14940
rect 10902 14888 10926 14922
rect 10962 14888 10982 14922
rect 10902 14874 10982 14888
rect 10524 14857 10807 14862
rect 10524 13955 10602 14857
rect 10712 14700 11172 14720
rect 10712 14689 10756 14700
rect 10824 14689 11172 14700
rect 10712 14655 10741 14689
rect 10824 14655 10833 14689
rect 10867 14655 10925 14689
rect 10959 14655 11017 14689
rect 11051 14655 11109 14689
rect 11143 14655 11172 14689
rect 10712 14638 10756 14655
rect 10824 14638 11172 14655
rect 10712 14624 11172 14638
rect 10786 14278 11430 14298
rect 10786 14267 11312 14278
rect 11380 14267 11430 14278
rect 10786 14233 10815 14267
rect 10849 14233 10907 14267
rect 10941 14233 10999 14267
rect 11033 14233 11091 14267
rect 11125 14233 11183 14267
rect 11217 14233 11275 14267
rect 11309 14233 11312 14267
rect 11401 14233 11430 14267
rect 10786 14216 11312 14233
rect 11380 14216 11430 14233
rect 10786 14202 11430 14216
rect 12309 14161 12359 15374
rect 13643 14697 13733 17497
rect 16187 16853 18657 16863
rect 16187 16847 20570 16853
rect 16187 16833 23479 16847
rect 16187 16367 16217 16833
rect 18512 16823 23479 16833
rect 19995 16817 23479 16823
rect 21207 16806 21237 16817
rect 16400 16400 16466 16420
rect 16400 16367 16416 16400
rect 16187 16366 16416 16367
rect 16452 16366 16466 16400
rect 16187 16337 16466 16366
rect 16496 16392 17234 16412
rect 16496 16388 17184 16392
rect 16496 16354 16502 16388
rect 16540 16358 17184 16388
rect 17222 16358 17234 16392
rect 16540 16354 17234 16358
rect 16496 16338 17234 16354
rect 17264 16396 18106 16418
rect 17264 16384 18048 16396
rect 17264 16350 17278 16384
rect 17312 16362 18048 16384
rect 18082 16362 18106 16396
rect 17312 16350 18106 16362
rect 16400 16336 16466 16337
rect 17264 16328 18106 16350
rect 18138 16392 18200 16416
rect 18138 16358 18150 16392
rect 18186 16390 18200 16392
rect 18656 16390 18722 16410
rect 18186 16388 18314 16390
rect 18656 16388 18672 16390
rect 18186 16358 18672 16388
rect 18138 16356 18672 16358
rect 18708 16356 18722 16390
rect 18138 16348 18722 16356
rect 18194 16342 18722 16348
rect 18512 16327 18722 16342
rect 18752 16382 19490 16402
rect 18752 16378 19440 16382
rect 18752 16344 18758 16378
rect 18796 16348 19440 16378
rect 19478 16348 19490 16382
rect 18796 16344 19490 16348
rect 18752 16328 19490 16344
rect 19520 16386 20362 16408
rect 19520 16374 20304 16386
rect 19520 16340 19534 16374
rect 19568 16352 20304 16374
rect 20338 16352 20362 16386
rect 19568 16340 20362 16352
rect 18656 16326 18722 16327
rect 19520 16318 20362 16340
rect 20394 16392 20456 16406
rect 21418 16392 21486 16404
rect 20394 16384 21486 16392
rect 20394 16382 21436 16384
rect 20394 16348 20406 16382
rect 20442 16350 21436 16382
rect 21472 16350 21486 16384
rect 20442 16348 21486 16350
rect 20394 16338 21486 16348
rect 20440 16336 21486 16338
rect 21418 16320 21486 16336
rect 21516 16376 22254 16396
rect 21516 16372 22204 16376
rect 21516 16338 21522 16372
rect 21560 16342 22204 16372
rect 22242 16342 22254 16376
rect 21560 16338 22254 16342
rect 21516 16322 22254 16338
rect 22284 16380 23126 16402
rect 22284 16368 23068 16380
rect 22284 16334 22298 16368
rect 22332 16346 23068 16368
rect 23102 16346 23126 16380
rect 22332 16334 23126 16346
rect 22284 16312 23126 16334
rect 23158 16376 23220 16400
rect 23158 16342 23170 16376
rect 23206 16374 23220 16376
rect 23449 16374 23479 16817
rect 23206 16344 23479 16374
rect 23206 16342 23220 16344
rect 23158 16332 23220 16342
rect 21575 16086 21605 16182
rect 23373 15607 23403 16344
rect 23372 15606 23403 15607
rect 22975 15577 23403 15606
rect 22975 14749 23005 15577
rect 22975 14719 23731 14749
rect 13643 14607 22797 14697
rect 23701 14614 23731 14719
rect 24138 14714 24198 14726
rect 24138 14662 24144 14714
rect 24196 14662 24198 14714
rect 24138 14650 24198 14662
rect 24138 14616 24150 14650
rect 24186 14616 24198 14650
rect 12604 14268 13156 14282
rect 12604 14251 12878 14268
rect 12946 14251 13156 14268
rect 12604 14217 12633 14251
rect 12667 14217 12725 14251
rect 12759 14217 12817 14251
rect 12851 14217 12878 14251
rect 12946 14217 13001 14251
rect 13035 14217 13093 14251
rect 13127 14217 13156 14251
rect 12604 14206 12878 14217
rect 12946 14206 13156 14217
rect 12604 14186 13156 14206
rect 12309 14156 12360 14161
rect 12309 14150 12956 14156
rect 12309 14116 12778 14150
rect 12814 14116 12956 14150
rect 12309 14109 12956 14116
rect 12352 14108 12956 14109
rect 13643 14098 13733 14607
rect 22618 14599 22797 14607
rect 22618 14580 23581 14599
rect 22618 14546 23530 14580
rect 23568 14546 23581 14580
rect 22618 14509 23581 14546
rect 23644 14562 23732 14614
rect 24138 14578 24198 14616
rect 23644 14528 23672 14562
rect 23708 14528 23732 14562
rect 22618 14508 22736 14509
rect 23644 14490 23732 14528
rect 24444 14564 24510 14620
rect 24444 14512 24452 14564
rect 24504 14512 24510 14564
rect 24444 14502 24510 14512
rect 24550 14588 24604 14620
rect 24550 14578 24556 14588
rect 24592 14578 24604 14588
rect 24550 14526 24552 14578
rect 24550 14502 24604 14526
rect 24684 14562 24770 14618
rect 24684 14536 24712 14562
rect 24746 14536 24770 14562
rect 25348 14598 28230 14610
rect 25348 14562 25364 14598
rect 25400 14562 28230 14598
rect 25348 14546 28230 14562
rect 24684 14484 24698 14536
rect 24750 14484 24770 14536
rect 24684 14434 24770 14484
rect 23850 14318 24212 14334
rect 23850 14258 23992 14318
rect 24054 14258 24212 14318
rect 23850 14240 24212 14258
rect 13142 14080 13733 14098
rect 12408 14014 12996 14074
rect 10785 13960 10863 14013
rect 12408 14002 12482 14014
rect 10785 13955 10812 13960
rect 10524 13926 10812 13955
rect 10846 13926 10863 13960
rect 10524 13877 10863 13926
rect 10252 13340 10338 13350
rect 9510 13044 9570 13290
rect 10252 13288 10260 13340
rect 10322 13288 10338 13340
rect 10252 13280 10338 13288
rect 10252 13212 10304 13280
rect 9998 13204 10304 13212
rect 9998 13170 10010 13204
rect 10044 13170 10304 13204
rect 9998 13160 10304 13170
rect 10524 13069 10602 13877
rect 10964 13874 11034 13920
rect 10964 13822 10974 13874
rect 11026 13822 11034 13874
rect 10964 13782 11034 13822
rect 11062 13914 11130 13970
rect 11062 13862 11072 13914
rect 11124 13862 11130 13914
rect 11062 13784 11130 13862
rect 11164 13954 11236 13972
rect 11164 13916 11174 13954
rect 11210 13916 11236 13954
rect 11164 13870 11236 13916
rect 11164 13814 11170 13870
rect 11222 13814 11236 13870
rect 11756 13902 12216 13924
rect 11756 13893 11790 13902
rect 11858 13893 12216 13902
rect 11756 13859 11785 13893
rect 11858 13859 11877 13893
rect 11911 13859 11969 13893
rect 12003 13859 12061 13893
rect 12095 13859 12153 13893
rect 12187 13859 12216 13893
rect 11164 13788 11236 13814
rect 11342 13836 11628 13856
rect 11342 13798 11356 13836
rect 11394 13798 11628 13836
rect 11756 13840 11790 13859
rect 11858 13840 12216 13859
rect 11756 13828 12216 13840
rect 12408 13914 12480 14002
rect 12718 13964 12858 13976
rect 12598 13932 12686 13958
rect 12598 13920 12636 13932
rect 11342 13782 11628 13798
rect 11547 13769 11628 13782
rect 12408 13770 12478 13914
rect 12598 13866 12614 13920
rect 12676 13898 12686 13932
rect 12666 13866 12686 13898
rect 12718 13888 12748 13964
rect 12828 13942 12858 13964
rect 12924 13956 12996 14014
rect 13080 14056 13733 14080
rect 13080 14016 13092 14056
rect 13134 14016 13733 14056
rect 13080 14008 13733 14016
rect 13080 14002 13726 14008
rect 12828 13888 12856 13942
rect 12902 13940 12996 13956
rect 12902 13904 12934 13940
rect 12972 13904 12996 13940
rect 12902 13888 12996 13904
rect 12718 13874 12856 13888
rect 12598 13840 12686 13866
rect 10786 13738 11430 13754
rect 10786 13723 10824 13738
rect 10892 13723 11430 13738
rect 10786 13689 10815 13723
rect 10892 13689 10907 13723
rect 10941 13689 10999 13723
rect 11033 13689 11091 13723
rect 11125 13689 11183 13723
rect 11217 13689 11275 13723
rect 11309 13689 11367 13723
rect 11401 13689 11430 13723
rect 11547 13695 12025 13769
rect 12082 13748 12478 13770
rect 12082 13714 12124 13748
rect 12158 13714 12478 13748
rect 12082 13698 12478 13714
rect 12604 13722 13156 13738
rect 10786 13676 10824 13689
rect 10892 13676 11430 13689
rect 10786 13658 11430 13676
rect 11951 13588 12025 13695
rect 12604 13660 12618 13722
rect 12686 13707 13156 13722
rect 12686 13673 12725 13707
rect 12759 13673 12817 13707
rect 12851 13673 12909 13707
rect 12943 13673 13001 13707
rect 13035 13673 13093 13707
rect 13127 13673 13156 13707
rect 12686 13660 13156 13673
rect 12604 13642 13156 13660
rect 11506 13538 11855 13561
rect 11506 13504 11796 13538
rect 11830 13504 11855 13538
rect 11506 13487 11855 13504
rect 11951 13554 11974 13588
rect 12008 13554 12025 13588
rect 10910 13434 11370 13456
rect 10910 13425 10946 13434
rect 11014 13425 11370 13434
rect 10910 13391 10939 13425
rect 11014 13391 11031 13425
rect 11065 13391 11123 13425
rect 11157 13391 11215 13425
rect 11249 13391 11307 13425
rect 11341 13391 11370 13425
rect 10910 13374 10946 13391
rect 11014 13374 11370 13391
rect 10910 13360 11370 13374
rect 11082 13322 11180 13328
rect 11082 13270 11102 13322
rect 11156 13270 11180 13322
rect 11506 13282 11580 13487
rect 11951 13473 12025 13554
rect 11756 13362 12216 13380
rect 11756 13349 12098 13362
rect 12166 13349 12216 13362
rect 11756 13315 11785 13349
rect 11819 13315 11877 13349
rect 11911 13315 11969 13349
rect 12003 13315 12061 13349
rect 12095 13315 12098 13349
rect 12187 13315 12216 13349
rect 11756 13300 12098 13315
rect 12166 13300 12216 13315
rect 11756 13284 12216 13300
rect 11082 13252 11180 13270
rect 11294 13262 11580 13282
rect 11294 13224 11304 13262
rect 11342 13224 11580 13262
rect 11294 13208 11580 13224
rect 9510 13010 9518 13044
rect 9552 13010 9570 13044
rect 9510 12990 9570 13010
rect 9600 13046 9710 13060
rect 9600 13012 9638 13046
rect 9672 13012 9710 13046
rect 9600 13004 9710 13012
rect 10524 13044 11043 13069
rect 10524 13010 10956 13044
rect 10990 13010 11043 13044
rect 9634 12842 9665 13004
rect 10524 12991 11043 13010
rect 11138 13066 11220 13138
rect 11138 13012 11158 13066
rect 11210 13012 11220 13066
rect 9432 12828 10076 12842
rect 9432 12811 9952 12828
rect 10024 12811 10076 12828
rect 9432 12777 9461 12811
rect 9495 12777 9553 12811
rect 9587 12777 9645 12811
rect 9679 12777 9737 12811
rect 9771 12777 9829 12811
rect 9863 12777 9921 12811
rect 10047 12777 10076 12811
rect 9432 12762 9952 12777
rect 10024 12762 10076 12777
rect 9432 12746 10076 12762
rect 9530 12626 9990 12642
rect 9530 12611 9596 12626
rect 9670 12611 9990 12626
rect 9530 12577 9559 12611
rect 9593 12577 9596 12611
rect 9685 12577 9743 12611
rect 9777 12577 9835 12611
rect 9869 12577 9927 12611
rect 9961 12577 9990 12611
rect 9530 12560 9596 12577
rect 9670 12560 9990 12577
rect 9530 12546 9990 12560
rect 9538 12322 9614 12348
rect 9738 12322 9788 12546
rect 9922 12374 10072 12388
rect 9922 12354 9968 12374
rect 9538 12282 9552 12322
rect 9594 12282 9614 12322
rect 9538 12266 9614 12282
rect 9730 12312 9798 12322
rect 9730 12272 9742 12312
rect 9784 12272 9798 12312
rect 9922 12320 9932 12354
rect 9922 12306 9968 12320
rect 10030 12306 10072 12374
rect 9922 12290 10072 12306
rect 9552 12098 9604 12266
rect 9730 12260 9798 12272
rect 10524 12105 10602 12991
rect 11138 12954 11220 13012
rect 10910 12900 11370 12912
rect 10910 12881 10958 12900
rect 11026 12881 11370 12900
rect 10910 12847 10939 12881
rect 11026 12847 11031 12881
rect 11065 12847 11123 12881
rect 11157 12847 11215 12881
rect 11249 12847 11307 12881
rect 11341 12847 11370 12881
rect 10910 12840 10958 12847
rect 11026 12840 11370 12847
rect 10910 12816 11370 12840
rect 10906 12416 11366 12436
rect 10906 12405 11242 12416
rect 11310 12405 11366 12416
rect 10906 12371 10935 12405
rect 10969 12371 11027 12405
rect 11061 12371 11119 12405
rect 11153 12371 11211 12405
rect 11337 12371 11366 12405
rect 10906 12354 11242 12371
rect 11310 12354 11366 12371
rect 10906 12340 11366 12354
rect 11296 12192 11364 12202
rect 11296 12140 11302 12192
rect 11354 12140 11364 12192
rect 11296 12134 11364 12140
rect 9530 12084 9990 12098
rect 9530 12067 9868 12084
rect 9942 12067 9990 12084
rect 9530 12033 9559 12067
rect 9593 12033 9651 12067
rect 9685 12033 9743 12067
rect 9777 12033 9835 12067
rect 9961 12033 9990 12067
rect 9530 12018 9868 12033
rect 9942 12018 9990 12033
rect 9530 12002 9990 12018
rect 10524 12096 11057 12105
rect 10524 12062 10980 12096
rect 11016 12062 11057 12096
rect 10524 12027 11057 12062
rect 11104 12102 11174 12110
rect 11104 12050 11112 12102
rect 11164 12050 11174 12102
rect 11104 12044 11174 12050
rect 9442 11804 10086 11822
rect 9442 11791 9522 11804
rect 9602 11791 10086 11804
rect 9442 11757 9471 11791
rect 9505 11757 9522 11791
rect 9602 11757 9655 11791
rect 9689 11757 9747 11791
rect 9781 11757 9839 11791
rect 9873 11757 9931 11791
rect 9965 11757 10023 11791
rect 10057 11757 10086 11791
rect 9442 11740 9522 11757
rect 9602 11740 10086 11757
rect 9442 11726 10086 11740
rect 9520 11480 9580 11726
rect 10524 11654 10602 12027
rect 10906 11876 11366 11892
rect 10906 11861 10964 11876
rect 11032 11861 11366 11876
rect 10906 11827 10935 11861
rect 11061 11827 11119 11861
rect 11153 11827 11211 11861
rect 11245 11827 11303 11861
rect 11337 11827 11366 11861
rect 10906 11814 10964 11827
rect 11032 11814 11366 11827
rect 10906 11796 11366 11814
rect 10004 11640 10602 11654
rect 10004 11606 10010 11640
rect 10046 11606 10602 11640
rect 10004 11576 10602 11606
rect 9520 11446 9528 11480
rect 9562 11446 9580 11480
rect 9520 11426 9580 11446
rect 9610 11482 9720 11496
rect 9610 11448 9648 11482
rect 9682 11448 9720 11482
rect 9610 11440 9720 11448
rect 9644 11278 9675 11440
rect 9442 11262 10086 11278
rect 9442 11247 9956 11262
rect 10036 11247 10086 11262
rect 9442 11213 9471 11247
rect 9505 11213 9563 11247
rect 9597 11213 9655 11247
rect 9689 11213 9747 11247
rect 9781 11213 9839 11247
rect 9873 11213 9931 11247
rect 10057 11213 10086 11247
rect 9442 11198 9956 11213
rect 10036 11198 10086 11213
rect 9442 11182 10086 11198
rect 9540 11058 10000 11078
rect 9540 11047 9588 11058
rect 9668 11047 10000 11058
rect 9540 11013 9569 11047
rect 9695 11013 9753 11047
rect 9787 11013 9845 11047
rect 9879 11013 9937 11047
rect 9971 11013 10000 11047
rect 9540 10994 9588 11013
rect 9668 10994 10000 11013
rect 9540 10982 10000 10994
rect 4970 10732 5202 10762
rect 4970 10730 5054 10732
rect 4970 10694 4982 10730
rect 5016 10694 5054 10730
rect 4970 10676 5054 10694
rect 5108 10676 5202 10732
rect 9548 10758 9624 10770
rect 9548 10718 9562 10758
rect 9604 10718 9624 10758
rect 9548 10702 9624 10718
rect 9738 10748 9810 10982
rect 9738 10714 9752 10748
rect 9740 10708 9752 10714
rect 9794 10714 9810 10748
rect 9932 10716 10164 10746
rect 9932 10714 10016 10716
rect 9794 10708 9808 10714
rect 4970 10652 5202 10676
rect 9568 10534 9618 10702
rect 9740 10692 9808 10708
rect 9932 10678 9944 10714
rect 9978 10678 10016 10714
rect 9932 10660 10016 10678
rect 10070 10660 10164 10716
rect 9932 10636 10164 10660
rect 9740 10534 9808 10538
rect 9540 10524 10000 10534
rect 9540 10503 9866 10524
rect 9946 10503 10000 10524
rect 9540 10469 9569 10503
rect 9603 10469 9661 10503
rect 9695 10469 9753 10503
rect 9787 10469 9845 10503
rect 9971 10469 10000 10503
rect 9540 10460 9866 10469
rect 9946 10460 10000 10469
rect 9540 10438 10000 10460
rect 6112 6638 6388 6648
rect 6112 6617 6226 6638
rect 6282 6617 6388 6638
rect 6112 6583 6141 6617
rect 6175 6583 6226 6617
rect 6282 6583 6325 6617
rect 6359 6583 6388 6617
rect 6112 6580 6226 6583
rect 6282 6580 6388 6583
rect 6112 6552 6388 6580
rect 6134 6390 6228 6398
rect 6134 6338 6168 6390
rect 6220 6338 6228 6390
rect 6262 6396 6328 6398
rect 6262 6344 6268 6396
rect 6320 6344 6328 6396
rect 6262 6338 6328 6344
rect 6134 6332 6228 6338
rect 6112 6088 6388 6104
rect 6112 6073 6170 6088
rect 6226 6073 6388 6088
rect 6112 6039 6141 6073
rect 6226 6039 6233 6073
rect 6267 6039 6325 6073
rect 6359 6039 6388 6073
rect 6112 6030 6170 6039
rect 6226 6030 6388 6039
rect 6112 6008 6388 6030
rect 9218 6002 10690 6016
rect 9218 5985 9606 6002
rect 9664 6000 10690 6002
rect 9664 5985 9974 6000
rect 10032 5985 10690 6000
rect 9218 5951 9247 5985
rect 9281 5951 9339 5985
rect 9373 5951 9431 5985
rect 9465 5951 9523 5985
rect 9557 5951 9606 5985
rect 9664 5951 9707 5985
rect 9741 5951 9799 5985
rect 9833 5951 9891 5985
rect 9925 5951 9974 5985
rect 10032 5951 10075 5985
rect 10109 5951 10167 5985
rect 10201 5951 10259 5985
rect 10293 5951 10351 5985
rect 10385 5951 10443 5985
rect 10477 5951 10535 5985
rect 10569 5951 10627 5985
rect 10661 5951 10690 5985
rect 9218 5940 9606 5951
rect 9664 5940 9974 5951
rect 9218 5936 9974 5940
rect 10032 5936 10690 5951
rect 9218 5920 10690 5936
rect 11088 5998 12560 6012
rect 11088 5981 11866 5998
rect 11924 5981 12560 5998
rect 11088 5947 11117 5981
rect 11151 5947 11209 5981
rect 11243 5947 11301 5981
rect 11335 5947 11393 5981
rect 11427 5947 11485 5981
rect 11519 5947 11577 5981
rect 11611 5947 11669 5981
rect 11703 5947 11761 5981
rect 11795 5947 11853 5981
rect 11924 5947 11945 5981
rect 11979 5947 12037 5981
rect 12071 5947 12129 5981
rect 12163 5947 12221 5981
rect 12255 5947 12313 5981
rect 12347 5947 12405 5981
rect 12439 5947 12497 5981
rect 12531 5947 12560 5981
rect 11088 5934 11866 5947
rect 11924 5934 12560 5947
rect 9414 5747 9472 5753
rect 9414 5713 9426 5747
rect 9460 5744 9472 5747
rect 9500 5744 9528 5920
rect 11088 5916 12560 5934
rect 12904 5988 14376 6008
rect 12904 5977 13652 5988
rect 13710 5977 14376 5988
rect 12904 5943 12933 5977
rect 12967 5943 13025 5977
rect 13059 5943 13117 5977
rect 13151 5943 13209 5977
rect 13243 5943 13301 5977
rect 13335 5943 13393 5977
rect 13427 5943 13485 5977
rect 13519 5943 13577 5977
rect 13611 5943 13652 5977
rect 13710 5943 13761 5977
rect 13795 5943 13853 5977
rect 13887 5943 13945 5977
rect 13979 5943 14037 5977
rect 14071 5943 14129 5977
rect 14163 5943 14221 5977
rect 14255 5943 14313 5977
rect 14347 5943 14376 5977
rect 12904 5924 13652 5943
rect 13710 5924 14376 5943
rect 9598 5815 9656 5821
rect 9598 5781 9610 5815
rect 9644 5812 9656 5815
rect 10338 5815 10396 5821
rect 10338 5812 10350 5815
rect 9644 5784 10350 5812
rect 9644 5781 9656 5784
rect 9598 5775 9656 5781
rect 10338 5781 10350 5784
rect 10384 5781 10396 5815
rect 10338 5775 10396 5781
rect 9782 5747 9840 5753
rect 9782 5744 9794 5747
rect 9460 5716 9794 5744
rect 9460 5713 9472 5716
rect 9414 5707 9472 5713
rect 9782 5713 9794 5716
rect 9828 5744 9840 5747
rect 10154 5747 10212 5753
rect 10154 5744 10166 5747
rect 9828 5716 10166 5744
rect 9828 5713 9840 5716
rect 9782 5707 9840 5713
rect 10154 5713 10166 5716
rect 10200 5744 10212 5747
rect 10430 5747 10488 5753
rect 10430 5744 10442 5747
rect 10200 5716 10442 5744
rect 10200 5713 10212 5716
rect 10154 5707 10212 5713
rect 10430 5713 10442 5716
rect 10476 5713 10488 5747
rect 10430 5707 10488 5713
rect 11284 5743 11342 5749
rect 11284 5709 11296 5743
rect 11330 5740 11342 5743
rect 11370 5740 11398 5916
rect 12904 5912 14376 5924
rect 14774 5992 16246 6004
rect 14774 5973 15534 5992
rect 15592 5973 16246 5992
rect 14774 5939 14803 5973
rect 14837 5939 14895 5973
rect 14929 5939 14987 5973
rect 15021 5939 15079 5973
rect 15113 5939 15171 5973
rect 15205 5939 15263 5973
rect 15297 5939 15355 5973
rect 15389 5939 15447 5973
rect 15481 5939 15534 5973
rect 15592 5939 15631 5973
rect 15665 5939 15723 5973
rect 15757 5939 15815 5973
rect 15849 5939 15907 5973
rect 15941 5939 15999 5973
rect 16033 5939 16091 5973
rect 16125 5939 16183 5973
rect 16217 5939 16246 5973
rect 14774 5928 15534 5939
rect 15592 5928 16246 5939
rect 11468 5811 11526 5817
rect 11468 5777 11480 5811
rect 11514 5808 11526 5811
rect 12208 5811 12266 5817
rect 12208 5808 12220 5811
rect 11514 5780 12220 5808
rect 11514 5777 11526 5780
rect 11468 5771 11526 5777
rect 12208 5777 12220 5780
rect 12254 5777 12266 5811
rect 12208 5771 12266 5777
rect 11652 5743 11710 5749
rect 11652 5740 11664 5743
rect 11330 5712 11664 5740
rect 11330 5709 11342 5712
rect 11284 5703 11342 5709
rect 11652 5709 11664 5712
rect 11698 5740 11710 5743
rect 12024 5743 12082 5749
rect 12024 5740 12036 5743
rect 11698 5712 12036 5740
rect 11698 5709 11710 5712
rect 11652 5703 11710 5709
rect 12024 5709 12036 5712
rect 12070 5740 12082 5743
rect 12300 5743 12358 5749
rect 12300 5740 12312 5743
rect 12070 5712 12312 5740
rect 12070 5709 12082 5712
rect 12024 5703 12082 5709
rect 12300 5709 12312 5712
rect 12346 5709 12358 5743
rect 12300 5703 12358 5709
rect 13100 5739 13158 5745
rect 13100 5705 13112 5739
rect 13146 5736 13158 5739
rect 13186 5736 13214 5912
rect 14774 5908 16246 5928
rect 13284 5807 13342 5813
rect 13284 5773 13296 5807
rect 13330 5804 13342 5807
rect 14024 5807 14082 5813
rect 14024 5804 14036 5807
rect 13330 5776 14036 5804
rect 13330 5773 13342 5776
rect 13284 5767 13342 5773
rect 14024 5773 14036 5776
rect 14070 5773 14082 5807
rect 14024 5767 14082 5773
rect 13468 5739 13526 5745
rect 13468 5736 13480 5739
rect 13146 5708 13480 5736
rect 13146 5705 13158 5708
rect 13100 5699 13158 5705
rect 13468 5705 13480 5708
rect 13514 5736 13526 5739
rect 13840 5739 13898 5745
rect 13840 5736 13852 5739
rect 13514 5708 13852 5736
rect 13514 5705 13526 5708
rect 13468 5699 13526 5705
rect 13840 5705 13852 5708
rect 13886 5736 13898 5739
rect 14116 5739 14174 5745
rect 14116 5736 14128 5739
rect 13886 5708 14128 5736
rect 13886 5705 13898 5708
rect 13840 5699 13898 5705
rect 14116 5705 14128 5708
rect 14162 5705 14174 5739
rect 14116 5699 14174 5705
rect 14970 5735 15028 5741
rect 14970 5701 14982 5735
rect 15016 5732 15028 5735
rect 15056 5732 15084 5908
rect 15154 5803 15212 5809
rect 15154 5769 15166 5803
rect 15200 5800 15212 5803
rect 15894 5803 15952 5809
rect 15894 5800 15906 5803
rect 15200 5772 15906 5800
rect 15200 5769 15212 5772
rect 15154 5763 15212 5769
rect 15894 5769 15906 5772
rect 15940 5769 15952 5803
rect 15894 5763 15952 5769
rect 28166 5774 28230 14546
rect 15338 5735 15396 5741
rect 15338 5732 15350 5735
rect 15016 5704 15350 5732
rect 15016 5701 15028 5704
rect 14970 5695 15028 5701
rect 15338 5701 15350 5704
rect 15384 5732 15396 5735
rect 15710 5735 15768 5741
rect 15710 5732 15722 5735
rect 15384 5704 15722 5732
rect 15384 5701 15396 5704
rect 15338 5695 15396 5701
rect 15710 5701 15722 5704
rect 15756 5732 15768 5735
rect 15986 5735 16044 5741
rect 15986 5732 15998 5735
rect 15756 5704 15998 5732
rect 15756 5701 15768 5704
rect 15710 5695 15768 5701
rect 15986 5701 15998 5704
rect 16032 5701 16044 5735
rect 28166 5710 30432 5774
rect 15986 5695 16044 5701
rect 9506 5679 9564 5685
rect 9506 5645 9518 5679
rect 9552 5676 9564 5679
rect 9966 5679 10024 5685
rect 9966 5676 9978 5679
rect 9552 5648 9978 5676
rect 9552 5645 9564 5648
rect 9506 5639 9564 5645
rect 9966 5645 9978 5648
rect 10012 5676 10024 5679
rect 10338 5679 10396 5685
rect 10338 5676 10350 5679
rect 10012 5648 10350 5676
rect 10012 5645 10024 5648
rect 9966 5639 10024 5645
rect 9604 5618 9670 5620
rect 1836 5578 3308 5596
rect 1836 5565 2564 5578
rect 2620 5565 3308 5578
rect 1836 5531 1865 5565
rect 1899 5531 1957 5565
rect 1991 5531 2049 5565
rect 2083 5531 2141 5565
rect 2175 5531 2233 5565
rect 2267 5531 2325 5565
rect 2359 5531 2417 5565
rect 2451 5531 2509 5565
rect 2543 5531 2564 5565
rect 2635 5531 2693 5565
rect 2727 5531 2785 5565
rect 2819 5531 2877 5565
rect 2911 5531 2969 5565
rect 3003 5531 3061 5565
rect 3095 5531 3153 5565
rect 3187 5531 3245 5565
rect 3279 5531 3308 5565
rect 1836 5520 2564 5531
rect 2620 5520 3308 5531
rect 1836 5500 3308 5520
rect 3706 5574 5178 5592
rect 3706 5561 4444 5574
rect 4500 5561 5178 5574
rect 3706 5527 3735 5561
rect 3769 5527 3827 5561
rect 3861 5527 3919 5561
rect 3953 5527 4011 5561
rect 4045 5527 4103 5561
rect 4137 5527 4195 5561
rect 4229 5527 4287 5561
rect 4321 5527 4379 5561
rect 4413 5527 4444 5561
rect 4505 5527 4563 5561
rect 4597 5527 4655 5561
rect 4689 5527 4747 5561
rect 4781 5527 4839 5561
rect 4873 5527 4931 5561
rect 4965 5527 5023 5561
rect 5057 5527 5115 5561
rect 5149 5527 5178 5561
rect 3706 5516 4444 5527
rect 4500 5516 5178 5527
rect 2032 5327 2090 5333
rect 2032 5293 2044 5327
rect 2078 5324 2090 5327
rect 2118 5324 2146 5500
rect 3706 5496 5178 5516
rect 5522 5576 6994 5588
rect 5522 5557 6166 5576
rect 6222 5557 6994 5576
rect 5522 5523 5551 5557
rect 5585 5523 5643 5557
rect 5677 5523 5735 5557
rect 5769 5523 5827 5557
rect 5861 5523 5919 5557
rect 5953 5523 6011 5557
rect 6045 5523 6103 5557
rect 6137 5523 6166 5557
rect 6229 5523 6287 5557
rect 6321 5523 6379 5557
rect 6413 5523 6471 5557
rect 6505 5523 6563 5557
rect 6597 5523 6655 5557
rect 6689 5523 6747 5557
rect 6781 5523 6839 5557
rect 6873 5523 6931 5557
rect 6965 5523 6994 5557
rect 5522 5518 6166 5523
rect 6222 5518 6994 5523
rect 2216 5395 2274 5401
rect 2216 5361 2228 5395
rect 2262 5392 2274 5395
rect 2956 5395 3014 5401
rect 2956 5392 2968 5395
rect 2262 5364 2968 5392
rect 2262 5361 2274 5364
rect 2216 5355 2274 5361
rect 2956 5361 2968 5364
rect 3002 5361 3014 5395
rect 2956 5355 3014 5361
rect 2400 5327 2458 5333
rect 2400 5324 2412 5327
rect 2078 5296 2412 5324
rect 2078 5293 2090 5296
rect 2032 5287 2090 5293
rect 2400 5293 2412 5296
rect 2446 5324 2458 5327
rect 2772 5327 2830 5333
rect 2772 5324 2784 5327
rect 2446 5296 2784 5324
rect 2446 5293 2458 5296
rect 2400 5287 2458 5293
rect 2772 5293 2784 5296
rect 2818 5324 2830 5327
rect 3048 5327 3106 5333
rect 3048 5324 3060 5327
rect 2818 5296 3060 5324
rect 2818 5293 2830 5296
rect 2772 5287 2830 5293
rect 3048 5293 3060 5296
rect 3094 5293 3106 5327
rect 3048 5287 3106 5293
rect 3902 5323 3960 5329
rect 3902 5289 3914 5323
rect 3948 5320 3960 5323
rect 3988 5320 4016 5496
rect 5522 5492 6994 5518
rect 7392 5566 8864 5584
rect 7392 5553 8076 5566
rect 8132 5553 8864 5566
rect 9604 5566 9610 5618
rect 9662 5566 9670 5618
rect 9604 5562 9670 5566
rect 7392 5519 7421 5553
rect 7455 5519 7513 5553
rect 7547 5519 7605 5553
rect 7639 5519 7697 5553
rect 7731 5519 7789 5553
rect 7823 5519 7881 5553
rect 7915 5519 7973 5553
rect 8007 5519 8065 5553
rect 8132 5519 8157 5553
rect 8191 5519 8249 5553
rect 8283 5519 8341 5553
rect 8375 5519 8433 5553
rect 8467 5519 8525 5553
rect 8559 5519 8617 5553
rect 8651 5519 8709 5553
rect 8743 5519 8801 5553
rect 8835 5519 8864 5553
rect 7392 5508 8076 5519
rect 8132 5508 8864 5519
rect 4086 5391 4144 5397
rect 4086 5357 4098 5391
rect 4132 5388 4144 5391
rect 4826 5391 4884 5397
rect 4826 5388 4838 5391
rect 4132 5360 4838 5388
rect 4132 5357 4144 5360
rect 4086 5351 4144 5357
rect 4826 5357 4838 5360
rect 4872 5357 4884 5391
rect 4826 5351 4884 5357
rect 4270 5323 4328 5329
rect 4270 5320 4282 5323
rect 3948 5292 4282 5320
rect 3948 5289 3960 5292
rect 3902 5283 3960 5289
rect 4270 5289 4282 5292
rect 4316 5320 4328 5323
rect 4642 5323 4700 5329
rect 4642 5320 4654 5323
rect 4316 5292 4654 5320
rect 4316 5289 4328 5292
rect 4270 5283 4328 5289
rect 4642 5289 4654 5292
rect 4688 5320 4700 5323
rect 4918 5323 4976 5329
rect 4918 5320 4930 5323
rect 4688 5292 4930 5320
rect 4688 5289 4700 5292
rect 4642 5283 4700 5289
rect 4918 5289 4930 5292
rect 4964 5289 4976 5323
rect 4918 5283 4976 5289
rect 5718 5319 5776 5325
rect 5718 5285 5730 5319
rect 5764 5316 5776 5319
rect 5804 5316 5832 5492
rect 7392 5488 8864 5508
rect 5902 5387 5960 5393
rect 5902 5353 5914 5387
rect 5948 5384 5960 5387
rect 6642 5387 6700 5393
rect 6642 5384 6654 5387
rect 5948 5356 6654 5384
rect 5948 5353 5960 5356
rect 5902 5347 5960 5353
rect 6642 5353 6654 5356
rect 6688 5353 6700 5387
rect 6642 5347 6700 5353
rect 6086 5319 6144 5325
rect 6086 5316 6098 5319
rect 5764 5288 6098 5316
rect 5764 5285 5776 5288
rect 5718 5279 5776 5285
rect 6086 5285 6098 5288
rect 6132 5316 6144 5319
rect 6458 5319 6516 5325
rect 6458 5316 6470 5319
rect 6132 5288 6470 5316
rect 6132 5285 6144 5288
rect 6086 5279 6144 5285
rect 6458 5285 6470 5288
rect 6504 5316 6516 5319
rect 6734 5319 6792 5325
rect 6734 5316 6746 5319
rect 6504 5288 6746 5316
rect 6504 5285 6516 5288
rect 6458 5279 6516 5285
rect 6734 5285 6746 5288
rect 6780 5285 6792 5319
rect 6734 5279 6792 5285
rect 7588 5315 7646 5321
rect 7588 5281 7600 5315
rect 7634 5312 7646 5315
rect 7674 5312 7702 5488
rect 10060 5472 10088 5648
rect 10338 5645 10350 5648
rect 10384 5645 10396 5679
rect 10338 5639 10396 5645
rect 11376 5675 11434 5681
rect 11376 5641 11388 5675
rect 11422 5672 11434 5675
rect 11836 5675 11894 5681
rect 11836 5672 11848 5675
rect 11422 5644 11848 5672
rect 11422 5641 11434 5644
rect 11376 5635 11434 5641
rect 11836 5641 11848 5644
rect 11882 5672 11894 5675
rect 12208 5675 12266 5681
rect 12208 5672 12220 5675
rect 11882 5644 12220 5672
rect 11882 5641 11894 5644
rect 11836 5635 11894 5641
rect 10612 5606 10672 5630
rect 10612 5570 10626 5606
rect 10666 5604 10672 5606
rect 11472 5608 11532 5614
rect 11472 5604 11486 5608
rect 10666 5574 11486 5604
rect 11520 5574 11532 5608
rect 10666 5570 11532 5574
rect 10612 5566 11532 5570
rect 10612 5554 10672 5566
rect 11472 5552 11532 5566
rect 9218 5452 10690 5472
rect 11930 5468 11958 5644
rect 12208 5641 12220 5644
rect 12254 5641 12266 5675
rect 12208 5635 12266 5641
rect 13192 5671 13250 5677
rect 13192 5637 13204 5671
rect 13238 5668 13250 5671
rect 13652 5671 13710 5677
rect 13652 5668 13664 5671
rect 13238 5640 13664 5668
rect 13238 5637 13250 5640
rect 13192 5631 13250 5637
rect 13652 5637 13664 5640
rect 13698 5668 13710 5671
rect 14024 5671 14082 5677
rect 14024 5668 14036 5671
rect 13698 5640 14036 5668
rect 13698 5637 13710 5640
rect 13652 5631 13710 5637
rect 12492 5602 12544 5626
rect 13288 5604 13348 5612
rect 13288 5602 13302 5604
rect 12492 5568 12502 5602
rect 12538 5570 13302 5602
rect 13336 5570 13348 5604
rect 12538 5568 13348 5570
rect 12492 5564 13348 5568
rect 12492 5550 12544 5564
rect 9218 5441 10414 5452
rect 10470 5441 10690 5452
rect 9218 5407 9247 5441
rect 9281 5407 9339 5441
rect 9373 5407 9431 5441
rect 9465 5407 9523 5441
rect 9557 5407 9615 5441
rect 9649 5407 9707 5441
rect 9741 5407 9799 5441
rect 9833 5407 9891 5441
rect 9925 5407 9983 5441
rect 10017 5407 10075 5441
rect 10109 5407 10167 5441
rect 10201 5407 10259 5441
rect 10293 5407 10351 5441
rect 10385 5407 10414 5441
rect 10477 5407 10535 5441
rect 10569 5407 10627 5441
rect 10661 5407 10690 5441
rect 9218 5394 10414 5407
rect 10470 5394 10690 5407
rect 7772 5383 7830 5389
rect 7772 5349 7784 5383
rect 7818 5380 7830 5383
rect 8512 5383 8570 5389
rect 8512 5380 8524 5383
rect 7818 5352 8524 5380
rect 7818 5349 7830 5352
rect 7772 5343 7830 5349
rect 8512 5349 8524 5352
rect 8558 5349 8570 5383
rect 9218 5376 10690 5394
rect 11088 5456 12560 5468
rect 13746 5464 13774 5640
rect 14024 5637 14036 5640
rect 14070 5637 14082 5671
rect 14024 5631 14082 5637
rect 15062 5667 15120 5673
rect 15062 5633 15074 5667
rect 15108 5664 15120 5667
rect 15522 5667 15580 5673
rect 15522 5664 15534 5667
rect 15108 5636 15534 5664
rect 15108 5633 15120 5636
rect 15062 5627 15120 5633
rect 15522 5633 15534 5636
rect 15568 5664 15580 5667
rect 15894 5667 15952 5673
rect 15894 5664 15906 5667
rect 15568 5636 15906 5664
rect 15568 5633 15580 5636
rect 15522 5627 15580 5633
rect 14298 5598 14358 5622
rect 14298 5562 14312 5598
rect 14352 5596 14358 5598
rect 15158 5600 15218 5606
rect 15158 5596 15172 5600
rect 14352 5566 15172 5596
rect 15206 5566 15218 5600
rect 14352 5562 15218 5566
rect 14298 5558 15218 5562
rect 14298 5546 14358 5558
rect 15158 5544 15218 5558
rect 11088 5437 11370 5456
rect 11428 5437 12560 5456
rect 11088 5403 11117 5437
rect 11151 5403 11209 5437
rect 11243 5403 11301 5437
rect 11335 5403 11370 5437
rect 11428 5403 11485 5437
rect 11519 5403 11577 5437
rect 11611 5403 11669 5437
rect 11703 5403 11761 5437
rect 11795 5403 11853 5437
rect 11887 5403 11945 5437
rect 11979 5403 12037 5437
rect 12071 5403 12129 5437
rect 12163 5403 12221 5437
rect 12255 5403 12313 5437
rect 12347 5403 12405 5437
rect 12439 5403 12497 5437
rect 12531 5403 12560 5437
rect 11088 5392 11370 5403
rect 11428 5392 12560 5403
rect 11088 5372 12560 5392
rect 12904 5450 14376 5464
rect 15616 5460 15644 5636
rect 15894 5633 15906 5636
rect 15940 5633 15952 5667
rect 15894 5627 15952 5633
rect 16166 5600 16228 5608
rect 16166 5564 16182 5600
rect 16216 5596 16228 5600
rect 16216 5564 16722 5596
rect 16166 5554 16228 5564
rect 12904 5433 14072 5450
rect 14130 5433 14376 5450
rect 12904 5399 12933 5433
rect 12967 5399 13025 5433
rect 13059 5399 13117 5433
rect 13151 5399 13209 5433
rect 13243 5399 13301 5433
rect 13335 5399 13393 5433
rect 13427 5399 13485 5433
rect 13519 5399 13577 5433
rect 13611 5399 13669 5433
rect 13703 5399 13761 5433
rect 13795 5399 13853 5433
rect 13887 5399 13945 5433
rect 13979 5399 14037 5433
rect 14071 5399 14072 5433
rect 14163 5399 14221 5433
rect 14255 5399 14313 5433
rect 14347 5399 14376 5433
rect 12904 5386 14072 5399
rect 14130 5386 14376 5399
rect 12904 5368 14376 5386
rect 14774 5442 16246 5460
rect 14774 5429 14992 5442
rect 15050 5429 16246 5442
rect 14774 5395 14803 5429
rect 14837 5395 14895 5429
rect 14929 5395 14987 5429
rect 15050 5395 15079 5429
rect 15113 5395 15171 5429
rect 15205 5395 15263 5429
rect 15297 5395 15355 5429
rect 15389 5395 15447 5429
rect 15481 5395 15539 5429
rect 15573 5395 15631 5429
rect 15665 5395 15723 5429
rect 15757 5395 15815 5429
rect 15849 5395 15907 5429
rect 15941 5395 15999 5429
rect 16033 5395 16091 5429
rect 16125 5395 16183 5429
rect 16217 5395 16246 5429
rect 14774 5378 14992 5395
rect 15050 5378 16246 5395
rect 14774 5364 16246 5378
rect 8512 5343 8570 5349
rect 7956 5315 8014 5321
rect 7956 5312 7968 5315
rect 7634 5284 7968 5312
rect 7634 5281 7646 5284
rect 7588 5275 7646 5281
rect 7956 5281 7968 5284
rect 8002 5312 8014 5315
rect 8328 5315 8386 5321
rect 8328 5312 8340 5315
rect 8002 5284 8340 5312
rect 8002 5281 8014 5284
rect 7956 5275 8014 5281
rect 8328 5281 8340 5284
rect 8374 5312 8386 5315
rect 8604 5315 8662 5321
rect 8604 5312 8616 5315
rect 8374 5284 8616 5312
rect 8374 5281 8386 5284
rect 8328 5275 8386 5281
rect 8604 5281 8616 5284
rect 8650 5281 8662 5315
rect 8604 5275 8662 5281
rect 16690 5302 16722 5564
rect 16690 5270 17232 5302
rect 2124 5259 2182 5265
rect 2124 5225 2136 5259
rect 2170 5256 2182 5259
rect 2584 5259 2642 5265
rect 2584 5256 2596 5259
rect 2170 5228 2596 5256
rect 2170 5225 2182 5228
rect 2124 5219 2182 5225
rect 2584 5225 2596 5228
rect 2630 5256 2642 5259
rect 2956 5259 3014 5265
rect 2956 5256 2968 5259
rect 2630 5228 2968 5256
rect 2630 5225 2642 5228
rect 2584 5219 2642 5225
rect 2222 5198 2288 5200
rect 2222 5146 2228 5198
rect 2280 5146 2288 5198
rect 2222 5142 2288 5146
rect 2678 5052 2706 5228
rect 2956 5225 2968 5228
rect 3002 5225 3014 5259
rect 2956 5219 3014 5225
rect 3994 5255 4052 5261
rect 3994 5221 4006 5255
rect 4040 5252 4052 5255
rect 4454 5255 4512 5261
rect 4454 5252 4466 5255
rect 4040 5224 4466 5252
rect 4040 5221 4052 5224
rect 3994 5215 4052 5221
rect 4454 5221 4466 5224
rect 4500 5252 4512 5255
rect 4826 5255 4884 5261
rect 4826 5252 4838 5255
rect 4500 5224 4838 5252
rect 4500 5221 4512 5224
rect 4454 5215 4512 5221
rect 3230 5186 3290 5210
rect 3230 5150 3244 5186
rect 3284 5184 3290 5186
rect 4090 5188 4150 5194
rect 4090 5184 4104 5188
rect 3284 5154 4104 5184
rect 4138 5154 4150 5188
rect 3284 5150 4150 5154
rect 3230 5146 4150 5150
rect 3230 5134 3290 5146
rect 4090 5132 4150 5146
rect 1836 5040 3308 5052
rect 4548 5048 4576 5224
rect 4826 5221 4838 5224
rect 4872 5221 4884 5255
rect 4826 5215 4884 5221
rect 5810 5251 5868 5257
rect 5100 5182 5164 5220
rect 5810 5217 5822 5251
rect 5856 5248 5868 5251
rect 6270 5251 6328 5257
rect 6270 5248 6282 5251
rect 5856 5220 6282 5248
rect 5856 5217 5868 5220
rect 5810 5211 5868 5217
rect 6270 5217 6282 5220
rect 6316 5248 6328 5251
rect 6642 5251 6700 5257
rect 6642 5248 6654 5251
rect 6316 5220 6654 5248
rect 6316 5217 6328 5220
rect 6270 5211 6328 5217
rect 5906 5184 5966 5192
rect 5906 5182 5920 5184
rect 5100 5144 5120 5182
rect 5156 5150 5920 5182
rect 5954 5150 5966 5184
rect 5156 5144 5966 5150
rect 5100 5124 5164 5144
rect 1836 5021 2584 5040
rect 2640 5021 3308 5040
rect 1836 4987 1865 5021
rect 1899 4987 1957 5021
rect 1991 4987 2049 5021
rect 2083 4987 2141 5021
rect 2175 4987 2233 5021
rect 2267 4987 2325 5021
rect 2359 4987 2417 5021
rect 2451 4987 2509 5021
rect 2543 4987 2584 5021
rect 2640 4987 2693 5021
rect 2727 4987 2785 5021
rect 2819 4987 2877 5021
rect 2911 4987 2969 5021
rect 3003 4987 3061 5021
rect 3095 4987 3153 5021
rect 3187 4987 3245 5021
rect 3279 4987 3308 5021
rect 1836 4982 2584 4987
rect 2640 4982 3308 4987
rect 1836 4956 3308 4982
rect 3706 5032 5178 5048
rect 6364 5044 6392 5220
rect 6642 5217 6654 5220
rect 6688 5217 6700 5251
rect 6642 5211 6700 5217
rect 7680 5247 7738 5253
rect 7680 5213 7692 5247
rect 7726 5244 7738 5247
rect 8140 5247 8198 5253
rect 8140 5244 8152 5247
rect 7726 5216 8152 5244
rect 7726 5213 7738 5216
rect 7680 5207 7738 5213
rect 8140 5213 8152 5216
rect 8186 5244 8198 5247
rect 8512 5247 8570 5253
rect 8512 5244 8524 5247
rect 8186 5216 8524 5244
rect 8186 5213 8198 5216
rect 8140 5207 8198 5213
rect 6916 5178 6976 5202
rect 6916 5142 6930 5178
rect 6970 5176 6976 5178
rect 7776 5180 7836 5186
rect 7776 5176 7790 5180
rect 6970 5146 7790 5176
rect 7824 5146 7836 5180
rect 6970 5142 7836 5146
rect 6916 5138 7836 5142
rect 6916 5126 6976 5138
rect 7776 5124 7836 5138
rect 3706 5017 4444 5032
rect 4500 5017 5178 5032
rect 3706 4983 3735 5017
rect 3769 4983 3827 5017
rect 3861 4983 3919 5017
rect 3953 4983 4011 5017
rect 4045 4983 4103 5017
rect 4137 4983 4195 5017
rect 4229 4983 4287 5017
rect 4321 4983 4379 5017
rect 4413 4983 4444 5017
rect 4505 4983 4563 5017
rect 4597 4983 4655 5017
rect 4689 4983 4747 5017
rect 4781 4983 4839 5017
rect 4873 4983 4931 5017
rect 4965 4983 5023 5017
rect 5057 4983 5115 5017
rect 5149 4983 5178 5017
rect 3706 4974 4444 4983
rect 4500 4974 5178 4983
rect 3706 4952 5178 4974
rect 5522 5028 6994 5044
rect 8234 5040 8262 5216
rect 8512 5213 8524 5216
rect 8558 5213 8570 5247
rect 8512 5207 8570 5213
rect 9106 5210 16590 5242
rect 8784 5180 8846 5188
rect 8784 5144 8800 5180
rect 8834 5176 8846 5180
rect 9106 5176 9138 5210
rect 8834 5144 9138 5176
rect 8784 5134 8846 5144
rect 9246 5120 10718 5142
rect 9246 5111 9388 5120
rect 9444 5111 10718 5120
rect 9246 5077 9275 5111
rect 9309 5077 9367 5111
rect 9444 5077 9459 5111
rect 9493 5077 9551 5111
rect 9585 5077 9643 5111
rect 9677 5077 9735 5111
rect 9769 5077 9827 5111
rect 9861 5077 9919 5111
rect 9953 5077 10011 5111
rect 10045 5077 10103 5111
rect 10137 5077 10195 5111
rect 10229 5077 10287 5111
rect 10321 5077 10379 5111
rect 10413 5077 10471 5111
rect 10505 5077 10563 5111
rect 10597 5077 10655 5111
rect 10689 5077 10718 5111
rect 9246 5062 9388 5077
rect 9444 5062 10718 5077
rect 9246 5046 10718 5062
rect 11116 5120 12588 5138
rect 11116 5107 12276 5120
rect 12334 5107 12588 5120
rect 11116 5073 11145 5107
rect 11179 5073 11237 5107
rect 11271 5073 11329 5107
rect 11363 5073 11421 5107
rect 11455 5073 11513 5107
rect 11547 5073 11605 5107
rect 11639 5073 11697 5107
rect 11731 5073 11789 5107
rect 11823 5073 11881 5107
rect 11915 5073 11973 5107
rect 12007 5073 12065 5107
rect 12099 5073 12157 5107
rect 12191 5073 12249 5107
rect 12334 5073 12341 5107
rect 12375 5073 12433 5107
rect 12467 5073 12525 5107
rect 12559 5073 12588 5107
rect 11116 5056 12276 5073
rect 12334 5056 12588 5073
rect 5522 5013 6148 5028
rect 6204 5013 6994 5028
rect 5522 4979 5551 5013
rect 5585 4979 5643 5013
rect 5677 4979 5735 5013
rect 5769 4979 5827 5013
rect 5861 4979 5919 5013
rect 5953 4979 6011 5013
rect 6045 4979 6103 5013
rect 6137 4979 6148 5013
rect 6229 4979 6287 5013
rect 6321 4979 6379 5013
rect 6413 4979 6471 5013
rect 6505 4979 6563 5013
rect 6597 4979 6655 5013
rect 6689 4979 6747 5013
rect 6781 4979 6839 5013
rect 6873 4979 6931 5013
rect 6965 4979 6994 5013
rect 5522 4970 6148 4979
rect 6204 4970 6994 4979
rect 5522 4948 6994 4970
rect 7392 5020 8864 5040
rect 7392 5009 8064 5020
rect 8120 5009 8864 5020
rect 7392 4975 7421 5009
rect 7455 4975 7513 5009
rect 7547 4975 7605 5009
rect 7639 4975 7697 5009
rect 7731 4975 7789 5009
rect 7823 4975 7881 5009
rect 7915 4975 7973 5009
rect 8007 4975 8064 5009
rect 8120 4975 8157 5009
rect 8191 4975 8249 5009
rect 8283 4975 8341 5009
rect 8375 4975 8433 5009
rect 8467 4975 8525 5009
rect 8559 4975 8617 5009
rect 8651 4975 8709 5009
rect 8743 4975 8801 5009
rect 8835 4975 8864 5009
rect 7392 4962 8064 4975
rect 8120 4962 8864 4975
rect 7392 4944 8864 4962
rect 9442 4873 9500 4879
rect 9442 4839 9454 4873
rect 9488 4870 9500 4873
rect 9528 4870 9556 5046
rect 11116 5042 12588 5056
rect 12932 5116 14404 5134
rect 12932 5103 13130 5116
rect 13188 5103 14404 5116
rect 12932 5069 12961 5103
rect 12995 5069 13053 5103
rect 13087 5069 13130 5103
rect 13188 5069 13237 5103
rect 13271 5069 13329 5103
rect 13363 5069 13421 5103
rect 13455 5069 13513 5103
rect 13547 5069 13605 5103
rect 13639 5069 13697 5103
rect 13731 5069 13789 5103
rect 13823 5069 13881 5103
rect 13915 5069 13973 5103
rect 14007 5069 14065 5103
rect 14099 5069 14157 5103
rect 14191 5069 14249 5103
rect 14283 5069 14341 5103
rect 14375 5069 14404 5103
rect 12932 5052 13130 5069
rect 13188 5052 14404 5069
rect 9626 4941 9684 4947
rect 9626 4907 9638 4941
rect 9672 4938 9684 4941
rect 10366 4941 10424 4947
rect 10366 4938 10378 4941
rect 9672 4910 10378 4938
rect 9672 4907 9684 4910
rect 9626 4901 9684 4907
rect 10366 4907 10378 4910
rect 10412 4907 10424 4941
rect 10366 4901 10424 4907
rect 9810 4873 9868 4879
rect 9810 4870 9822 4873
rect 9488 4842 9822 4870
rect 9488 4839 9500 4842
rect 9442 4833 9500 4839
rect 9810 4839 9822 4842
rect 9856 4870 9868 4873
rect 10182 4873 10240 4879
rect 10182 4870 10194 4873
rect 9856 4842 10194 4870
rect 9856 4839 9868 4842
rect 9810 4833 9868 4839
rect 10182 4839 10194 4842
rect 10228 4870 10240 4873
rect 10458 4873 10516 4879
rect 10458 4870 10470 4873
rect 10228 4842 10470 4870
rect 10228 4839 10240 4842
rect 10182 4833 10240 4839
rect 10458 4839 10470 4842
rect 10504 4839 10516 4873
rect 10458 4833 10516 4839
rect 11312 4869 11370 4875
rect 11312 4835 11324 4869
rect 11358 4866 11370 4869
rect 11398 4866 11426 5042
rect 12932 5038 14404 5052
rect 14802 5114 16274 5130
rect 14802 5099 15922 5114
rect 15980 5099 16274 5114
rect 14802 5065 14831 5099
rect 14865 5065 14923 5099
rect 14957 5065 15015 5099
rect 15049 5065 15107 5099
rect 15141 5065 15199 5099
rect 15233 5065 15291 5099
rect 15325 5065 15383 5099
rect 15417 5065 15475 5099
rect 15509 5065 15567 5099
rect 15601 5065 15659 5099
rect 15693 5065 15751 5099
rect 15785 5065 15843 5099
rect 15877 5065 15922 5099
rect 15980 5065 16027 5099
rect 16061 5065 16119 5099
rect 16153 5065 16211 5099
rect 16245 5065 16274 5099
rect 16521 5108 16590 5210
rect 17098 5222 17148 5242
rect 17098 5188 17108 5222
rect 17142 5188 17148 5222
rect 17098 5134 17148 5188
rect 17178 5194 17232 5270
rect 17178 5160 17190 5194
rect 17224 5160 17232 5194
rect 16926 5108 16980 5120
rect 16521 5070 16932 5108
rect 16970 5070 17072 5108
rect 14802 5050 15922 5065
rect 15980 5050 16274 5065
rect 16926 5054 16980 5070
rect 11496 4937 11554 4943
rect 11496 4903 11508 4937
rect 11542 4934 11554 4937
rect 12236 4937 12294 4943
rect 12236 4934 12248 4937
rect 11542 4906 12248 4934
rect 11542 4903 11554 4906
rect 11496 4897 11554 4903
rect 12236 4903 12248 4906
rect 12282 4903 12294 4937
rect 12236 4897 12294 4903
rect 11680 4869 11738 4875
rect 11680 4866 11692 4869
rect 11358 4838 11692 4866
rect 11358 4835 11370 4838
rect 11312 4829 11370 4835
rect 11680 4835 11692 4838
rect 11726 4866 11738 4869
rect 12052 4869 12110 4875
rect 12052 4866 12064 4869
rect 11726 4838 12064 4866
rect 11726 4835 11738 4838
rect 11680 4829 11738 4835
rect 12052 4835 12064 4838
rect 12098 4866 12110 4869
rect 12328 4869 12386 4875
rect 12328 4866 12340 4869
rect 12098 4838 12340 4866
rect 12098 4835 12110 4838
rect 12052 4829 12110 4835
rect 12328 4835 12340 4838
rect 12374 4835 12386 4869
rect 12328 4829 12386 4835
rect 13128 4865 13186 4871
rect 13128 4831 13140 4865
rect 13174 4862 13186 4865
rect 13214 4862 13242 5038
rect 14802 5034 16274 5050
rect 13312 4933 13370 4939
rect 13312 4899 13324 4933
rect 13358 4930 13370 4933
rect 14052 4933 14110 4939
rect 14052 4930 14064 4933
rect 13358 4902 14064 4930
rect 13358 4899 13370 4902
rect 13312 4893 13370 4899
rect 14052 4899 14064 4902
rect 14098 4899 14110 4933
rect 14052 4893 14110 4899
rect 13496 4865 13554 4871
rect 13496 4862 13508 4865
rect 13174 4834 13508 4862
rect 13174 4831 13186 4834
rect 13128 4825 13186 4831
rect 13496 4831 13508 4834
rect 13542 4862 13554 4865
rect 13868 4865 13926 4871
rect 13868 4862 13880 4865
rect 13542 4834 13880 4862
rect 13542 4831 13554 4834
rect 13496 4825 13554 4831
rect 13868 4831 13880 4834
rect 13914 4862 13926 4865
rect 14144 4865 14202 4871
rect 14144 4862 14156 4865
rect 13914 4834 14156 4862
rect 13914 4831 13926 4834
rect 13868 4825 13926 4831
rect 14144 4831 14156 4834
rect 14190 4831 14202 4865
rect 14144 4825 14202 4831
rect 14998 4861 15056 4867
rect 14998 4827 15010 4861
rect 15044 4858 15056 4861
rect 15084 4858 15112 5034
rect 17108 5024 17140 5134
rect 17178 5114 17232 5160
rect 17178 5110 17216 5114
rect 16558 4992 17140 5024
rect 17546 5050 17612 5098
rect 17546 4998 17556 5050
rect 17608 4998 17612 5050
rect 15182 4929 15240 4935
rect 15182 4895 15194 4929
rect 15228 4926 15240 4929
rect 15922 4929 15980 4935
rect 15922 4926 15934 4929
rect 15228 4898 15934 4926
rect 15228 4895 15240 4898
rect 15182 4889 15240 4895
rect 15922 4895 15934 4898
rect 15968 4895 15980 4929
rect 15922 4889 15980 4895
rect 15366 4861 15424 4867
rect 15366 4858 15378 4861
rect 15044 4830 15378 4858
rect 15044 4827 15056 4830
rect 14998 4821 15056 4827
rect 15366 4827 15378 4830
rect 15412 4858 15424 4861
rect 15738 4861 15796 4867
rect 15738 4858 15750 4861
rect 15412 4830 15750 4858
rect 15412 4827 15424 4830
rect 15366 4821 15424 4827
rect 15738 4827 15750 4830
rect 15784 4858 15796 4861
rect 16014 4861 16072 4867
rect 16014 4858 16026 4861
rect 15784 4830 16026 4858
rect 15784 4827 15796 4830
rect 15738 4821 15796 4827
rect 16014 4827 16026 4830
rect 16060 4827 16072 4861
rect 16014 4821 16072 4827
rect 9534 4805 9592 4811
rect 9534 4771 9546 4805
rect 9580 4802 9592 4805
rect 9994 4805 10052 4811
rect 9994 4802 10006 4805
rect 9580 4774 10006 4802
rect 9580 4771 9592 4774
rect 9534 4765 9592 4771
rect 9994 4771 10006 4774
rect 10040 4802 10052 4805
rect 10366 4805 10424 4811
rect 10366 4802 10378 4805
rect 10040 4774 10378 4802
rect 10040 4771 10052 4774
rect 9994 4765 10052 4771
rect 9632 4744 9698 4746
rect 9632 4692 9638 4744
rect 9690 4692 9698 4744
rect 9632 4688 9698 4692
rect 10088 4598 10116 4774
rect 10366 4771 10378 4774
rect 10412 4771 10424 4805
rect 10366 4765 10424 4771
rect 11404 4801 11462 4807
rect 11404 4767 11416 4801
rect 11450 4798 11462 4801
rect 11864 4801 11922 4807
rect 11864 4798 11876 4801
rect 11450 4770 11876 4798
rect 11450 4767 11462 4770
rect 11404 4761 11462 4767
rect 11864 4767 11876 4770
rect 11910 4798 11922 4801
rect 12236 4801 12294 4807
rect 12236 4798 12248 4801
rect 11910 4770 12248 4798
rect 11910 4767 11922 4770
rect 11864 4761 11922 4767
rect 10640 4732 10700 4756
rect 10640 4696 10654 4732
rect 10694 4730 10700 4732
rect 11500 4734 11560 4740
rect 11500 4730 11514 4734
rect 10694 4700 11514 4730
rect 11548 4700 11560 4734
rect 10694 4696 11560 4700
rect 10640 4692 11560 4696
rect 10640 4680 10700 4692
rect 11500 4678 11560 4692
rect 9246 4580 10718 4598
rect 11958 4594 11986 4770
rect 12236 4767 12248 4770
rect 12282 4767 12294 4801
rect 12236 4761 12294 4767
rect 13220 4797 13278 4803
rect 13220 4763 13232 4797
rect 13266 4794 13278 4797
rect 13680 4797 13738 4803
rect 13680 4794 13692 4797
rect 13266 4766 13692 4794
rect 13266 4763 13278 4766
rect 13220 4757 13278 4763
rect 13680 4763 13692 4766
rect 13726 4794 13738 4797
rect 14052 4797 14110 4803
rect 14052 4794 14064 4797
rect 13726 4766 14064 4794
rect 13726 4763 13738 4766
rect 13680 4757 13738 4763
rect 12518 4728 12572 4742
rect 13316 4730 13376 4738
rect 13316 4728 13330 4730
rect 12518 4718 13330 4728
rect 12518 4684 12530 4718
rect 12564 4696 13330 4718
rect 13364 4696 13376 4730
rect 12564 4690 13376 4696
rect 12564 4684 12572 4690
rect 12518 4670 12572 4684
rect 9246 4567 9988 4580
rect 10044 4567 10718 4580
rect 9246 4533 9275 4567
rect 9309 4533 9367 4567
rect 9401 4533 9459 4567
rect 9493 4533 9551 4567
rect 9585 4566 9643 4567
rect 9677 4566 9735 4567
rect 9585 4533 9640 4566
rect 9692 4533 9735 4566
rect 9769 4533 9827 4567
rect 9861 4533 9919 4567
rect 9953 4533 9988 4567
rect 10045 4533 10103 4567
rect 10137 4533 10195 4567
rect 10229 4533 10287 4567
rect 10321 4533 10379 4567
rect 10413 4533 10471 4567
rect 10505 4533 10563 4567
rect 10597 4533 10655 4567
rect 10689 4533 10718 4567
rect 9246 4512 9640 4533
rect 9692 4522 9988 4533
rect 10044 4522 10718 4533
rect 9692 4512 10718 4522
rect 9246 4502 10718 4512
rect 11116 4578 12588 4594
rect 13774 4590 13802 4766
rect 14052 4763 14064 4766
rect 14098 4763 14110 4797
rect 14052 4757 14110 4763
rect 15090 4793 15148 4799
rect 15090 4759 15102 4793
rect 15136 4790 15148 4793
rect 15550 4793 15608 4799
rect 15550 4790 15562 4793
rect 15136 4762 15562 4790
rect 15136 4759 15148 4762
rect 15090 4753 15148 4759
rect 15550 4759 15562 4762
rect 15596 4790 15608 4793
rect 15922 4793 15980 4799
rect 15922 4790 15934 4793
rect 15596 4762 15934 4790
rect 15596 4759 15608 4762
rect 15550 4753 15608 4759
rect 14326 4724 14386 4748
rect 14326 4688 14340 4724
rect 14380 4722 14386 4724
rect 15186 4726 15246 4732
rect 15186 4722 15200 4726
rect 14380 4692 15200 4722
rect 15234 4692 15246 4726
rect 14380 4688 15246 4692
rect 14326 4684 15246 4688
rect 14326 4672 14386 4684
rect 15186 4670 15246 4684
rect 11116 4563 11894 4578
rect 11952 4563 12588 4578
rect 11116 4529 11145 4563
rect 11179 4529 11237 4563
rect 11271 4529 11329 4563
rect 11363 4529 11421 4563
rect 11455 4529 11513 4563
rect 11547 4529 11605 4563
rect 11639 4529 11697 4563
rect 11731 4529 11789 4563
rect 11823 4529 11881 4563
rect 11952 4529 11973 4563
rect 12007 4529 12065 4563
rect 12099 4529 12157 4563
rect 12191 4529 12249 4563
rect 12283 4529 12341 4563
rect 12375 4529 12433 4563
rect 12467 4529 12525 4563
rect 12559 4529 12588 4563
rect 11116 4514 11894 4529
rect 11952 4514 12588 4529
rect 11116 4498 12588 4514
rect 12932 4574 14404 4590
rect 15644 4586 15672 4762
rect 15922 4759 15934 4762
rect 15968 4759 15980 4793
rect 15922 4753 15980 4759
rect 16194 4726 16256 4734
rect 16194 4690 16210 4726
rect 16244 4722 16256 4726
rect 16558 4722 16590 4992
rect 17546 4944 17612 4998
rect 16244 4690 16590 4722
rect 16194 4680 16256 4690
rect 12932 4559 13698 4574
rect 13756 4559 14404 4574
rect 12932 4525 12961 4559
rect 12995 4525 13053 4559
rect 13087 4525 13145 4559
rect 13179 4525 13237 4559
rect 13271 4525 13329 4559
rect 13363 4525 13421 4559
rect 13455 4525 13513 4559
rect 13547 4525 13605 4559
rect 13639 4525 13697 4559
rect 13756 4525 13789 4559
rect 13823 4525 13881 4559
rect 13915 4525 13973 4559
rect 14007 4525 14065 4559
rect 14099 4525 14157 4559
rect 14191 4525 14249 4559
rect 14283 4525 14341 4559
rect 14375 4525 14404 4559
rect 12932 4510 13698 4525
rect 13756 4510 14404 4525
rect 12932 4494 14404 4510
rect 14802 4566 16274 4586
rect 14802 4555 15628 4566
rect 15686 4555 16274 4566
rect 14802 4521 14831 4555
rect 14865 4521 14923 4555
rect 14957 4521 15015 4555
rect 15049 4521 15107 4555
rect 15141 4521 15199 4555
rect 15233 4521 15291 4555
rect 15325 4521 15383 4555
rect 15417 4521 15475 4555
rect 15509 4521 15567 4555
rect 15601 4521 15628 4555
rect 15693 4521 15751 4555
rect 15785 4521 15843 4555
rect 15877 4521 15935 4555
rect 15969 4521 16027 4555
rect 16061 4521 16119 4555
rect 16153 4521 16211 4555
rect 16245 4521 16274 4555
rect 14802 4502 15628 4521
rect 15686 4502 16274 4521
rect 14802 4490 16274 4502
rect 6104 3130 6198 3138
rect 6104 3078 6138 3130
rect 6190 3078 6198 3130
rect 6232 3136 6298 3138
rect 6232 3084 6238 3136
rect 6290 3084 6298 3136
rect 6232 3078 6298 3084
rect 6104 3072 6198 3078
rect 1806 2318 3278 2336
rect 1806 2305 2604 2318
rect 2660 2305 3278 2318
rect 1806 2271 1835 2305
rect 1869 2271 1927 2305
rect 1961 2271 2019 2305
rect 2053 2271 2111 2305
rect 2145 2271 2203 2305
rect 2237 2271 2295 2305
rect 2329 2271 2387 2305
rect 2421 2271 2479 2305
rect 2513 2271 2571 2305
rect 2660 2271 2663 2305
rect 2697 2271 2755 2305
rect 2789 2271 2847 2305
rect 2881 2271 2939 2305
rect 2973 2271 3031 2305
rect 3065 2271 3123 2305
rect 3157 2271 3215 2305
rect 3249 2271 3278 2305
rect 1806 2260 2604 2271
rect 2660 2260 3278 2271
rect 1806 2240 3278 2260
rect 3676 2314 5148 2332
rect 3676 2301 4392 2314
rect 4448 2301 5148 2314
rect 3676 2267 3705 2301
rect 3739 2267 3797 2301
rect 3831 2267 3889 2301
rect 3923 2267 3981 2301
rect 4015 2267 4073 2301
rect 4107 2267 4165 2301
rect 4199 2267 4257 2301
rect 4291 2267 4349 2301
rect 4383 2267 4392 2301
rect 4475 2267 4533 2301
rect 4567 2267 4625 2301
rect 4659 2267 4717 2301
rect 4751 2267 4809 2301
rect 4843 2267 4901 2301
rect 4935 2267 4993 2301
rect 5027 2267 5085 2301
rect 5119 2267 5148 2301
rect 3676 2256 4392 2267
rect 4448 2256 5148 2267
rect 2002 2067 2060 2073
rect 2002 2033 2014 2067
rect 2048 2064 2060 2067
rect 2088 2064 2116 2240
rect 3676 2236 5148 2256
rect 5492 2310 6964 2328
rect 5492 2297 6220 2310
rect 6276 2297 6964 2310
rect 5492 2263 5521 2297
rect 5555 2263 5613 2297
rect 5647 2263 5705 2297
rect 5739 2263 5797 2297
rect 5831 2263 5889 2297
rect 5923 2263 5981 2297
rect 6015 2263 6073 2297
rect 6107 2263 6165 2297
rect 6199 2263 6220 2297
rect 6291 2263 6349 2297
rect 6383 2263 6441 2297
rect 6475 2263 6533 2297
rect 6567 2263 6625 2297
rect 6659 2263 6717 2297
rect 6751 2263 6809 2297
rect 6843 2263 6901 2297
rect 6935 2263 6964 2297
rect 5492 2252 6220 2263
rect 6276 2252 6964 2263
rect 2186 2135 2244 2141
rect 2186 2101 2198 2135
rect 2232 2132 2244 2135
rect 2926 2135 2984 2141
rect 2926 2132 2938 2135
rect 2232 2104 2938 2132
rect 2232 2101 2244 2104
rect 2186 2095 2244 2101
rect 2926 2101 2938 2104
rect 2972 2101 2984 2135
rect 2926 2095 2984 2101
rect 2370 2067 2428 2073
rect 2370 2064 2382 2067
rect 2048 2036 2382 2064
rect 2048 2033 2060 2036
rect 2002 2027 2060 2033
rect 2370 2033 2382 2036
rect 2416 2064 2428 2067
rect 2742 2067 2800 2073
rect 2742 2064 2754 2067
rect 2416 2036 2754 2064
rect 2416 2033 2428 2036
rect 2370 2027 2428 2033
rect 2742 2033 2754 2036
rect 2788 2064 2800 2067
rect 3018 2067 3076 2073
rect 3018 2064 3030 2067
rect 2788 2036 3030 2064
rect 2788 2033 2800 2036
rect 2742 2027 2800 2033
rect 3018 2033 3030 2036
rect 3064 2033 3076 2067
rect 3018 2027 3076 2033
rect 3872 2063 3930 2069
rect 3872 2029 3884 2063
rect 3918 2060 3930 2063
rect 3958 2060 3986 2236
rect 5492 2232 6964 2252
rect 7362 2308 8834 2324
rect 7362 2293 8060 2308
rect 8116 2293 8834 2308
rect 7362 2259 7391 2293
rect 7425 2259 7483 2293
rect 7517 2259 7575 2293
rect 7609 2259 7667 2293
rect 7701 2259 7759 2293
rect 7793 2259 7851 2293
rect 7885 2259 7943 2293
rect 7977 2259 8035 2293
rect 8116 2259 8127 2293
rect 8161 2259 8219 2293
rect 8253 2259 8311 2293
rect 8345 2259 8403 2293
rect 8437 2259 8495 2293
rect 8529 2259 8587 2293
rect 8621 2259 8679 2293
rect 8713 2259 8771 2293
rect 8805 2259 8834 2293
rect 7362 2250 8060 2259
rect 8116 2250 8834 2259
rect 4056 2131 4114 2137
rect 4056 2097 4068 2131
rect 4102 2128 4114 2131
rect 4796 2131 4854 2137
rect 4796 2128 4808 2131
rect 4102 2100 4808 2128
rect 4102 2097 4114 2100
rect 4056 2091 4114 2097
rect 4796 2097 4808 2100
rect 4842 2097 4854 2131
rect 4796 2091 4854 2097
rect 4240 2063 4298 2069
rect 4240 2060 4252 2063
rect 3918 2032 4252 2060
rect 3918 2029 3930 2032
rect 3872 2023 3930 2029
rect 4240 2029 4252 2032
rect 4286 2060 4298 2063
rect 4612 2063 4670 2069
rect 4612 2060 4624 2063
rect 4286 2032 4624 2060
rect 4286 2029 4298 2032
rect 4240 2023 4298 2029
rect 4612 2029 4624 2032
rect 4658 2060 4670 2063
rect 4888 2063 4946 2069
rect 4888 2060 4900 2063
rect 4658 2032 4900 2060
rect 4658 2029 4670 2032
rect 4612 2023 4670 2029
rect 4888 2029 4900 2032
rect 4934 2029 4946 2063
rect 4888 2023 4946 2029
rect 5688 2059 5746 2065
rect 5688 2025 5700 2059
rect 5734 2056 5746 2059
rect 5774 2056 5802 2232
rect 7362 2228 8834 2250
rect 9176 2312 10648 2322
rect 9176 2291 9870 2312
rect 9926 2291 10648 2312
rect 9176 2257 9205 2291
rect 9239 2257 9297 2291
rect 9331 2257 9389 2291
rect 9423 2257 9481 2291
rect 9515 2257 9573 2291
rect 9607 2257 9665 2291
rect 9699 2257 9757 2291
rect 9791 2257 9849 2291
rect 9926 2257 9941 2291
rect 9975 2257 10033 2291
rect 10067 2257 10125 2291
rect 10159 2257 10217 2291
rect 10251 2257 10309 2291
rect 10343 2257 10401 2291
rect 10435 2257 10493 2291
rect 10527 2257 10585 2291
rect 10619 2257 10648 2291
rect 9176 2254 9870 2257
rect 9926 2254 10648 2257
rect 5872 2127 5930 2133
rect 5872 2093 5884 2127
rect 5918 2124 5930 2127
rect 6612 2127 6670 2133
rect 6612 2124 6624 2127
rect 5918 2096 6624 2124
rect 5918 2093 5930 2096
rect 5872 2087 5930 2093
rect 6612 2093 6624 2096
rect 6658 2093 6670 2127
rect 6612 2087 6670 2093
rect 6056 2059 6114 2065
rect 6056 2056 6068 2059
rect 5734 2028 6068 2056
rect 5734 2025 5746 2028
rect 5688 2019 5746 2025
rect 6056 2025 6068 2028
rect 6102 2056 6114 2059
rect 6428 2059 6486 2065
rect 6428 2056 6440 2059
rect 6102 2028 6440 2056
rect 6102 2025 6114 2028
rect 6056 2019 6114 2025
rect 6428 2025 6440 2028
rect 6474 2056 6486 2059
rect 6704 2059 6762 2065
rect 6704 2056 6716 2059
rect 6474 2028 6716 2056
rect 6474 2025 6486 2028
rect 6428 2019 6486 2025
rect 6704 2025 6716 2028
rect 6750 2025 6762 2059
rect 6704 2019 6762 2025
rect 7558 2055 7616 2061
rect 7558 2021 7570 2055
rect 7604 2052 7616 2055
rect 7644 2052 7672 2228
rect 9176 2226 10648 2254
rect 11046 2302 12518 2318
rect 11046 2287 11686 2302
rect 11742 2287 12518 2302
rect 11046 2253 11075 2287
rect 11109 2253 11167 2287
rect 11201 2253 11259 2287
rect 11293 2253 11351 2287
rect 11385 2253 11443 2287
rect 11477 2253 11535 2287
rect 11569 2253 11627 2287
rect 11661 2253 11686 2287
rect 11753 2253 11811 2287
rect 11845 2253 11903 2287
rect 11937 2253 11995 2287
rect 12029 2253 12087 2287
rect 12121 2253 12179 2287
rect 12213 2253 12271 2287
rect 12305 2253 12363 2287
rect 12397 2253 12455 2287
rect 12489 2253 12518 2287
rect 11046 2244 11686 2253
rect 11742 2244 12518 2253
rect 7742 2123 7800 2129
rect 7742 2089 7754 2123
rect 7788 2120 7800 2123
rect 8482 2123 8540 2129
rect 8482 2120 8494 2123
rect 7788 2092 8494 2120
rect 7788 2089 7800 2092
rect 7742 2083 7800 2089
rect 8482 2089 8494 2092
rect 8528 2089 8540 2123
rect 8482 2083 8540 2089
rect 7926 2055 7984 2061
rect 7926 2052 7938 2055
rect 7604 2024 7938 2052
rect 7604 2021 7616 2024
rect 7558 2015 7616 2021
rect 7926 2021 7938 2024
rect 7972 2052 7984 2055
rect 8298 2055 8356 2061
rect 8298 2052 8310 2055
rect 7972 2024 8310 2052
rect 7972 2021 7984 2024
rect 7926 2015 7984 2021
rect 8298 2021 8310 2024
rect 8344 2052 8356 2055
rect 8574 2055 8632 2061
rect 8574 2052 8586 2055
rect 8344 2024 8586 2052
rect 8344 2021 8356 2024
rect 8298 2015 8356 2021
rect 8574 2021 8586 2024
rect 8620 2021 8632 2055
rect 8574 2015 8632 2021
rect 9372 2053 9430 2059
rect 9372 2019 9384 2053
rect 9418 2050 9430 2053
rect 9458 2050 9486 2226
rect 11046 2222 12518 2244
rect 12862 2300 14334 2314
rect 12862 2283 13594 2300
rect 13650 2283 14334 2300
rect 12862 2249 12891 2283
rect 12925 2249 12983 2283
rect 13017 2249 13075 2283
rect 13109 2249 13167 2283
rect 13201 2249 13259 2283
rect 13293 2249 13351 2283
rect 13385 2249 13443 2283
rect 13477 2249 13535 2283
rect 13569 2249 13594 2283
rect 13661 2249 13719 2283
rect 13753 2249 13811 2283
rect 13845 2249 13903 2283
rect 13937 2249 13995 2283
rect 14029 2249 14087 2283
rect 14121 2249 14179 2283
rect 14213 2249 14271 2283
rect 14305 2249 14334 2283
rect 12862 2242 13594 2249
rect 13650 2242 14334 2249
rect 9556 2121 9614 2127
rect 9556 2087 9568 2121
rect 9602 2118 9614 2121
rect 10296 2121 10354 2127
rect 10296 2118 10308 2121
rect 9602 2090 10308 2118
rect 9602 2087 9614 2090
rect 9556 2081 9614 2087
rect 10296 2087 10308 2090
rect 10342 2087 10354 2121
rect 10296 2081 10354 2087
rect 9740 2053 9798 2059
rect 9740 2050 9752 2053
rect 9418 2022 9752 2050
rect 9418 2019 9430 2022
rect 9372 2013 9430 2019
rect 9740 2019 9752 2022
rect 9786 2050 9798 2053
rect 10112 2053 10170 2059
rect 10112 2050 10124 2053
rect 9786 2022 10124 2050
rect 9786 2019 9798 2022
rect 9740 2013 9798 2019
rect 10112 2019 10124 2022
rect 10158 2050 10170 2053
rect 10388 2053 10446 2059
rect 10388 2050 10400 2053
rect 10158 2022 10400 2050
rect 10158 2019 10170 2022
rect 10112 2013 10170 2019
rect 10388 2019 10400 2022
rect 10434 2019 10446 2053
rect 10388 2013 10446 2019
rect 11242 2049 11300 2055
rect 11242 2015 11254 2049
rect 11288 2046 11300 2049
rect 11328 2046 11356 2222
rect 12862 2218 14334 2242
rect 14732 2296 16204 2310
rect 14732 2279 15534 2296
rect 15592 2279 16204 2296
rect 14732 2245 14761 2279
rect 14795 2245 14853 2279
rect 14887 2245 14945 2279
rect 14979 2245 15037 2279
rect 15071 2245 15129 2279
rect 15163 2245 15221 2279
rect 15255 2245 15313 2279
rect 15347 2245 15405 2279
rect 15439 2245 15497 2279
rect 15531 2245 15534 2279
rect 15623 2245 15681 2279
rect 15715 2245 15773 2279
rect 15807 2245 15865 2279
rect 15899 2245 15957 2279
rect 15991 2245 16049 2279
rect 16083 2245 16141 2279
rect 16175 2245 16204 2279
rect 14732 2238 15534 2245
rect 15592 2238 16204 2245
rect 11426 2117 11484 2123
rect 11426 2083 11438 2117
rect 11472 2114 11484 2117
rect 12166 2117 12224 2123
rect 12166 2114 12178 2117
rect 11472 2086 12178 2114
rect 11472 2083 11484 2086
rect 11426 2077 11484 2083
rect 12166 2083 12178 2086
rect 12212 2083 12224 2117
rect 12166 2077 12224 2083
rect 11610 2049 11668 2055
rect 11610 2046 11622 2049
rect 11288 2018 11622 2046
rect 11288 2015 11300 2018
rect 11242 2009 11300 2015
rect 11610 2015 11622 2018
rect 11656 2046 11668 2049
rect 11982 2049 12040 2055
rect 11982 2046 11994 2049
rect 11656 2018 11994 2046
rect 11656 2015 11668 2018
rect 11610 2009 11668 2015
rect 11982 2015 11994 2018
rect 12028 2046 12040 2049
rect 12258 2049 12316 2055
rect 12258 2046 12270 2049
rect 12028 2018 12270 2046
rect 12028 2015 12040 2018
rect 11982 2009 12040 2015
rect 12258 2015 12270 2018
rect 12304 2015 12316 2049
rect 12258 2009 12316 2015
rect 13058 2045 13116 2051
rect 13058 2011 13070 2045
rect 13104 2042 13116 2045
rect 13144 2042 13172 2218
rect 14732 2214 16204 2238
rect 13242 2113 13300 2119
rect 13242 2079 13254 2113
rect 13288 2110 13300 2113
rect 13982 2113 14040 2119
rect 13982 2110 13994 2113
rect 13288 2082 13994 2110
rect 13288 2079 13300 2082
rect 13242 2073 13300 2079
rect 13982 2079 13994 2082
rect 14028 2079 14040 2113
rect 13982 2073 14040 2079
rect 13426 2045 13484 2051
rect 13426 2042 13438 2045
rect 13104 2014 13438 2042
rect 13104 2011 13116 2014
rect 13058 2005 13116 2011
rect 13426 2011 13438 2014
rect 13472 2042 13484 2045
rect 13798 2045 13856 2051
rect 13798 2042 13810 2045
rect 13472 2014 13810 2042
rect 13472 2011 13484 2014
rect 13426 2005 13484 2011
rect 13798 2011 13810 2014
rect 13844 2042 13856 2045
rect 14074 2045 14132 2051
rect 14074 2042 14086 2045
rect 13844 2014 14086 2042
rect 13844 2011 13856 2014
rect 13798 2005 13856 2011
rect 14074 2011 14086 2014
rect 14120 2011 14132 2045
rect 14074 2005 14132 2011
rect 14928 2041 14986 2047
rect 14928 2007 14940 2041
rect 14974 2038 14986 2041
rect 15014 2038 15042 2214
rect 15112 2109 15170 2115
rect 15112 2075 15124 2109
rect 15158 2106 15170 2109
rect 15852 2109 15910 2115
rect 15852 2106 15864 2109
rect 15158 2078 15864 2106
rect 15158 2075 15170 2078
rect 15112 2069 15170 2075
rect 15852 2075 15864 2078
rect 15898 2075 15910 2109
rect 15852 2069 15910 2075
rect 15296 2041 15354 2047
rect 15296 2038 15308 2041
rect 14974 2010 15308 2038
rect 14974 2007 14986 2010
rect 2094 1999 2152 2005
rect 2094 1965 2106 1999
rect 2140 1996 2152 1999
rect 2554 1999 2612 2005
rect 2554 1996 2566 1999
rect 2140 1968 2566 1996
rect 2140 1965 2152 1968
rect 2094 1959 2152 1965
rect 2554 1965 2566 1968
rect 2600 1996 2612 1999
rect 2926 1999 2984 2005
rect 14928 2001 14986 2007
rect 15296 2007 15308 2010
rect 15342 2038 15354 2041
rect 15668 2041 15726 2047
rect 15668 2038 15680 2041
rect 15342 2010 15680 2038
rect 15342 2007 15354 2010
rect 15296 2001 15354 2007
rect 15668 2007 15680 2010
rect 15714 2038 15726 2041
rect 15944 2041 16002 2047
rect 15944 2038 15956 2041
rect 15714 2010 15956 2038
rect 15714 2007 15726 2010
rect 15668 2001 15726 2007
rect 15944 2007 15956 2010
rect 15990 2007 16002 2041
rect 15944 2001 16002 2007
rect 2926 1996 2938 1999
rect 2600 1968 2938 1996
rect 2600 1965 2612 1968
rect 2554 1959 2612 1965
rect 2192 1938 2258 1940
rect 2192 1886 2198 1938
rect 2250 1886 2258 1938
rect 2192 1882 2258 1886
rect 2648 1792 2676 1968
rect 2926 1965 2938 1968
rect 2972 1965 2984 1999
rect 2926 1959 2984 1965
rect 3964 1995 4022 2001
rect 3964 1961 3976 1995
rect 4010 1992 4022 1995
rect 4424 1995 4482 2001
rect 4424 1992 4436 1995
rect 4010 1964 4436 1992
rect 4010 1961 4022 1964
rect 3964 1955 4022 1961
rect 4424 1961 4436 1964
rect 4470 1992 4482 1995
rect 4796 1995 4854 2001
rect 4796 1992 4808 1995
rect 4470 1964 4808 1992
rect 4470 1961 4482 1964
rect 4424 1955 4482 1961
rect 3200 1926 3260 1950
rect 3200 1890 3214 1926
rect 3254 1924 3260 1926
rect 4060 1928 4120 1934
rect 4060 1924 4074 1928
rect 3254 1894 4074 1924
rect 4108 1894 4120 1928
rect 3254 1890 4120 1894
rect 3200 1886 4120 1890
rect 3200 1874 3260 1886
rect 4060 1872 4120 1886
rect 1806 1778 3278 1792
rect 4518 1788 4546 1964
rect 4796 1961 4808 1964
rect 4842 1961 4854 1995
rect 4796 1955 4854 1961
rect 5780 1991 5838 1997
rect 5780 1957 5792 1991
rect 5826 1988 5838 1991
rect 6240 1991 6298 1997
rect 6240 1988 6252 1991
rect 5826 1960 6252 1988
rect 5826 1957 5838 1960
rect 5780 1951 5838 1957
rect 6240 1957 6252 1960
rect 6286 1988 6298 1991
rect 6612 1991 6670 1997
rect 6612 1988 6624 1991
rect 6286 1960 6624 1988
rect 6286 1957 6298 1960
rect 6240 1951 6298 1957
rect 5078 1922 5130 1940
rect 5876 1924 5936 1932
rect 5876 1922 5890 1924
rect 5078 1886 5090 1922
rect 5124 1890 5890 1922
rect 5924 1890 5936 1924
rect 5124 1886 5936 1890
rect 5078 1884 5936 1886
rect 5078 1874 5130 1884
rect 1806 1761 2604 1778
rect 2656 1761 3278 1778
rect 1806 1727 1835 1761
rect 1869 1727 1927 1761
rect 1961 1727 2019 1761
rect 2053 1727 2111 1761
rect 2145 1727 2203 1761
rect 2237 1727 2295 1761
rect 2329 1727 2387 1761
rect 2421 1727 2479 1761
rect 2513 1727 2571 1761
rect 2656 1727 2663 1761
rect 2697 1727 2755 1761
rect 2789 1727 2847 1761
rect 2881 1727 2939 1761
rect 2973 1727 3031 1761
rect 3065 1727 3123 1761
rect 3157 1727 3215 1761
rect 3249 1727 3278 1761
rect 1806 1720 2604 1727
rect 2656 1720 3278 1727
rect 1806 1696 3278 1720
rect 3676 1768 5148 1788
rect 6334 1784 6362 1960
rect 6612 1957 6624 1960
rect 6658 1957 6670 1991
rect 6612 1951 6670 1957
rect 7650 1987 7708 1993
rect 7650 1953 7662 1987
rect 7696 1984 7708 1987
rect 8110 1987 8168 1993
rect 8110 1984 8122 1987
rect 7696 1956 8122 1984
rect 7696 1953 7708 1956
rect 7650 1947 7708 1953
rect 8110 1953 8122 1956
rect 8156 1984 8168 1987
rect 8482 1987 8540 1993
rect 8482 1984 8494 1987
rect 8156 1956 8494 1984
rect 8156 1953 8168 1956
rect 8110 1947 8168 1953
rect 6886 1918 6946 1942
rect 6886 1882 6900 1918
rect 6940 1916 6946 1918
rect 7746 1920 7806 1926
rect 7746 1916 7760 1920
rect 6940 1886 7760 1916
rect 7794 1886 7806 1920
rect 6940 1882 7806 1886
rect 6886 1878 7806 1882
rect 6886 1866 6946 1878
rect 7746 1864 7806 1878
rect 3676 1757 4396 1768
rect 4452 1757 5148 1768
rect 3676 1723 3705 1757
rect 3739 1723 3797 1757
rect 3831 1723 3889 1757
rect 3923 1723 3981 1757
rect 4015 1723 4073 1757
rect 4107 1723 4165 1757
rect 4199 1723 4257 1757
rect 4291 1723 4349 1757
rect 4383 1723 4396 1757
rect 4475 1723 4533 1757
rect 4567 1723 4625 1757
rect 4659 1723 4717 1757
rect 4751 1723 4809 1757
rect 4843 1723 4901 1757
rect 4935 1723 4993 1757
rect 5027 1723 5085 1757
rect 5119 1723 5148 1757
rect 3676 1710 4396 1723
rect 4452 1710 5148 1723
rect 3676 1692 5148 1710
rect 5492 1760 6964 1784
rect 8204 1780 8232 1956
rect 8482 1953 8494 1956
rect 8528 1953 8540 1987
rect 8482 1947 8540 1953
rect 9464 1985 9522 1991
rect 9464 1951 9476 1985
rect 9510 1982 9522 1985
rect 9924 1985 9982 1991
rect 9924 1982 9936 1985
rect 9510 1954 9936 1982
rect 9510 1951 9522 1954
rect 9464 1945 9522 1951
rect 9924 1951 9936 1954
rect 9970 1982 9982 1985
rect 10296 1985 10354 1991
rect 10296 1982 10308 1985
rect 9970 1954 10308 1982
rect 9970 1951 9982 1954
rect 9924 1945 9982 1951
rect 8754 1920 8816 1928
rect 8754 1884 8770 1920
rect 8804 1916 8816 1920
rect 9562 1918 9628 1926
rect 9562 1916 9574 1918
rect 8804 1884 9574 1916
rect 9610 1884 9628 1918
rect 8754 1874 8816 1884
rect 9562 1876 9628 1884
rect 5492 1753 6238 1760
rect 6294 1753 6964 1760
rect 5492 1719 5521 1753
rect 5555 1719 5613 1753
rect 5647 1719 5705 1753
rect 5739 1719 5797 1753
rect 5831 1719 5889 1753
rect 5923 1719 5981 1753
rect 6015 1719 6073 1753
rect 6107 1719 6165 1753
rect 6199 1719 6238 1753
rect 6294 1719 6349 1753
rect 6383 1719 6441 1753
rect 6475 1719 6533 1753
rect 6567 1719 6625 1753
rect 6659 1719 6717 1753
rect 6751 1719 6809 1753
rect 6843 1719 6901 1753
rect 6935 1719 6964 1753
rect 5492 1702 6238 1719
rect 6294 1702 6964 1719
rect 5492 1688 6964 1702
rect 7362 1762 8834 1780
rect 10018 1778 10046 1954
rect 10296 1951 10308 1954
rect 10342 1951 10354 1985
rect 10296 1945 10354 1951
rect 11334 1981 11392 1987
rect 11334 1947 11346 1981
rect 11380 1978 11392 1981
rect 11794 1981 11852 1987
rect 11794 1978 11806 1981
rect 11380 1950 11806 1978
rect 11380 1947 11392 1950
rect 11334 1941 11392 1947
rect 11794 1947 11806 1950
rect 11840 1978 11852 1981
rect 12166 1981 12224 1987
rect 12166 1978 12178 1981
rect 11840 1950 12178 1978
rect 11840 1947 11852 1950
rect 11794 1941 11852 1947
rect 10570 1912 10630 1936
rect 10570 1876 10584 1912
rect 10624 1910 10630 1912
rect 11430 1914 11490 1920
rect 11430 1910 11444 1914
rect 10624 1880 11444 1910
rect 11478 1880 11490 1914
rect 10624 1876 11490 1880
rect 10570 1872 11490 1876
rect 10570 1860 10630 1872
rect 11430 1858 11490 1872
rect 7362 1749 8056 1762
rect 8112 1749 8834 1762
rect 7362 1715 7391 1749
rect 7425 1715 7483 1749
rect 7517 1715 7575 1749
rect 7609 1715 7667 1749
rect 7701 1715 7759 1749
rect 7793 1715 7851 1749
rect 7885 1715 7943 1749
rect 7977 1715 8035 1749
rect 8112 1715 8127 1749
rect 8161 1715 8219 1749
rect 8253 1715 8311 1749
rect 8345 1715 8403 1749
rect 8437 1715 8495 1749
rect 8529 1715 8587 1749
rect 8621 1715 8679 1749
rect 8713 1715 8771 1749
rect 8805 1715 8834 1749
rect 7362 1704 8056 1715
rect 8112 1704 8834 1715
rect 7362 1684 8834 1704
rect 9176 1762 10648 1778
rect 11888 1774 11916 1950
rect 12166 1947 12178 1950
rect 12212 1947 12224 1981
rect 12166 1941 12224 1947
rect 13150 1977 13208 1983
rect 13150 1943 13162 1977
rect 13196 1974 13208 1977
rect 13610 1977 13668 1983
rect 13610 1974 13622 1977
rect 13196 1946 13622 1974
rect 13196 1943 13208 1946
rect 13150 1937 13208 1943
rect 13610 1943 13622 1946
rect 13656 1974 13668 1977
rect 13982 1977 14040 1983
rect 13982 1974 13994 1977
rect 13656 1946 13994 1974
rect 13656 1943 13668 1946
rect 13610 1937 13668 1943
rect 12444 1912 12500 1930
rect 12444 1878 12454 1912
rect 12488 1908 12500 1912
rect 13246 1910 13306 1918
rect 13246 1908 13260 1910
rect 12488 1878 13260 1908
rect 12444 1876 13260 1878
rect 13294 1876 13306 1910
rect 12444 1870 13306 1876
rect 12444 1864 12500 1870
rect 9176 1747 9908 1762
rect 9964 1747 10648 1762
rect 9176 1713 9205 1747
rect 9239 1713 9297 1747
rect 9331 1713 9389 1747
rect 9423 1713 9481 1747
rect 9515 1713 9573 1747
rect 9607 1713 9665 1747
rect 9699 1713 9757 1747
rect 9791 1713 9849 1747
rect 9883 1713 9908 1747
rect 9975 1713 10033 1747
rect 10067 1713 10125 1747
rect 10159 1713 10217 1747
rect 10251 1713 10309 1747
rect 10343 1713 10401 1747
rect 10435 1713 10493 1747
rect 10527 1713 10585 1747
rect 10619 1713 10648 1747
rect 9176 1704 9908 1713
rect 9964 1704 10648 1713
rect 9176 1682 10648 1704
rect 11046 1758 12518 1774
rect 13704 1770 13732 1946
rect 13982 1943 13994 1946
rect 14028 1943 14040 1977
rect 13982 1937 14040 1943
rect 15020 1973 15078 1979
rect 15020 1939 15032 1973
rect 15066 1970 15078 1973
rect 15480 1973 15538 1979
rect 15480 1970 15492 1973
rect 15066 1942 15492 1970
rect 15066 1939 15078 1942
rect 15020 1933 15078 1939
rect 15480 1939 15492 1942
rect 15526 1970 15538 1973
rect 15852 1973 15910 1979
rect 15852 1970 15864 1973
rect 15526 1942 15864 1970
rect 15526 1939 15538 1942
rect 15480 1933 15538 1939
rect 14256 1904 14316 1928
rect 14256 1868 14270 1904
rect 14310 1902 14316 1904
rect 15116 1906 15176 1912
rect 15116 1902 15130 1906
rect 14310 1872 15130 1902
rect 15164 1872 15176 1906
rect 14310 1868 15176 1872
rect 14256 1864 15176 1868
rect 14256 1852 14316 1864
rect 15116 1850 15176 1864
rect 11046 1743 11676 1758
rect 11732 1743 12518 1758
rect 11046 1709 11075 1743
rect 11109 1709 11167 1743
rect 11201 1709 11259 1743
rect 11293 1709 11351 1743
rect 11385 1709 11443 1743
rect 11477 1709 11535 1743
rect 11569 1709 11627 1743
rect 11661 1709 11676 1743
rect 11753 1709 11811 1743
rect 11845 1709 11903 1743
rect 11937 1709 11995 1743
rect 12029 1709 12087 1743
rect 12121 1709 12179 1743
rect 12213 1709 12271 1743
rect 12305 1709 12363 1743
rect 12397 1709 12455 1743
rect 12489 1709 12518 1743
rect 11046 1700 11676 1709
rect 11732 1700 12518 1709
rect 11046 1678 12518 1700
rect 12862 1756 14334 1770
rect 15574 1766 15602 1942
rect 15852 1939 15864 1942
rect 15898 1939 15910 1973
rect 15852 1933 15910 1939
rect 16136 1926 16410 1930
rect 16136 1918 16316 1926
rect 16136 1884 16150 1918
rect 16186 1884 16316 1918
rect 16136 1874 16316 1884
rect 16368 1874 16410 1926
rect 16136 1868 16410 1874
rect 12862 1739 13570 1756
rect 12862 1705 12891 1739
rect 12925 1705 12983 1739
rect 13017 1705 13075 1739
rect 13109 1705 13167 1739
rect 13201 1705 13259 1739
rect 13293 1705 13351 1739
rect 13385 1705 13443 1739
rect 13477 1705 13535 1739
rect 13569 1705 13570 1739
rect 12862 1698 13570 1705
rect 13626 1739 14334 1756
rect 13626 1705 13627 1739
rect 13661 1705 13719 1739
rect 13753 1705 13811 1739
rect 13845 1705 13903 1739
rect 13937 1705 13995 1739
rect 14029 1705 14087 1739
rect 14121 1705 14179 1739
rect 14213 1705 14271 1739
rect 14305 1705 14334 1739
rect 13626 1698 14334 1705
rect 12862 1674 14334 1698
rect 14732 1752 16204 1766
rect 14732 1735 15516 1752
rect 15574 1735 16204 1752
rect 14732 1701 14761 1735
rect 14795 1701 14853 1735
rect 14887 1701 14945 1735
rect 14979 1701 15037 1735
rect 15071 1701 15129 1735
rect 15163 1701 15221 1735
rect 15255 1701 15313 1735
rect 15347 1701 15405 1735
rect 15439 1701 15497 1735
rect 15574 1701 15589 1735
rect 15623 1701 15681 1735
rect 15715 1701 15773 1735
rect 15807 1701 15865 1735
rect 15899 1701 15957 1735
rect 15991 1701 16049 1735
rect 16083 1701 16141 1735
rect 16175 1701 16204 1735
rect 14732 1694 15516 1701
rect 15574 1694 16204 1701
rect 14732 1670 16204 1694
rect 30368 862 30432 5710
rect 30230 820 30578 862
rect 30230 716 30332 820
rect 30436 716 30578 820
rect 30230 638 30578 716
<< via1 >>
rect 9540 17762 9600 17822
rect 6646 17504 6722 17576
rect 9536 17218 9594 17278
rect 11414 16986 11474 17042
rect 4590 16570 4642 16624
rect 4976 16020 5034 16074
rect 4746 15814 4808 15874
rect 6712 15706 6780 15768
rect 6608 15356 6660 15408
rect 4898 15270 4966 15332
rect 6130 15202 6198 15264
rect 7114 15156 7182 15218
rect 4582 14986 4648 15052
rect 5794 14654 5862 14716
rect 5012 14442 5078 14508
rect 4682 14244 4754 14314
rect 6350 14232 6418 14294
rect 7916 14222 7984 14284
rect 9552 16587 9604 16608
rect 9552 16554 9585 16587
rect 9585 16554 9604 16587
rect 10968 16324 11038 16390
rect 9938 16043 9996 16058
rect 9938 16009 9953 16043
rect 9953 16009 9996 16043
rect 9938 16004 9996 16009
rect 9708 15843 9770 15858
rect 9708 15809 9741 15843
rect 9741 15809 9770 15843
rect 9708 15798 9770 15809
rect 11674 15733 11742 15752
rect 11674 15699 11691 15733
rect 11691 15699 11725 15733
rect 11725 15699 11742 15733
rect 11674 15690 11742 15699
rect 9938 15474 9992 15486
rect 9938 15440 9968 15474
rect 9968 15440 9992 15474
rect 9938 15432 9992 15440
rect 9860 15299 9928 15316
rect 9860 15265 9867 15299
rect 9867 15265 9925 15299
rect 9925 15265 9928 15299
rect 9860 15254 9928 15265
rect 9544 15023 9610 15036
rect 9544 14989 9561 15023
rect 9561 14989 9595 15023
rect 9595 14989 9610 15023
rect 9544 14970 9610 14989
rect 11570 15384 11622 15392
rect 11570 15348 11594 15384
rect 11594 15348 11622 15384
rect 11570 15340 11622 15348
rect 11092 15233 11160 15248
rect 11092 15199 11109 15233
rect 11109 15199 11143 15233
rect 11143 15199 11160 15233
rect 11092 15186 11160 15199
rect 12076 15189 12144 15202
rect 12076 15155 12093 15189
rect 12093 15155 12144 15189
rect 12076 15140 12144 15155
rect 9974 14479 10040 14492
rect 9974 14445 10021 14479
rect 10021 14445 10040 14479
rect 9974 14426 10040 14445
rect 9644 14279 9716 14298
rect 9644 14245 9659 14279
rect 9659 14245 9693 14279
rect 9693 14245 9716 14279
rect 9644 14228 9716 14245
rect 6828 13856 6896 13918
rect 7652 13914 7674 13936
rect 7674 13914 7704 13936
rect 7652 13882 7704 13914
rect 4884 13700 4956 13770
rect 9992 13822 10052 13884
rect 5862 13692 5930 13754
rect 7656 13676 7724 13738
rect 9846 13735 9918 13754
rect 9846 13701 9877 13735
rect 9877 13701 9918 13735
rect 9846 13684 9918 13701
rect 5984 13390 6052 13450
rect 4576 13318 4648 13384
rect 7136 13316 7204 13378
rect 9538 13355 9610 13368
rect 9538 13321 9553 13355
rect 9553 13321 9587 13355
rect 9587 13321 9610 13355
rect 9538 13302 9610 13321
rect 10756 14689 10824 14700
rect 10756 14655 10775 14689
rect 10775 14655 10824 14689
rect 10756 14638 10824 14655
rect 11312 14267 11380 14278
rect 11312 14233 11367 14267
rect 11367 14233 11380 14267
rect 11312 14216 11380 14233
rect 16430 16660 16498 16722
rect 17188 16652 17256 16714
rect 18078 16654 18146 16716
rect 18686 16650 18754 16712
rect 19444 16642 19512 16704
rect 20334 16644 20402 16706
rect 21450 16644 21518 16706
rect 22208 16636 22276 16698
rect 23098 16638 23166 16700
rect 16410 16122 16478 16184
rect 17196 16112 17264 16174
rect 18076 16112 18144 16174
rect 18666 16112 18734 16174
rect 19452 16102 19520 16164
rect 20332 16102 20400 16164
rect 21430 16106 21498 16168
rect 22216 16096 22284 16158
rect 23096 16096 23164 16158
rect 24400 14810 24462 14870
rect 24144 14662 24196 14714
rect 12878 14251 12946 14268
rect 12878 14217 12909 14251
rect 12909 14217 12943 14251
rect 12943 14217 12946 14251
rect 12878 14206 12946 14217
rect 24452 14552 24504 14564
rect 24452 14518 24456 14552
rect 24456 14518 24492 14552
rect 24492 14518 24504 14552
rect 24452 14512 24504 14518
rect 24552 14554 24556 14578
rect 24556 14554 24592 14578
rect 24592 14554 24604 14578
rect 24552 14526 24604 14554
rect 24698 14528 24712 14536
rect 24712 14528 24746 14536
rect 24746 14528 24750 14536
rect 24698 14484 24750 14528
rect 23992 14258 24054 14318
rect 10260 13288 10322 13340
rect 10974 13864 11026 13874
rect 10974 13830 10982 13864
rect 10982 13830 11016 13864
rect 11016 13830 11026 13864
rect 10974 13822 11026 13830
rect 11072 13904 11124 13914
rect 11072 13870 11080 13904
rect 11080 13870 11114 13904
rect 11114 13870 11124 13904
rect 11072 13862 11124 13870
rect 11170 13814 11222 13870
rect 11790 13893 11858 13902
rect 11790 13859 11819 13893
rect 11819 13859 11858 13893
rect 11790 13840 11858 13859
rect 12614 13898 12636 13920
rect 12636 13898 12666 13920
rect 12614 13866 12666 13898
rect 12748 13944 12828 13964
rect 12748 13902 12762 13944
rect 12762 13902 12812 13944
rect 12812 13902 12828 13944
rect 12748 13888 12828 13902
rect 10824 13723 10892 13738
rect 10824 13689 10849 13723
rect 10849 13689 10892 13723
rect 10824 13676 10892 13689
rect 12618 13707 12686 13722
rect 12618 13673 12633 13707
rect 12633 13673 12667 13707
rect 12667 13673 12686 13707
rect 12618 13660 12686 13673
rect 10946 13425 11014 13434
rect 10946 13391 10973 13425
rect 10973 13391 11014 13425
rect 10946 13374 11014 13391
rect 11102 13318 11156 13322
rect 11102 13282 11108 13318
rect 11108 13282 11144 13318
rect 11144 13282 11156 13318
rect 11102 13270 11156 13282
rect 12098 13349 12166 13362
rect 12098 13315 12153 13349
rect 12153 13315 12166 13349
rect 12098 13300 12166 13315
rect 5996 12856 6064 12916
rect 4990 12778 5062 12844
rect 11158 13050 11210 13066
rect 11158 13016 11194 13050
rect 11194 13016 11210 13050
rect 11158 13012 11210 13016
rect 9952 12811 10024 12828
rect 9952 12777 9955 12811
rect 9955 12777 10013 12811
rect 10013 12777 10024 12811
rect 9952 12762 10024 12777
rect 4634 12576 4708 12642
rect 9596 12611 9670 12626
rect 9596 12577 9651 12611
rect 9651 12577 9670 12611
rect 9596 12560 9670 12577
rect 6280 12370 6348 12432
rect 9968 12306 10030 12374
rect 4906 12034 4980 12100
rect 10958 12881 11026 12900
rect 10958 12847 10973 12881
rect 10973 12847 11026 12881
rect 10958 12840 11026 12847
rect 11242 12405 11310 12416
rect 11242 12371 11245 12405
rect 11245 12371 11303 12405
rect 11303 12371 11310 12405
rect 11242 12354 11310 12371
rect 11302 12180 11354 12192
rect 11302 12146 11308 12180
rect 11308 12146 11342 12180
rect 11342 12146 11354 12180
rect 11302 12140 11354 12146
rect 9868 12067 9942 12084
rect 9868 12033 9869 12067
rect 9869 12033 9927 12067
rect 9927 12033 9942 12067
rect 9868 12018 9942 12033
rect 11112 12094 11164 12102
rect 11112 12060 11120 12094
rect 11120 12060 11156 12094
rect 11156 12060 11164 12094
rect 11112 12050 11164 12060
rect 6002 11830 6070 11892
rect 4560 11756 4640 11820
rect 9522 11791 9602 11804
rect 9522 11757 9563 11791
rect 9563 11757 9597 11791
rect 9597 11757 9602 11791
rect 9522 11740 9602 11757
rect 10964 11861 11032 11876
rect 10964 11827 10969 11861
rect 10969 11827 11027 11861
rect 11027 11827 11032 11861
rect 10964 11814 11032 11827
rect 4994 11214 5074 11278
rect 9956 11247 10036 11262
rect 9956 11213 9965 11247
rect 9965 11213 10023 11247
rect 10023 11213 10036 11247
rect 9956 11198 10036 11213
rect 4626 11010 4706 11074
rect 9588 11047 9668 11058
rect 9588 11013 9603 11047
rect 9603 11013 9661 11047
rect 9661 11013 9668 11047
rect 9588 10994 9668 11013
rect 5054 10676 5108 10732
rect 4904 10476 4984 10540
rect 10016 10660 10070 10716
rect 9866 10503 9946 10524
rect 9866 10469 9879 10503
rect 9879 10469 9937 10503
rect 9937 10469 9946 10503
rect 9866 10460 9946 10469
rect 6226 6617 6282 6638
rect 6226 6583 6233 6617
rect 6233 6583 6267 6617
rect 6267 6583 6282 6617
rect 6226 6580 6282 6583
rect 6168 6382 6220 6390
rect 6168 6348 6178 6382
rect 6178 6348 6212 6382
rect 6212 6348 6220 6382
rect 6168 6338 6220 6348
rect 6268 6384 6320 6396
rect 6268 6350 6274 6384
rect 6274 6350 6308 6384
rect 6308 6350 6320 6384
rect 6268 6344 6320 6350
rect 6170 6073 6226 6088
rect 6170 6039 6175 6073
rect 6175 6039 6226 6073
rect 6170 6030 6226 6039
rect 9606 5985 9664 6002
rect 9974 5985 10032 6000
rect 9606 5951 9615 5985
rect 9615 5951 9649 5985
rect 9649 5951 9664 5985
rect 9974 5951 9983 5985
rect 9983 5951 10017 5985
rect 10017 5951 10032 5985
rect 9606 5940 9664 5951
rect 9974 5936 10032 5951
rect 11866 5981 11924 5998
rect 11866 5947 11887 5981
rect 11887 5947 11924 5981
rect 11866 5934 11924 5947
rect 13652 5977 13710 5988
rect 13652 5943 13669 5977
rect 13669 5943 13703 5977
rect 13703 5943 13710 5977
rect 13652 5924 13710 5943
rect 15534 5973 15592 5992
rect 15534 5939 15539 5973
rect 15539 5939 15573 5973
rect 15573 5939 15592 5973
rect 15534 5928 15592 5939
rect 2564 5565 2620 5578
rect 2564 5531 2601 5565
rect 2601 5531 2620 5565
rect 2564 5520 2620 5531
rect 4444 5561 4500 5574
rect 4444 5527 4471 5561
rect 4471 5527 4500 5561
rect 4444 5516 4500 5527
rect 6166 5557 6222 5576
rect 6166 5523 6195 5557
rect 6195 5523 6222 5557
rect 6166 5518 6222 5523
rect 8076 5553 8132 5566
rect 9610 5614 9662 5618
rect 9610 5580 9618 5614
rect 9618 5580 9652 5614
rect 9652 5580 9662 5614
rect 9610 5566 9662 5580
rect 8076 5519 8099 5553
rect 8099 5519 8132 5553
rect 8076 5508 8132 5519
rect 10414 5441 10470 5452
rect 10414 5407 10443 5441
rect 10443 5407 10470 5441
rect 10414 5394 10470 5407
rect 11370 5437 11428 5456
rect 11370 5403 11393 5437
rect 11393 5403 11427 5437
rect 11427 5403 11428 5437
rect 11370 5392 11428 5403
rect 14072 5433 14130 5450
rect 14072 5399 14129 5433
rect 14129 5399 14130 5433
rect 14072 5386 14130 5399
rect 14992 5429 15050 5442
rect 14992 5395 15021 5429
rect 15021 5395 15050 5429
rect 14992 5378 15050 5395
rect 17226 5364 17284 5428
rect 2228 5194 2280 5198
rect 2228 5160 2236 5194
rect 2236 5160 2270 5194
rect 2270 5160 2280 5194
rect 2228 5146 2280 5160
rect 2584 5021 2640 5040
rect 2584 4987 2601 5021
rect 2601 4987 2635 5021
rect 2635 4987 2640 5021
rect 2584 4982 2640 4987
rect 4444 5017 4500 5032
rect 4444 4983 4471 5017
rect 4471 4983 4500 5017
rect 4444 4974 4500 4983
rect 9388 5111 9444 5120
rect 9388 5077 9401 5111
rect 9401 5077 9444 5111
rect 9388 5062 9444 5077
rect 12276 5107 12334 5120
rect 12276 5073 12283 5107
rect 12283 5073 12334 5107
rect 12276 5056 12334 5073
rect 6148 5013 6204 5028
rect 6148 4979 6195 5013
rect 6195 4979 6204 5013
rect 6148 4970 6204 4979
rect 8064 5009 8120 5020
rect 8064 4975 8065 5009
rect 8065 4975 8099 5009
rect 8099 4975 8120 5009
rect 8064 4962 8120 4975
rect 13130 5103 13188 5116
rect 13130 5069 13145 5103
rect 13145 5069 13179 5103
rect 13179 5069 13188 5103
rect 13130 5052 13188 5069
rect 15922 5099 15980 5114
rect 15922 5065 15935 5099
rect 15935 5065 15969 5099
rect 15969 5065 15980 5099
rect 15922 5050 15980 5065
rect 17556 5042 17608 5050
rect 17556 5004 17564 5042
rect 17564 5004 17602 5042
rect 17602 5004 17608 5042
rect 17556 4998 17608 5004
rect 9638 4740 9690 4744
rect 9638 4706 9646 4740
rect 9646 4706 9680 4740
rect 9680 4706 9690 4740
rect 9638 4692 9690 4706
rect 9988 4567 10044 4580
rect 9640 4533 9643 4566
rect 9643 4533 9677 4566
rect 9677 4533 9692 4566
rect 9988 4533 10011 4567
rect 10011 4533 10044 4567
rect 9640 4512 9692 4533
rect 9988 4522 10044 4533
rect 11894 4563 11952 4578
rect 11894 4529 11915 4563
rect 11915 4529 11952 4563
rect 11894 4514 11952 4529
rect 17220 4816 17278 4880
rect 13698 4559 13756 4574
rect 13698 4525 13731 4559
rect 13731 4525 13756 4559
rect 13698 4510 13756 4525
rect 15628 4555 15686 4566
rect 15628 4521 15659 4555
rect 15659 4521 15686 4555
rect 15628 4502 15686 4521
rect 6194 3320 6254 3382
rect 6138 3122 6190 3130
rect 6138 3088 6148 3122
rect 6148 3088 6182 3122
rect 6182 3088 6190 3122
rect 6138 3078 6190 3088
rect 6238 3124 6290 3136
rect 6238 3090 6244 3124
rect 6244 3090 6278 3124
rect 6278 3090 6290 3124
rect 6238 3084 6290 3090
rect 6176 2766 6236 2828
rect 2604 2305 2660 2318
rect 2604 2271 2605 2305
rect 2605 2271 2660 2305
rect 2604 2260 2660 2271
rect 4392 2301 4448 2314
rect 4392 2267 4441 2301
rect 4441 2267 4448 2301
rect 4392 2256 4448 2267
rect 6220 2297 6276 2310
rect 6220 2263 6257 2297
rect 6257 2263 6276 2297
rect 6220 2252 6276 2263
rect 8060 2293 8116 2308
rect 8060 2259 8069 2293
rect 8069 2259 8116 2293
rect 8060 2250 8116 2259
rect 9870 2291 9926 2312
rect 9870 2257 9883 2291
rect 9883 2257 9926 2291
rect 9870 2254 9926 2257
rect 11686 2287 11742 2302
rect 11686 2253 11719 2287
rect 11719 2253 11742 2287
rect 11686 2244 11742 2253
rect 13594 2283 13650 2300
rect 13594 2249 13627 2283
rect 13627 2249 13650 2283
rect 13594 2242 13650 2249
rect 15534 2279 15592 2296
rect 15534 2245 15589 2279
rect 15589 2245 15592 2279
rect 15534 2238 15592 2245
rect 2198 1934 2250 1938
rect 2198 1900 2206 1934
rect 2206 1900 2240 1934
rect 2240 1900 2250 1934
rect 2198 1886 2250 1900
rect 2604 1761 2656 1778
rect 2604 1727 2605 1761
rect 2605 1727 2656 1761
rect 2604 1720 2656 1727
rect 4396 1757 4452 1768
rect 4396 1723 4441 1757
rect 4441 1723 4452 1757
rect 4396 1710 4452 1723
rect 6238 1753 6294 1760
rect 6238 1719 6257 1753
rect 6257 1719 6291 1753
rect 6291 1719 6294 1753
rect 6238 1702 6294 1719
rect 8056 1749 8112 1762
rect 8056 1715 8069 1749
rect 8069 1715 8112 1749
rect 8056 1704 8112 1715
rect 9908 1747 9964 1762
rect 9908 1713 9941 1747
rect 9941 1713 9964 1747
rect 9908 1704 9964 1713
rect 11676 1743 11732 1758
rect 11676 1709 11719 1743
rect 11719 1709 11732 1743
rect 11676 1700 11732 1709
rect 16316 1874 16368 1926
rect 13570 1698 13626 1756
rect 15516 1735 15574 1752
rect 15516 1701 15531 1735
rect 15531 1701 15574 1735
rect 15516 1694 15574 1701
rect 30332 716 30436 820
<< metal2 >>
rect 9430 17822 9706 17844
rect 9430 17762 9540 17822
rect 9600 17762 9706 17822
rect 9430 17746 9706 17762
rect 6463 17587 6545 17588
rect 6463 17586 6759 17587
rect 6463 17576 6760 17586
rect 6463 17505 6646 17576
rect 4472 16624 4732 16636
rect 4472 16614 4590 16624
rect 4472 16558 4552 16614
rect 4642 16570 4732 16624
rect 4608 16558 4732 16570
rect 4472 16536 4732 16558
rect 4886 16076 5106 16090
rect 4886 16020 4976 16076
rect 5034 16020 5106 16076
rect 4886 15994 5106 16020
rect 4562 15874 4938 15880
rect 4562 15814 4746 15874
rect 4808 15814 4938 15874
rect 4562 15792 4938 15814
rect 6463 15424 6545 17505
rect 6604 17504 6646 17505
rect 6722 17504 6760 17576
rect 6604 17498 6760 17504
rect 9432 17278 9706 17302
rect 9432 17218 9536 17278
rect 9594 17218 9706 17278
rect 9432 17202 9706 17218
rect 11401 17054 11483 17055
rect 11400 17042 11506 17054
rect 11400 16986 11414 17042
rect 11474 17033 11506 17042
rect 11474 16986 11507 17033
rect 11400 16762 11507 16986
rect 9434 16608 9694 16620
rect 9434 16598 9552 16608
rect 9434 16542 9514 16598
rect 9604 16554 9694 16608
rect 9570 16542 9694 16554
rect 9434 16520 9694 16542
rect 10908 16390 11110 16422
rect 10908 16324 10968 16390
rect 11038 16324 11110 16390
rect 10908 16296 11110 16324
rect 9848 16060 10068 16074
rect 9848 16004 9938 16060
rect 9996 16004 10068 16060
rect 9848 15978 10068 16004
rect 9524 15858 9900 15864
rect 9524 15798 9708 15858
rect 9770 15798 9900 15858
rect 6608 15768 6894 15780
rect 9524 15776 9900 15798
rect 6608 15706 6712 15768
rect 6780 15706 6894 15768
rect 6608 15684 6894 15706
rect 9920 15486 10028 15494
rect 9920 15432 9938 15486
rect 9992 15456 10028 15486
rect 9992 15432 10420 15456
rect 6463 15408 6682 15424
rect 9920 15420 10420 15432
rect 6463 15356 6608 15408
rect 6660 15356 6682 15408
rect 4836 15332 5028 15350
rect 6463 15342 6682 15356
rect 4836 15270 4898 15332
rect 4966 15270 5028 15332
rect 9798 15316 9990 15334
rect 4836 15254 5028 15270
rect 6108 15264 6254 15280
rect 6108 15202 6130 15264
rect 6198 15202 6254 15264
rect 9798 15254 9860 15316
rect 9928 15254 9990 15316
rect 9798 15238 9990 15254
rect 6108 15184 6254 15202
rect 7046 15218 7252 15238
rect 7046 15156 7114 15218
rect 7182 15156 7252 15218
rect 7046 15140 7252 15156
rect 4476 15052 4750 15070
rect 4476 14986 4582 15052
rect 4648 14986 4750 15052
rect 4476 14978 4750 14986
rect 9438 15036 9712 15054
rect 9438 14970 9544 15036
rect 9610 14970 9712 15036
rect 9438 14962 9712 14970
rect 5748 14716 5908 14736
rect 5748 14654 5794 14716
rect 5862 14654 5908 14716
rect 5748 14640 5908 14654
rect 4946 14508 5118 14524
rect 4946 14442 5012 14508
rect 5078 14442 5118 14508
rect 4946 14434 5118 14442
rect 7635 14487 8531 14581
rect 4576 14314 4870 14320
rect 4576 14244 4682 14314
rect 4754 14244 4870 14314
rect 4576 14232 4870 14244
rect 6322 14294 6470 14316
rect 6322 14232 6350 14294
rect 6418 14232 6470 14294
rect 6322 14218 6470 14232
rect 6794 13918 6946 13938
rect 6794 13856 6828 13918
rect 6896 13856 6946 13918
rect 7635 13936 7729 14487
rect 7840 14284 8072 14296
rect 7840 14222 7916 14284
rect 7984 14222 8072 14284
rect 7840 14204 8072 14222
rect 7635 13882 7652 13936
rect 7704 13882 7729 13936
rect 7635 13857 7729 13882
rect 6794 13842 6946 13856
rect 4820 13770 5040 13780
rect 4820 13700 4884 13770
rect 4956 13700 5040 13770
rect 4820 13684 5040 13700
rect 5824 13754 5974 13770
rect 5824 13692 5862 13754
rect 5930 13692 5974 13754
rect 5824 13672 5974 13692
rect 7642 13738 7744 13754
rect 7642 13676 7656 13738
rect 7724 13676 7744 13738
rect 7642 13658 7744 13676
rect 5950 13450 6084 13470
rect 4468 13384 4738 13396
rect 4468 13318 4576 13384
rect 4648 13318 4738 13384
rect 5950 13390 5984 13450
rect 6052 13390 6084 13450
rect 5950 13378 6084 13390
rect 7096 13378 7248 13396
rect 4468 13310 4738 13318
rect 7096 13316 7136 13378
rect 7204 13316 7248 13378
rect 7096 13300 7248 13316
rect 5948 12916 6100 12928
rect 5948 12856 5996 12916
rect 6064 12856 6100 12916
rect 4922 12844 5112 12854
rect 4922 12778 4990 12844
rect 5062 12778 5112 12844
rect 5948 12834 6100 12856
rect 4922 12766 5112 12778
rect 4574 12642 4780 12654
rect 4574 12576 4634 12642
rect 4708 12576 4780 12642
rect 4574 12560 4780 12576
rect 6230 12432 6402 12452
rect 6230 12370 6280 12432
rect 6348 12370 6402 12432
rect 6230 12356 6402 12370
rect 4858 12100 5024 12116
rect 4858 12034 4906 12100
rect 4980 12034 5024 12100
rect 4858 12022 5024 12034
rect 5944 11892 6100 11908
rect 4510 11820 4690 11834
rect 4510 11756 4560 11820
rect 4640 11756 4690 11820
rect 5944 11830 6002 11892
rect 6070 11830 6100 11892
rect 5944 11812 6100 11830
rect 4510 11746 4690 11756
rect 4938 11278 5118 11292
rect 4938 11214 4994 11278
rect 5074 11214 5118 11278
rect 4938 11204 5118 11214
rect 4580 11074 4776 11092
rect 4580 11010 4626 11074
rect 4706 11010 4776 11074
rect 4580 10996 4776 11010
rect 8437 10762 8531 14487
rect 9908 14492 10080 14508
rect 9908 14426 9974 14492
rect 10040 14426 10080 14492
rect 9908 14418 10080 14426
rect 9538 14298 9832 14304
rect 9538 14228 9644 14298
rect 9716 14228 9832 14298
rect 9538 14216 9832 14228
rect 10384 14082 10420 15420
rect 10710 14700 10870 14720
rect 10710 14638 10756 14700
rect 10824 14638 10870 14700
rect 10710 14624 10870 14638
rect 10972 14494 11040 16296
rect 11425 15408 11507 16762
rect 16346 16722 16558 16738
rect 16346 16660 16430 16722
rect 16498 16660 16558 16722
rect 16346 16646 16558 16660
rect 17116 16714 17328 16732
rect 17116 16652 17188 16714
rect 17256 16652 17328 16714
rect 17116 16640 17328 16652
rect 18008 16716 18220 16732
rect 18008 16654 18078 16716
rect 18146 16654 18220 16716
rect 18008 16640 18220 16654
rect 18602 16712 18814 16728
rect 18602 16650 18686 16712
rect 18754 16650 18814 16712
rect 18602 16636 18814 16650
rect 19372 16704 19584 16722
rect 19372 16642 19444 16704
rect 19512 16642 19584 16704
rect 19372 16630 19584 16642
rect 20264 16706 20476 16722
rect 20264 16644 20334 16706
rect 20402 16644 20476 16706
rect 20264 16630 20476 16644
rect 21366 16706 21578 16722
rect 21366 16644 21450 16706
rect 21518 16644 21578 16706
rect 21366 16630 21578 16644
rect 22136 16698 22348 16716
rect 22136 16636 22208 16698
rect 22276 16636 22348 16698
rect 22136 16624 22348 16636
rect 23028 16700 23240 16716
rect 23028 16638 23098 16700
rect 23166 16638 23240 16700
rect 23028 16624 23240 16638
rect 16336 16184 16548 16194
rect 16336 16122 16410 16184
rect 16478 16122 16548 16184
rect 16336 16102 16548 16122
rect 17126 16174 17338 16186
rect 17126 16112 17196 16174
rect 17264 16112 17338 16174
rect 17126 16094 17338 16112
rect 17996 16174 18208 16186
rect 17996 16112 18076 16174
rect 18144 16112 18208 16174
rect 17996 16094 18208 16112
rect 18592 16174 18804 16184
rect 18592 16112 18666 16174
rect 18734 16112 18804 16174
rect 18592 16092 18804 16112
rect 19382 16164 19594 16176
rect 19382 16102 19452 16164
rect 19520 16102 19594 16164
rect 19382 16084 19594 16102
rect 20252 16164 20464 16176
rect 20252 16102 20332 16164
rect 20400 16102 20464 16164
rect 20252 16084 20464 16102
rect 21356 16168 21568 16178
rect 21356 16106 21430 16168
rect 21498 16106 21568 16168
rect 21356 16086 21568 16106
rect 22146 16158 22358 16170
rect 22146 16096 22216 16158
rect 22284 16096 22358 16158
rect 22146 16078 22358 16096
rect 23016 16158 23228 16170
rect 23016 16096 23096 16158
rect 23164 16096 23228 16158
rect 23016 16078 23228 16096
rect 11570 15752 11856 15764
rect 11570 15690 11674 15752
rect 11742 15690 11856 15752
rect 11570 15668 11856 15690
rect 11425 15392 11644 15408
rect 11425 15340 11570 15392
rect 11622 15340 11644 15392
rect 11425 15326 11644 15340
rect 11070 15248 11216 15264
rect 11070 15186 11092 15248
rect 11160 15186 11216 15248
rect 11070 15168 11216 15186
rect 12008 15202 12214 15222
rect 12008 15140 12076 15202
rect 12144 15140 12214 15202
rect 12008 15124 12214 15140
rect 24312 14870 24542 14880
rect 24312 14810 24400 14870
rect 24462 14810 24542 14870
rect 24312 14788 24542 14810
rect 26389 14843 27464 14921
rect 26389 14740 26467 14843
rect 26948 14766 27172 14794
rect 26389 14726 26466 14740
rect 24138 14714 26466 14726
rect 24138 14662 24144 14714
rect 24196 14662 26466 14714
rect 24138 14658 26466 14662
rect 13142 14565 13434 14581
rect 10972 14426 11130 14494
rect 10384 14046 10994 14082
rect 10958 13920 10994 14046
rect 9930 13884 10100 13896
rect 9930 13822 9992 13884
rect 10052 13864 10100 13884
rect 10958 13874 11034 13920
rect 10958 13864 10974 13874
rect 10052 13822 10676 13864
rect 9930 13816 10676 13822
rect 10956 13822 10974 13864
rect 11026 13822 11034 13874
rect 10956 13816 11034 13822
rect 9930 13802 10100 13816
rect 9782 13754 10002 13764
rect 9782 13684 9846 13754
rect 9918 13684 10002 13754
rect 9782 13668 10002 13684
rect 10626 13576 10674 13816
rect 10964 13778 11034 13816
rect 11062 13914 11130 14426
rect 12597 14471 13493 14565
rect 24138 14488 24198 14658
rect 26389 14657 26466 14658
rect 26948 14646 27000 14766
rect 27122 14726 27172 14766
rect 27122 14658 27176 14726
rect 27122 14646 27172 14658
rect 24448 14564 24504 14620
rect 24448 14512 24452 14564
rect 11284 14278 11432 14300
rect 11284 14216 11312 14278
rect 11380 14216 11432 14278
rect 11284 14202 11432 14216
rect 11062 13862 11072 13914
rect 11124 13862 11130 13914
rect 11062 13776 11130 13862
rect 11163 13870 11237 13969
rect 11163 13814 11170 13870
rect 11222 13814 11237 13870
rect 11756 13902 11908 13922
rect 11756 13840 11790 13902
rect 11858 13840 11908 13902
rect 12597 13920 12691 14471
rect 12802 14268 13034 14280
rect 12802 14206 12878 14268
rect 12946 14206 13034 14268
rect 12802 14188 13034 14206
rect 12597 13866 12614 13920
rect 12666 13866 12691 13920
rect 12720 13964 12858 13976
rect 12720 13888 12748 13964
rect 12828 13888 12858 13964
rect 12720 13874 12858 13888
rect 12597 13841 12691 13866
rect 11756 13826 11908 13840
rect 11163 13785 11237 13814
rect 10786 13738 10936 13754
rect 10786 13676 10824 13738
rect 10892 13676 10936 13738
rect 11163 13711 11305 13785
rect 10786 13656 10936 13676
rect 10626 13528 11136 13576
rect 10912 13434 11046 13454
rect 9430 13368 9700 13380
rect 9430 13302 9538 13368
rect 9610 13302 9700 13368
rect 10912 13374 10946 13434
rect 11014 13374 11046 13434
rect 10912 13362 11046 13374
rect 11088 13356 11136 13528
rect 10322 13350 10728 13352
rect 9430 13294 9700 13302
rect 10252 13340 10728 13350
rect 10252 13288 10260 13340
rect 10322 13288 10728 13340
rect 10252 13280 10728 13288
rect 10656 13154 10728 13280
rect 11082 13322 11180 13356
rect 11082 13270 11102 13322
rect 11156 13270 11180 13322
rect 11082 13252 11180 13270
rect 11231 13156 11305 13711
rect 12604 13722 12706 13738
rect 12604 13660 12618 13722
rect 12686 13660 12706 13722
rect 12604 13642 12706 13660
rect 12058 13362 12210 13380
rect 12058 13300 12098 13362
rect 12166 13300 12210 13362
rect 12058 13284 12210 13300
rect 11102 13154 11305 13156
rect 10656 13082 11305 13154
rect 11148 13066 11220 13082
rect 11148 13012 11158 13066
rect 11210 13012 11220 13066
rect 11148 12928 11220 13012
rect 10910 12900 11062 12912
rect 10910 12840 10958 12900
rect 11026 12840 11062 12900
rect 9884 12828 10074 12838
rect 9884 12762 9952 12828
rect 10024 12762 10074 12828
rect 10910 12818 11062 12840
rect 9884 12750 10074 12762
rect 9536 12626 9742 12638
rect 9536 12560 9596 12626
rect 9670 12560 9742 12626
rect 9536 12544 9742 12560
rect 11192 12416 11364 12436
rect 9922 12374 10072 12388
rect 9922 12306 9968 12374
rect 10030 12322 10072 12374
rect 11192 12354 11242 12416
rect 11310 12354 11364 12416
rect 11192 12340 11364 12354
rect 10030 12306 11152 12322
rect 9922 12290 11152 12306
rect 11120 12110 11152 12290
rect 12740 12202 12808 13874
rect 11296 12192 12808 12202
rect 11296 12140 11302 12192
rect 11354 12140 12808 12192
rect 11296 12134 12808 12140
rect 11104 12102 11174 12110
rect 9820 12084 9986 12100
rect 9820 12018 9868 12084
rect 9942 12018 9986 12084
rect 11104 12050 11112 12102
rect 11164 12050 11174 12102
rect 11104 12044 11174 12050
rect 9820 12006 9986 12018
rect 10906 11876 11062 11892
rect 9472 11804 9652 11818
rect 9472 11740 9522 11804
rect 9602 11740 9652 11804
rect 10906 11814 10964 11876
rect 11032 11814 11062 11876
rect 10906 11796 11062 11814
rect 9472 11730 9652 11740
rect 9900 11262 10080 11276
rect 9900 11198 9956 11262
rect 10036 11198 10080 11262
rect 9900 11188 10080 11198
rect 9542 11058 9738 11076
rect 9542 10994 9588 11058
rect 9668 10994 9738 11058
rect 9542 10980 9738 10994
rect 13341 10762 13493 14471
rect 23850 14318 24212 14334
rect 23850 14258 23992 14318
rect 24054 14258 24212 14318
rect 23850 14240 24212 14258
rect 24448 14112 24504 14512
rect 24546 14578 24606 14622
rect 24546 14526 24552 14578
rect 24604 14526 24606 14578
rect 24448 14056 24502 14112
rect 4970 10732 8531 10762
rect 13142 10746 13493 10762
rect 4970 10676 5054 10732
rect 5108 10676 8531 10732
rect 4970 10668 8531 10676
rect 9932 10716 13493 10746
rect 4970 10652 5202 10668
rect 9932 10660 10016 10716
rect 10070 10660 13493 10716
rect 9932 10652 13493 10660
rect 23258 14000 24502 14056
rect 9932 10636 10164 10652
rect 4856 10540 5036 10546
rect 4856 10476 4904 10540
rect 4984 10476 5036 10540
rect 4856 10458 5036 10476
rect 9818 10524 9998 10530
rect 9818 10460 9866 10524
rect 9946 10460 9998 10524
rect 9818 10442 9998 10460
rect 6112 6638 6388 6648
rect 6112 6580 6226 6638
rect 6282 6580 6388 6638
rect 6112 6558 6388 6580
rect 5585 6398 5651 6404
rect 2222 6390 6228 6398
rect 2222 6338 6168 6390
rect 6220 6338 6228 6390
rect 6262 6396 13156 6398
rect 6262 6344 6268 6396
rect 6320 6394 13156 6396
rect 23258 6394 23314 14000
rect 24546 13290 24606 14526
rect 24684 14536 24776 14624
rect 26948 14604 27172 14646
rect 24684 14484 24698 14536
rect 24750 14514 24776 14536
rect 26993 14514 27071 14604
rect 24750 14484 27071 14514
rect 24684 14436 27071 14484
rect 27386 14514 27464 14843
rect 27386 14510 27604 14514
rect 27386 14492 27730 14510
rect 27386 14436 27550 14492
rect 27512 14372 27550 14436
rect 27682 14372 27730 14492
rect 27512 14336 27730 14372
rect 6320 6344 23314 6394
rect 6262 6338 23314 6344
rect 24252 13230 24608 13290
rect 2222 6332 6228 6338
rect 2222 5198 2290 6332
rect 6110 6088 6274 6104
rect 6110 6030 6170 6088
rect 6226 6030 6274 6088
rect 6110 6018 6274 6030
rect 9604 6002 9672 6018
rect 9604 5940 9606 6002
rect 9664 5940 9672 6002
rect 9604 5618 9672 5940
rect 9908 6000 10088 6016
rect 9908 5936 9974 6000
rect 10032 5936 10088 6000
rect 9908 5922 10088 5936
rect 11800 5998 11982 6006
rect 11800 5934 11866 5998
rect 11924 5934 11982 5998
rect 11800 5910 11982 5934
rect 13570 5988 13752 6010
rect 13570 5924 13652 5988
rect 13710 5924 13752 5988
rect 13570 5914 13752 5924
rect 15464 5992 15644 6004
rect 15464 5928 15534 5992
rect 15592 5928 15644 5992
rect 15464 5912 15644 5928
rect 2510 5578 2690 5596
rect 2510 5520 2564 5578
rect 2620 5520 2690 5578
rect 2510 5502 2690 5520
rect 4378 5574 4558 5592
rect 4378 5516 4444 5574
rect 4500 5516 4558 5574
rect 4378 5498 4558 5516
rect 6102 5576 6282 5588
rect 6102 5518 6166 5576
rect 6222 5518 6282 5576
rect 6102 5494 6282 5518
rect 8010 5566 8190 5584
rect 8010 5508 8076 5566
rect 8132 5508 8190 5566
rect 9604 5566 9610 5618
rect 9662 5566 9672 5618
rect 9604 5562 9672 5566
rect 8010 5490 8190 5508
rect 10342 5452 10524 5474
rect 10342 5394 10414 5452
rect 10470 5394 10524 5452
rect 10342 5378 10524 5394
rect 11312 5456 11494 5468
rect 11312 5392 11370 5456
rect 11428 5392 11494 5456
rect 11312 5372 11494 5392
rect 14016 5450 14198 5462
rect 14016 5386 14072 5450
rect 14130 5386 14198 5450
rect 14016 5366 14198 5386
rect 14936 5442 15118 5458
rect 14936 5378 14992 5442
rect 15050 5378 15118 5442
rect 14936 5362 15118 5378
rect 17158 5428 17338 5444
rect 17158 5364 17226 5428
rect 17284 5364 17338 5428
rect 17158 5348 17338 5364
rect 2222 5146 2228 5198
rect 2280 5146 2290 5198
rect 17693 5175 17748 6338
rect 2222 5142 2290 5146
rect 9328 5120 9508 5142
rect 9328 5062 9388 5120
rect 9444 5062 9508 5120
rect 2520 5040 2700 5050
rect 9328 5046 9508 5062
rect 12208 5120 12390 5136
rect 12208 5056 12276 5120
rect 12334 5056 12390 5120
rect 2520 4982 2584 5040
rect 2640 4982 2700 5040
rect 2520 4956 2700 4982
rect 4378 5032 4558 5046
rect 4378 4974 4444 5032
rect 4500 4974 4558 5032
rect 4378 4952 4558 4974
rect 6092 5028 6272 5044
rect 12208 5040 12390 5056
rect 13070 5116 13252 5134
rect 13070 5052 13130 5116
rect 13188 5052 13252 5116
rect 6092 4970 6148 5028
rect 6204 4970 6272 5028
rect 6092 4950 6272 4970
rect 8004 5020 8184 5040
rect 13070 5038 13252 5052
rect 15866 5114 16048 5130
rect 15866 5050 15922 5114
rect 15980 5050 16048 5114
rect 17696 5098 17744 5175
rect 15866 5036 16048 5050
rect 17548 5050 17744 5098
rect 8004 4962 8064 5020
rect 8120 4962 8184 5020
rect 8004 4946 8184 4962
rect 17548 4998 17556 5050
rect 17608 4998 17612 5050
rect 17548 4942 17612 4998
rect 17162 4880 17342 4894
rect 17162 4816 17220 4880
rect 17278 4816 17342 4880
rect 9632 4744 9700 4802
rect 17162 4798 17342 4816
rect 9632 4692 9638 4744
rect 9690 4692 9700 4744
rect 9632 4566 9700 4692
rect 9632 4512 9640 4566
rect 9692 4512 9700 4566
rect 9632 4502 9700 4512
rect 9934 4580 10114 4594
rect 9934 4522 9988 4580
rect 10044 4522 10114 4580
rect 9934 4498 10114 4522
rect 11828 4578 12010 4592
rect 11828 4514 11894 4578
rect 11952 4514 12010 4578
rect 11828 4496 12010 4514
rect 13630 4574 13812 4590
rect 13630 4510 13698 4574
rect 13756 4510 13812 4574
rect 13630 4494 13812 4510
rect 15560 4566 15742 4584
rect 15560 4502 15628 4566
rect 15686 4502 15742 4566
rect 15560 4488 15742 4502
rect 6082 3382 6354 3386
rect 6082 3320 6194 3382
rect 6254 3320 6354 3382
rect 6082 3292 6354 3320
rect 24252 3138 24312 13230
rect 2192 3130 6198 3138
rect 2192 3078 6138 3130
rect 6190 3078 6198 3130
rect 6232 3136 24312 3138
rect 6232 3084 6238 3136
rect 6290 3084 24312 3136
rect 6232 3078 24312 3084
rect 2192 3072 6198 3078
rect 2192 1938 2260 3072
rect 6080 2828 6300 2842
rect 6080 2766 6176 2828
rect 6236 2766 6300 2828
rect 6080 2752 6300 2766
rect 2540 2318 2720 2336
rect 2540 2260 2604 2318
rect 2660 2260 2720 2318
rect 2540 2242 2720 2260
rect 4334 2314 4514 2330
rect 4334 2256 4392 2314
rect 4448 2256 4514 2314
rect 4334 2236 4514 2256
rect 6154 2310 6334 2326
rect 6154 2252 6220 2310
rect 6276 2252 6334 2310
rect 6154 2232 6334 2252
rect 7992 2308 8172 2322
rect 7992 2250 8060 2308
rect 8116 2250 8172 2308
rect 7992 2228 8172 2250
rect 9804 2312 9984 2320
rect 9804 2254 9870 2312
rect 9926 2254 9984 2312
rect 9804 2226 9984 2254
rect 11620 2302 11800 2318
rect 11620 2244 11686 2302
rect 11742 2244 11800 2302
rect 11620 2224 11800 2244
rect 13534 2300 13714 2312
rect 13534 2242 13594 2300
rect 13650 2242 13714 2300
rect 13534 2218 13714 2242
rect 15470 2296 15650 2310
rect 15470 2238 15534 2296
rect 15592 2238 15650 2296
rect 15470 2216 15650 2238
rect 2192 1886 2198 1938
rect 2250 1886 2260 1938
rect 2192 1882 2260 1886
rect 16306 1926 16376 3078
rect 16306 1874 16316 1926
rect 16368 1874 16376 1926
rect 16306 1866 16376 1874
rect 2538 1778 2718 1794
rect 2538 1720 2604 1778
rect 2660 1720 2718 1778
rect 2538 1700 2718 1720
rect 4334 1768 4514 1786
rect 4334 1710 4396 1768
rect 4452 1710 4514 1768
rect 4334 1692 4514 1710
rect 6190 1760 6370 1784
rect 6190 1702 6238 1760
rect 6294 1702 6370 1760
rect 6190 1690 6370 1702
rect 7994 1762 8174 1778
rect 7994 1704 8056 1762
rect 8112 1704 8174 1762
rect 7994 1684 8174 1704
rect 9846 1762 10026 1776
rect 9846 1704 9908 1762
rect 9964 1704 10026 1762
rect 9846 1682 10026 1704
rect 11616 1758 11796 1772
rect 11616 1700 11676 1758
rect 11732 1700 11796 1758
rect 11616 1678 11796 1700
rect 13504 1756 13684 1768
rect 13504 1698 13570 1756
rect 13626 1698 13684 1756
rect 13504 1674 13684 1698
rect 15452 1752 15632 1766
rect 15452 1694 15516 1752
rect 15574 1694 15632 1752
rect 15452 1672 15632 1694
rect 30230 820 30578 862
rect 30230 716 30332 820
rect 30436 716 30578 820
rect 30230 638 30578 716
<< via2 >>
rect 9540 17762 9600 17822
rect 4552 16570 4590 16614
rect 4590 16570 4608 16614
rect 4552 16558 4608 16570
rect 4976 16074 5034 16076
rect 4976 16020 5034 16074
rect 4746 15814 4808 15874
rect 9536 17218 9594 17278
rect 9514 16554 9552 16598
rect 9552 16554 9570 16598
rect 9514 16542 9570 16554
rect 9938 16058 9996 16060
rect 9938 16004 9996 16058
rect 9708 15798 9770 15858
rect 6712 15706 6780 15768
rect 4898 15270 4966 15332
rect 6130 15202 6198 15264
rect 9860 15254 9928 15316
rect 7114 15156 7182 15218
rect 4582 14986 4648 15052
rect 9544 14970 9610 15036
rect 5794 14654 5862 14716
rect 5012 14442 5078 14508
rect 4682 14244 4754 14314
rect 6350 14232 6418 14294
rect 6828 13856 6896 13918
rect 7916 14222 7984 14284
rect 4884 13700 4956 13770
rect 5862 13692 5930 13754
rect 7656 13676 7724 13738
rect 4576 13318 4648 13384
rect 5984 13390 6052 13450
rect 7136 13316 7204 13378
rect 5996 12856 6064 12916
rect 4990 12778 5062 12844
rect 4634 12576 4708 12642
rect 6280 12370 6348 12432
rect 4906 12034 4980 12100
rect 4560 11756 4640 11820
rect 6002 11830 6070 11892
rect 4994 11214 5074 11278
rect 4626 11010 4706 11074
rect 9974 14426 10040 14492
rect 9644 14228 9716 14298
rect 10756 14638 10824 14700
rect 16430 16660 16498 16722
rect 17188 16652 17256 16714
rect 18078 16654 18146 16716
rect 18686 16650 18754 16712
rect 19444 16642 19512 16704
rect 20334 16644 20402 16706
rect 21450 16644 21518 16706
rect 22208 16636 22276 16698
rect 23098 16638 23166 16700
rect 16410 16122 16478 16184
rect 17196 16112 17264 16174
rect 18076 16112 18144 16174
rect 18666 16112 18734 16174
rect 19452 16102 19520 16164
rect 20332 16102 20400 16164
rect 21430 16106 21498 16168
rect 22216 16096 22284 16158
rect 23096 16096 23164 16158
rect 11674 15690 11742 15752
rect 11092 15186 11160 15248
rect 12076 15140 12144 15202
rect 24400 14810 24462 14870
rect 9846 13684 9918 13754
rect 27000 14646 27122 14766
rect 11312 14216 11380 14278
rect 11790 13840 11858 13902
rect 12878 14206 12946 14268
rect 10824 13676 10892 13738
rect 9538 13302 9610 13368
rect 10946 13374 11014 13434
rect 12618 13660 12686 13722
rect 12098 13300 12166 13362
rect 10958 12840 11026 12900
rect 9952 12762 10024 12828
rect 9596 12560 9670 12626
rect 11242 12354 11310 12416
rect 9868 12018 9942 12084
rect 9522 11740 9602 11804
rect 10964 11814 11032 11876
rect 9956 11198 10036 11262
rect 9588 10994 9668 11058
rect 23992 14258 24054 14318
rect 4904 10476 4984 10540
rect 9866 10460 9946 10524
rect 6226 6580 6282 6638
rect 27550 14372 27682 14492
rect 6170 6030 6226 6088
rect 9974 5936 10032 6000
rect 11866 5934 11924 5998
rect 13652 5924 13710 5988
rect 15534 5928 15592 5992
rect 2564 5520 2620 5578
rect 4444 5516 4500 5574
rect 6166 5518 6222 5576
rect 8076 5508 8132 5566
rect 10414 5394 10470 5452
rect 11370 5392 11428 5456
rect 14072 5386 14130 5450
rect 14992 5378 15050 5442
rect 17226 5364 17284 5428
rect 9388 5062 9444 5120
rect 12276 5056 12334 5120
rect 2584 4982 2640 5040
rect 4444 4974 4500 5032
rect 13130 5052 13188 5116
rect 6148 4970 6204 5028
rect 15922 5050 15980 5114
rect 8064 4962 8120 5020
rect 17220 4816 17278 4880
rect 9988 4522 10044 4580
rect 11894 4514 11952 4578
rect 13698 4510 13756 4574
rect 15628 4502 15686 4566
rect 6194 3320 6254 3382
rect 6176 2766 6236 2828
rect 2604 2260 2660 2318
rect 4392 2256 4448 2314
rect 6220 2252 6276 2310
rect 8060 2250 8116 2308
rect 9870 2254 9926 2312
rect 11686 2244 11742 2302
rect 13594 2242 13650 2300
rect 15534 2238 15592 2296
rect 2604 1720 2656 1778
rect 2656 1720 2660 1778
rect 4396 1710 4452 1768
rect 6238 1702 6294 1760
rect 8056 1704 8112 1762
rect 9908 1704 9964 1762
rect 11676 1700 11732 1758
rect 13570 1698 13626 1756
rect 15516 1694 15574 1752
rect 30332 716 30436 820
<< metal3 >>
rect 814 17848 23871 17936
rect 814 17780 996 17848
rect 1066 17822 23871 17848
rect 1066 17780 9540 17822
rect 814 17762 9540 17780
rect 9600 17762 23871 17822
rect 814 17722 23871 17762
rect 18799 17720 19013 17722
rect 200 17278 13306 17330
rect 200 17218 9536 17278
rect 9594 17218 13306 17278
rect 200 17104 13306 17218
rect 200 16942 322 17104
rect 474 17038 13306 17104
rect 474 17022 21152 17038
rect 474 16942 23276 17022
rect 200 16810 23276 16942
rect 200 16808 13306 16810
rect 4036 16628 4280 16808
rect 4036 16614 4844 16628
rect 4036 16558 4552 16614
rect 4608 16558 4844 16614
rect 4036 16536 4844 16558
rect 4036 15884 4280 16536
rect 4880 16076 5584 16082
rect 4880 16020 4976 16076
rect 5034 16020 5584 16076
rect 4880 15994 5584 16020
rect 5342 15912 5584 15994
rect 4036 15874 4938 15884
rect 4036 15814 4746 15874
rect 4808 15814 4938 15874
rect 4036 15792 4938 15814
rect 4036 15066 4280 15792
rect 5340 15344 5584 15912
rect 4834 15332 5584 15344
rect 4834 15270 4898 15332
rect 4966 15270 5584 15332
rect 6320 15780 6502 16808
rect 6320 15768 6896 15780
rect 6320 15706 6712 15768
rect 6780 15706 6896 15768
rect 6320 15684 6896 15706
rect 6320 15278 6502 15684
rect 4834 15256 5584 15270
rect 4036 15052 4900 15066
rect 4036 14986 4582 15052
rect 4648 14986 4900 15052
rect 4036 14974 4900 14986
rect 4036 14324 4280 14974
rect 5340 14738 5584 15256
rect 6088 15264 6502 15278
rect 6088 15202 6130 15264
rect 6198 15202 6502 15264
rect 6088 15180 6502 15202
rect 5340 14716 6026 14738
rect 5340 14654 5794 14716
rect 5862 14654 6026 14716
rect 5340 14642 6026 14654
rect 5340 14522 5584 14642
rect 4942 14508 5584 14522
rect 4942 14442 5012 14508
rect 5078 14442 5584 14508
rect 4942 14434 5584 14442
rect 4036 14314 4880 14324
rect 4036 14244 4682 14314
rect 4754 14244 4880 14314
rect 4036 14232 4880 14244
rect 4036 13404 4280 14232
rect 5340 13776 5584 14434
rect 6320 14433 6502 15180
rect 7050 15218 7552 15236
rect 7050 15156 7114 15218
rect 7182 15156 7552 15218
rect 7050 15140 7552 15156
rect 6321 14430 6502 14433
rect 6321 14334 6684 14430
rect 6321 14328 6502 14334
rect 6320 14294 6502 14328
rect 6320 14232 6350 14294
rect 6418 14232 6502 14294
rect 6320 14213 6502 14232
rect 6589 13938 6684 14334
rect 6584 13918 6948 13938
rect 6584 13856 6828 13918
rect 6896 13856 6948 13918
rect 6584 13846 6948 13856
rect 4822 13772 5584 13776
rect 4822 13770 6086 13772
rect 4822 13700 4884 13770
rect 4956 13754 6086 13770
rect 4956 13700 5862 13754
rect 4822 13692 5862 13700
rect 5930 13692 6086 13754
rect 4822 13688 6086 13692
rect 5340 13676 6086 13688
rect 4036 13384 4884 13404
rect 4036 13318 4576 13384
rect 4648 13318 4884 13384
rect 4036 13312 4884 13318
rect 4036 12658 4280 13312
rect 5340 12928 5584 13676
rect 6589 13470 6684 13846
rect 5948 13450 6684 13470
rect 5948 13390 5984 13450
rect 6052 13390 6684 13450
rect 7348 13752 7552 15140
rect 7838 14284 8072 16808
rect 8940 16772 9242 16808
rect 11224 16772 11464 16808
rect 12742 16772 13034 16808
rect 7838 14222 7916 14284
rect 7984 14222 8072 14284
rect 7838 14188 8072 14222
rect 8998 16612 9242 16772
rect 8998 16598 9806 16612
rect 8998 16542 9514 16598
rect 9570 16542 9806 16598
rect 8998 16520 9806 16542
rect 8998 15868 9242 16520
rect 9842 16060 10546 16066
rect 9842 16004 9938 16060
rect 9996 16004 10546 16060
rect 9842 15978 10546 16004
rect 10304 15896 10546 15978
rect 8998 15858 9900 15868
rect 8998 15798 9708 15858
rect 9770 15798 9900 15858
rect 8998 15776 9900 15798
rect 8998 15050 9242 15776
rect 10302 15328 10546 15896
rect 9796 15316 10546 15328
rect 9796 15254 9860 15316
rect 9928 15254 10546 15316
rect 11282 15764 11464 16772
rect 11282 15752 11858 15764
rect 11282 15690 11674 15752
rect 11742 15690 11858 15752
rect 11282 15668 11858 15690
rect 11282 15262 11464 15668
rect 9796 15240 10546 15254
rect 8998 15036 9862 15050
rect 8998 14970 9544 15036
rect 9610 14970 9862 15036
rect 8998 14958 9862 14970
rect 8998 14308 9242 14958
rect 10302 14722 10546 15240
rect 11050 15248 11464 15262
rect 11050 15186 11092 15248
rect 11160 15186 11464 15248
rect 11050 15164 11464 15186
rect 10302 14700 10988 14722
rect 10302 14638 10756 14700
rect 10824 14638 10988 14700
rect 10302 14626 10988 14638
rect 10302 14506 10546 14626
rect 9904 14492 10546 14506
rect 9904 14426 9974 14492
rect 10040 14426 10546 14492
rect 9904 14418 10546 14426
rect 8998 14298 9842 14308
rect 8998 14228 9644 14298
rect 9716 14228 9842 14298
rect 8998 14216 9842 14228
rect 7348 13738 7746 13752
rect 7348 13676 7656 13738
rect 7724 13676 7746 13738
rect 7348 13656 7746 13676
rect 7348 13394 7552 13656
rect 5948 13378 6684 13390
rect 5340 12916 6098 12928
rect 5340 12856 5996 12916
rect 6064 12856 6098 12916
rect 5340 12854 6098 12856
rect 4926 12844 6098 12854
rect 4926 12778 4990 12844
rect 5062 12832 6098 12844
rect 5062 12778 5584 12832
rect 4926 12766 5584 12778
rect 4036 12642 4952 12658
rect 4036 12576 4634 12642
rect 4708 12576 4952 12642
rect 4036 12566 4952 12576
rect 4036 11840 4280 12566
rect 5340 12110 5584 12766
rect 6589 12454 6684 13378
rect 7092 13378 7552 13394
rect 7092 13316 7136 13378
rect 7204 13316 7552 13378
rect 7092 13298 7552 13316
rect 6193 12432 6684 12454
rect 6193 12370 6280 12432
rect 6348 12370 6684 12432
rect 6193 12359 6684 12370
rect 4850 12100 5584 12110
rect 4850 12034 4906 12100
rect 4980 12034 5584 12100
rect 4850 12022 5584 12034
rect 5340 11906 5584 12022
rect 5340 11892 6100 11906
rect 4036 11820 4838 11840
rect 4036 11756 4560 11820
rect 4640 11756 4838 11820
rect 4036 11748 4838 11756
rect 5340 11830 6002 11892
rect 6070 11830 6100 11892
rect 5340 11810 6100 11830
rect 4036 11090 4280 11748
rect 5340 11294 5584 11810
rect 4936 11278 5584 11294
rect 4936 11214 4994 11278
rect 5074 11214 5584 11278
rect 4936 11200 5584 11214
rect 4036 11074 4904 11090
rect 4036 11010 4626 11074
rect 4706 11010 4904 11074
rect 4036 10998 4904 11010
rect 4036 10996 4280 10998
rect 5340 10554 5584 11200
rect 4852 10540 5584 10554
rect 4852 10476 4904 10540
rect 4984 10476 5584 10540
rect 4852 10448 5584 10476
rect 5340 9882 5584 10448
rect 7348 9882 7552 13298
rect 8998 13388 9242 14216
rect 10302 13760 10546 14418
rect 11282 14417 11464 15164
rect 12012 15202 12514 15220
rect 12012 15140 12076 15202
rect 12144 15140 12514 15202
rect 12012 15124 12514 15140
rect 11283 14414 11464 14417
rect 11283 14318 11646 14414
rect 11283 14312 11464 14318
rect 11282 14278 11464 14312
rect 11282 14216 11312 14278
rect 11380 14216 11464 14278
rect 11282 14197 11464 14216
rect 11551 13922 11646 14318
rect 11546 13902 11910 13922
rect 11546 13840 11790 13902
rect 11858 13840 11910 13902
rect 11546 13830 11910 13840
rect 9784 13756 10546 13760
rect 9784 13754 11048 13756
rect 9784 13684 9846 13754
rect 9918 13738 11048 13754
rect 9918 13684 10824 13738
rect 9784 13676 10824 13684
rect 10892 13676 11048 13738
rect 9784 13672 11048 13676
rect 10302 13660 11048 13672
rect 8998 13368 9846 13388
rect 8998 13302 9538 13368
rect 9610 13302 9846 13368
rect 8998 13296 9846 13302
rect 8998 12642 9242 13296
rect 10302 12912 10546 13660
rect 11551 13454 11646 13830
rect 10910 13434 11646 13454
rect 10910 13374 10946 13434
rect 11014 13374 11646 13434
rect 12310 13736 12514 15124
rect 12800 14268 13034 16772
rect 15198 15406 15426 16810
rect 16340 16722 16568 16810
rect 16340 16660 16430 16722
rect 16498 16660 16568 16722
rect 16340 16652 16568 16660
rect 17108 16714 17336 16810
rect 17108 16652 17188 16714
rect 17256 16652 17336 16714
rect 17108 16642 17336 16652
rect 17998 16716 18226 16810
rect 18452 16800 20542 16810
rect 17998 16654 18078 16716
rect 18146 16654 18226 16716
rect 17998 16638 18226 16654
rect 18596 16712 18824 16800
rect 18596 16650 18686 16712
rect 18754 16650 18824 16712
rect 18596 16642 18824 16650
rect 19364 16704 19592 16800
rect 19364 16642 19444 16704
rect 19512 16642 19592 16704
rect 19364 16632 19592 16642
rect 20254 16706 20482 16800
rect 20990 16794 23276 16810
rect 20254 16644 20334 16706
rect 20402 16644 20482 16706
rect 20254 16628 20482 16644
rect 21360 16706 21588 16794
rect 21360 16644 21450 16706
rect 21518 16644 21588 16706
rect 21360 16636 21588 16644
rect 22128 16698 22356 16794
rect 22128 16636 22208 16698
rect 22276 16636 22356 16698
rect 22128 16626 22356 16636
rect 23018 16700 23246 16794
rect 23018 16638 23098 16700
rect 23166 16638 23246 16700
rect 23018 16622 23246 16638
rect 16333 16184 16547 16199
rect 16333 16122 16410 16184
rect 16478 16122 16547 16184
rect 16333 16027 16547 16122
rect 17127 16174 17341 16185
rect 17127 16112 17196 16174
rect 17264 16112 17341 16174
rect 17127 16027 17341 16112
rect 17993 16174 18207 16191
rect 17993 16112 18076 16174
rect 18144 16112 18207 16174
rect 17993 16027 18207 16112
rect 18589 16174 18803 16189
rect 18589 16112 18666 16174
rect 18734 16112 18803 16174
rect 16197 16018 18300 16027
rect 16197 16017 18510 16018
rect 18589 16017 18803 16112
rect 19383 16164 19597 16175
rect 19383 16102 19452 16164
rect 19520 16102 19597 16164
rect 19383 16017 19597 16102
rect 20249 16164 20463 16181
rect 20249 16102 20332 16164
rect 20400 16102 20463 16164
rect 20249 16017 20463 16102
rect 21353 16168 21567 16183
rect 21353 16106 21430 16168
rect 21498 16106 21567 16168
rect 21353 16017 21567 16106
rect 16197 16011 21567 16017
rect 22147 16158 22361 16169
rect 22147 16096 22216 16158
rect 22284 16096 22361 16158
rect 22147 16011 22361 16096
rect 23013 16158 23227 16175
rect 23013 16096 23096 16158
rect 23164 16096 23227 16158
rect 23013 16027 23227 16096
rect 23657 16027 23871 17722
rect 22627 16011 23871 16027
rect 16197 16010 21710 16011
rect 21790 16010 21966 16011
rect 16197 16006 21966 16010
rect 22094 16006 23871 16011
rect 16197 15896 23871 16006
rect 16197 15813 23874 15896
rect 18292 15803 23874 15813
rect 20597 15797 23874 15803
rect 23270 15794 23874 15797
rect 15198 15178 24536 15406
rect 24310 15150 24536 15178
rect 24310 14870 24538 15150
rect 24310 14810 24400 14870
rect 24462 14810 24538 14870
rect 24310 14790 24538 14810
rect 26956 14766 27174 14788
rect 26956 14646 27000 14766
rect 27122 14646 27174 14766
rect 26956 14604 27174 14646
rect 27512 14492 27730 14510
rect 27512 14372 27550 14492
rect 27682 14372 27730 14492
rect 27512 14336 27730 14372
rect 12800 14206 12878 14268
rect 12946 14206 13034 14268
rect 12800 14172 13034 14206
rect 23852 14318 24212 14334
rect 23852 14258 23992 14318
rect 24054 14258 24212 14318
rect 23852 14128 24212 14258
rect 23852 13946 24204 14128
rect 12310 13722 12708 13736
rect 12310 13660 12618 13722
rect 12686 13660 12708 13722
rect 12310 13640 12708 13660
rect 15110 13726 24204 13946
rect 12310 13378 12514 13640
rect 10910 13362 11646 13374
rect 10302 12900 11060 12912
rect 10302 12840 10958 12900
rect 11026 12840 11060 12900
rect 10302 12838 11060 12840
rect 9888 12828 11060 12838
rect 9888 12762 9952 12828
rect 10024 12816 11060 12828
rect 10024 12762 10546 12816
rect 9888 12750 10546 12762
rect 8998 12626 9914 12642
rect 8998 12560 9596 12626
rect 9670 12560 9914 12626
rect 8998 12550 9914 12560
rect 8998 11824 9242 12550
rect 10302 12094 10546 12750
rect 11551 12438 11646 13362
rect 12054 13362 12514 13378
rect 12054 13300 12098 13362
rect 12166 13300 12514 13362
rect 12054 13282 12514 13300
rect 11155 12416 11646 12438
rect 11155 12354 11242 12416
rect 11310 12354 11646 12416
rect 11155 12343 11646 12354
rect 9812 12084 10546 12094
rect 9812 12018 9868 12084
rect 9942 12018 10546 12084
rect 9812 12006 10546 12018
rect 10302 11890 10546 12006
rect 10302 11876 11062 11890
rect 8998 11804 9800 11824
rect 8998 11740 9522 11804
rect 9602 11740 9800 11804
rect 8998 11732 9800 11740
rect 10302 11814 10964 11876
rect 11032 11814 11062 11876
rect 10302 11794 11062 11814
rect 8998 11074 9242 11732
rect 10302 11278 10546 11794
rect 9898 11262 10546 11278
rect 9898 11198 9956 11262
rect 10036 11198 10546 11262
rect 9898 11184 10546 11198
rect 8998 11058 9866 11074
rect 8998 10994 9588 11058
rect 9668 10994 9866 11058
rect 8998 10982 9866 10994
rect 8998 10980 9242 10982
rect 10302 10538 10546 11184
rect 9814 10524 10546 10538
rect 9814 10460 9866 10524
rect 9946 10460 10546 10524
rect 9814 10432 10546 10460
rect 800 9864 8764 9882
rect 10302 9864 10546 10432
rect 12310 9864 12514 13282
rect 15110 13586 24208 13726
rect 15110 9890 15470 13586
rect 13142 9864 15470 9890
rect 800 9724 15470 9864
rect 800 9562 994 9724
rect 1146 9562 15470 9724
rect 800 9530 15470 9562
rect 800 9376 13253 9530
rect 6108 6638 6646 6736
rect 6108 6580 6226 6638
rect 6282 6580 6646 6638
rect 6108 6556 6646 6580
rect 372 6088 6274 6108
rect 372 6074 6170 6088
rect 372 5986 392 6074
rect 498 6030 6170 6074
rect 6226 6030 6274 6088
rect 498 5986 6274 6030
rect 372 5954 6274 5986
rect 6466 5814 6646 6556
rect 8852 6042 17338 6222
rect 8852 5814 9032 6042
rect 802 5774 9032 5814
rect 802 5670 936 5774
rect 1052 5670 9032 5774
rect 802 5634 9032 5670
rect 2512 5578 2692 5634
rect 2512 5520 2564 5578
rect 2620 5520 2692 5578
rect 2512 5506 2692 5520
rect 4378 5574 4558 5634
rect 4378 5516 4444 5574
rect 4500 5516 4558 5574
rect 4378 5496 4558 5516
rect 6104 5576 6284 5634
rect 6104 5518 6166 5576
rect 6222 5518 6284 5576
rect 6104 5490 6284 5518
rect 8010 5566 8190 5634
rect 8010 5508 8076 5566
rect 8132 5508 8190 5566
rect 8010 5492 8190 5508
rect 9328 5120 9508 6042
rect 9908 6000 10088 6042
rect 9908 5936 9974 6000
rect 10032 5936 10088 6000
rect 9908 5924 10088 5936
rect 11798 5998 11978 6042
rect 11798 5934 11866 5998
rect 11924 5934 11978 5998
rect 11798 5918 11978 5934
rect 10172 5456 11640 5480
rect 10172 5452 11370 5456
rect 10172 5394 10414 5452
rect 10470 5394 11370 5452
rect 10172 5392 11370 5394
rect 11428 5392 11640 5456
rect 10172 5300 11640 5392
rect 9328 5062 9388 5120
rect 9444 5062 9508 5120
rect 2520 5040 2700 5048
rect 9328 5046 9508 5062
rect 2520 4982 2584 5040
rect 2640 4982 2700 5040
rect 2520 4850 2700 4982
rect 4380 5032 4560 5046
rect 4380 4974 4444 5032
rect 4500 4974 4560 5032
rect 4380 4850 4560 4974
rect 6092 5028 6272 5038
rect 6092 4970 6148 5028
rect 6204 4970 6272 5028
rect 6092 4850 6272 4970
rect 8002 5020 8182 5042
rect 8002 4962 8064 5020
rect 8120 4962 8182 5020
rect 8002 4850 8182 4962
rect 198 4814 9032 4850
rect 198 4710 330 4814
rect 446 4710 9032 4814
rect 198 4670 9032 4710
rect 8852 4496 9032 4670
rect 9932 4580 10112 4598
rect 9932 4522 9988 4580
rect 10044 4522 10112 4580
rect 8852 4376 9034 4496
rect 9932 4376 10112 4522
rect 10776 4376 10956 5300
rect 12630 5216 12810 6042
rect 13570 5988 13750 6042
rect 13570 5924 13652 5988
rect 13710 5924 13750 5988
rect 13570 5916 13750 5924
rect 15464 5992 15644 6042
rect 15866 6036 16046 6042
rect 15464 5928 15534 5992
rect 15592 5928 15644 5992
rect 15464 5912 15644 5928
rect 13828 5450 15242 5458
rect 13828 5386 14072 5450
rect 14130 5442 15242 5450
rect 14130 5386 14992 5442
rect 13828 5378 14992 5386
rect 15050 5378 15242 5442
rect 13828 5278 15242 5378
rect 12044 5120 13380 5216
rect 12044 5056 12276 5120
rect 12334 5116 13380 5120
rect 12334 5056 13130 5116
rect 12044 5052 13130 5056
rect 13188 5052 13380 5116
rect 12044 5036 13380 5052
rect 11828 4578 12008 4594
rect 11828 4514 11894 4578
rect 11952 4514 12008 4578
rect 11828 4376 12008 4514
rect 13636 4574 13816 4588
rect 13636 4510 13698 4574
rect 13756 4510 13816 4574
rect 13636 4376 13816 4510
rect 14502 4376 14682 5278
rect 15866 5130 16046 5878
rect 17158 5428 17338 6042
rect 17158 5364 17226 5428
rect 17284 5364 17338 5428
rect 17158 5354 17338 5364
rect 15866 5114 16048 5130
rect 15866 5050 15922 5114
rect 15980 5050 16048 5114
rect 15866 5034 16048 5050
rect 17162 4880 17342 4888
rect 17162 4816 17220 4880
rect 17278 4816 17342 4880
rect 15556 4566 15736 4582
rect 15556 4502 15628 4566
rect 15686 4502 15736 4566
rect 15556 4376 15736 4502
rect 17162 4376 17342 4816
rect 8852 4196 17342 4376
rect 6082 3382 6656 3408
rect 6082 3320 6194 3382
rect 6254 3320 6656 3382
rect 6082 3228 6656 3320
rect 294 2828 6298 2858
rect 294 2808 6176 2828
rect 294 2714 384 2808
rect 484 2766 6176 2808
rect 6236 2766 6298 2828
rect 484 2714 6298 2766
rect 294 2664 6298 2714
rect 6476 2554 6656 3228
rect 794 2518 16220 2554
rect 794 2410 936 2518
rect 1068 2410 16220 2518
rect 794 2374 16220 2410
rect 2540 2318 2720 2374
rect 2540 2260 2604 2318
rect 2660 2260 2720 2318
rect 2540 2244 2720 2260
rect 4336 2314 4516 2374
rect 4336 2256 4392 2314
rect 4448 2256 4516 2314
rect 4336 2236 4516 2256
rect 6154 2310 6334 2374
rect 6154 2252 6220 2310
rect 6276 2252 6334 2310
rect 6154 2234 6334 2252
rect 7992 2308 8172 2374
rect 7992 2250 8060 2308
rect 8116 2250 8172 2308
rect 7992 2232 8172 2250
rect 9804 2312 9984 2374
rect 9804 2254 9870 2312
rect 9926 2254 9984 2312
rect 9804 2226 9984 2254
rect 11620 2302 11800 2374
rect 11620 2244 11686 2302
rect 11742 2244 11800 2302
rect 11620 2224 11800 2244
rect 13534 2300 13714 2374
rect 13534 2242 13594 2300
rect 13650 2242 13714 2300
rect 15470 2296 15650 2374
rect 15470 2280 15534 2296
rect 13534 2224 13714 2242
rect 15468 2238 15534 2280
rect 15592 2238 15650 2296
rect 15468 2216 15650 2238
rect 2542 1778 2722 1790
rect 2542 1720 2604 1778
rect 2660 1720 2722 1778
rect 2542 1590 2722 1720
rect 4334 1768 4514 1792
rect 4334 1710 4396 1768
rect 4452 1710 4514 1768
rect 4334 1590 4514 1710
rect 6190 1760 6370 1784
rect 6190 1702 6238 1760
rect 6294 1702 6370 1760
rect 6190 1590 6370 1702
rect 7996 1762 8176 1780
rect 7996 1704 8056 1762
rect 8112 1704 8176 1762
rect 7996 1590 8176 1704
rect 9844 1762 10024 1774
rect 9844 1704 9908 1762
rect 9964 1704 10024 1762
rect 9844 1590 10024 1704
rect 11616 1758 11796 1780
rect 11616 1700 11676 1758
rect 11732 1700 11796 1758
rect 11616 1590 11796 1700
rect 13506 1756 13686 1772
rect 13506 1698 13570 1756
rect 13626 1698 13686 1756
rect 13506 1590 13686 1698
rect 15456 1752 15636 1766
rect 15456 1694 15516 1752
rect 15574 1694 15636 1752
rect 15456 1590 15636 1694
rect 210 1548 15636 1590
rect 210 1438 336 1548
rect 456 1438 15636 1548
rect 210 1410 15636 1438
rect 30230 820 30578 862
rect 30230 716 30332 820
rect 30436 716 30578 820
rect 30230 638 30578 716
<< via3 >>
rect 996 17780 1066 17848
rect 322 16942 474 17104
rect 27000 14646 27122 14766
rect 27550 14372 27682 14492
rect 994 9562 1146 9724
rect 392 5986 498 6074
rect 936 5670 1052 5774
rect 330 4710 446 4814
rect 384 2714 484 2808
rect 936 2410 1068 2518
rect 336 1438 456 1548
rect 30332 716 30436 820
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 200 17104 600 44152
rect 200 16942 322 17104
rect 474 16942 600 17104
rect 200 6074 600 16942
rect 200 5986 392 6074
rect 498 5986 600 6074
rect 200 4814 600 5986
rect 200 4710 330 4814
rect 446 4710 600 4814
rect 200 2808 600 4710
rect 200 2714 384 2808
rect 484 2714 600 2808
rect 200 1548 600 2714
rect 200 1438 336 1548
rect 456 1438 600 1548
rect 200 1000 600 1438
rect 800 17848 1200 44152
rect 800 17780 996 17848
rect 1066 17780 1200 17848
rect 800 9724 1200 17780
rect 27110 14788 27170 45152
rect 26956 14766 27174 14788
rect 26956 14646 27000 14766
rect 27122 14646 27174 14766
rect 26956 14604 27174 14646
rect 27662 14510 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 27512 14492 27730 14510
rect 27512 14372 27550 14492
rect 27682 14372 27730 14492
rect 27512 14336 27730 14372
rect 800 9562 994 9724
rect 1146 9562 1200 9724
rect 800 5774 1200 9562
rect 800 5670 936 5774
rect 1052 5670 1200 5774
rect 800 2518 1200 5670
rect 800 2410 936 2518
rect 1068 2410 1200 2518
rect 800 1000 1200 2410
rect 30230 820 30578 862
rect 30230 716 30332 820
rect 30436 716 30578 820
rect 30230 638 30578 716
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 0 30542 638
use CLA  CLA_0
timestamp 1754418791
transform 1 0 4568 0 1 15292
box -138 -4838 3664 1342
use CLA  CLA_1
timestamp 1754418791
transform 1 0 9530 0 1 15276
box -138 -4838 3664 1342
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 3278 0 -1 2288
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_1
timestamp 1723858470
transform -1 0 5148 0 -1 2284
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_2
timestamp 1723858470
transform -1 0 6964 0 -1 2280
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_3
timestamp 1723858470
transform -1 0 8834 0 -1 2276
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_4
timestamp 1723858470
transform -1 0 16204 0 -1 2262
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_5
timestamp 1723858470
transform -1 0 14334 0 -1 2266
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_6
timestamp 1723858470
transform -1 0 10648 0 -1 2274
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_7
timestamp 1723858470
transform -1 0 12518 0 -1 2270
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_8
timestamp 1723858470
transform -1 0 8864 0 -1 5536
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_9
timestamp 1723858470
transform -1 0 6994 0 -1 5540
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_10
timestamp 1723858470
transform -1 0 3308 0 -1 5548
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_11
timestamp 1723858470
transform -1 0 5178 0 -1 5544
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_12
timestamp 1723858470
transform -1 0 12560 0 -1 5964
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_13
timestamp 1723858470
transform -1 0 10690 0 -1 5968
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_14
timestamp 1723858470
transform -1 0 14376 0 -1 5960
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_15
timestamp 1723858470
transform -1 0 16246 0 -1 5956
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_16
timestamp 1723858470
transform -1 0 12588 0 -1 5090
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_17
timestamp 1723858470
transform -1 0 10718 0 -1 5094
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_18
timestamp 1723858470
transform -1 0 14404 0 -1 5086
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_19
timestamp 1723858470
transform -1 0 16274 0 -1 5082
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 6358 0 -1 3340
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1723858470
transform -1 0 6388 0 -1 6600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1723858470
transform -1 0 9706 0 -1 17794
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1723858470
transform 1 0 16336 0 1 16150
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_4
timestamp 1723858470
transform 1 0 17104 0 1 16140
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_5
timestamp 1723858470
transform 1 0 17978 0 1 16142
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_6
timestamp 1723858470
transform 1 0 18592 0 1 16140
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_7
timestamp 1723858470
transform 1 0 19360 0 1 16130
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_8
timestamp 1723858470
transform 1 0 20234 0 1 16132
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_9
timestamp 1723858470
transform 1 0 21356 0 1 16134
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_10
timestamp 1723858470
transform 1 0 22124 0 1 16124
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_11
timestamp 1723858470
transform 1 0 22998 0 1 16126
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sky130_fd_sc_hd__mux2_1_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 17630 0 -1 5396
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 23484 0 1 14288
box -38 -48 1970 592
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
rlabel metal1 s 3676 1692 5148 1788 5 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 3676 2236 5148 2332 5 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4796 1992 4854 2001 5 B
port 2 nsew signal input
rlabel metal1 s 3964 1964 4854 1992 5 B
port 2 nsew signal input
rlabel metal1 s 4796 1955 4854 1964 5 B
port 2 nsew signal input
rlabel metal1 s 4424 1992 4482 2001 5 B
port 2 nsew signal input
rlabel metal1 s 4424 1955 4482 1964 5 B
port 2 nsew signal input
rlabel metal1 s 3964 1992 4022 2001 5 B
port 2 nsew signal input
rlabel metal1 s 3964 1955 4022 1964 5 B
port 2 nsew signal input
rlabel locali s 3937 1931 4021 1995 5 B
port 2 nsew signal input
rlabel locali s 4436 1931 4508 1997 5 B
port 2 nsew signal input
rlabel metal1 s 4888 2060 4946 2069 5 A
port 1 nsew signal input
rlabel metal1 s 3872 2032 4946 2060 5 A
port 1 nsew signal input
rlabel metal1 s 4888 2023 4946 2032 5 A
port 1 nsew signal input
rlabel metal1 s 4612 2060 4670 2069 5 A
port 1 nsew signal input
rlabel metal1 s 4612 2023 4670 2032 5 A
port 1 nsew signal input
rlabel metal1 s 4240 2060 4298 2069 5 A
port 1 nsew signal input
rlabel metal1 s 4240 2023 4298 2032 5 A
port 1 nsew signal input
rlabel metal1 s 3872 2060 3930 2069 5 A
port 1 nsew signal input
rlabel metal1 s 3872 2023 3930 2032 5 A
port 1 nsew signal input
rlabel locali s 3883 2029 3971 2077 5 A
port 1 nsew signal input
rlabel locali s 4223 2029 4298 2093 5 A
port 1 nsew signal input
rlabel locali s 4624 2012 4702 2078 5 A
port 1 nsew signal input
rlabel comment s 5148 2284 5148 2284 8 fa_1
flabel metal1 s 5084 1723 5118 1757 0 FreeSans 200 180 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 5084 2267 5118 2301 0 FreeSans 200 180 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel pwell s 5084 2267 5118 2301 0 FreeSans 200 180 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 5084 1723 5118 1757 0 FreeSans 200 180 0 0 VPB
port 6 nsew power bidirectional
flabel locali s 4808 1961 4842 1995 0 FreeSans 200 180 0 0 B
port 2 nsew signal input
flabel locali s 4900 2029 4934 2063 0 FreeSans 200 180 0 0 A
port 1 nsew signal input
flabel locali s 3700 1825 3734 1859 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 3700 1893 3734 1927 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 3700 1961 3734 1995 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 3700 2029 3734 2063 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 3700 2097 3734 2131 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 3700 2165 3734 2199 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 4068 1893 4102 1927 0 FreeSans 200 180 0 0 CIN
port 3 nsew signal input
flabel locali s 5084 2165 5118 2199 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 5084 1893 5118 1927 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 5084 1825 5118 1859 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
rlabel metal1 s 1806 1696 3278 1792 5 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 1806 2240 3278 2336 5 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2926 1996 2984 2005 5 B
port 2 nsew signal input
rlabel metal1 s 2094 1968 2984 1996 5 B
port 2 nsew signal input
rlabel metal1 s 2926 1959 2984 1968 5 B
port 2 nsew signal input
rlabel metal1 s 2554 1996 2612 2005 5 B
port 2 nsew signal input
rlabel metal1 s 2554 1959 2612 1968 5 B
port 2 nsew signal input
rlabel metal1 s 2094 1996 2152 2005 5 B
port 2 nsew signal input
rlabel metal1 s 2094 1959 2152 1968 5 B
port 2 nsew signal input
rlabel locali s 2067 1935 2151 1999 5 B
port 2 nsew signal input
rlabel locali s 2566 1935 2638 2001 5 B
port 2 nsew signal input
rlabel metal1 s 3018 2064 3076 2073 5 A
port 1 nsew signal input
rlabel metal1 s 2002 2036 3076 2064 5 A
port 1 nsew signal input
rlabel metal1 s 3018 2027 3076 2036 5 A
port 1 nsew signal input
rlabel metal1 s 2742 2064 2800 2073 5 A
port 1 nsew signal input
rlabel metal1 s 2742 2027 2800 2036 5 A
port 1 nsew signal input
rlabel metal1 s 2370 2064 2428 2073 5 A
port 1 nsew signal input
rlabel metal1 s 2370 2027 2428 2036 5 A
port 1 nsew signal input
rlabel metal1 s 2002 2064 2060 2073 5 A
port 1 nsew signal input
rlabel metal1 s 2002 2027 2060 2036 5 A
port 1 nsew signal input
rlabel locali s 2013 2033 2101 2081 5 A
port 1 nsew signal input
rlabel locali s 2353 2033 2428 2097 5 A
port 1 nsew signal input
rlabel locali s 2754 2016 2832 2082 5 A
port 1 nsew signal input
rlabel comment s 3278 2288 3278 2288 8 fa_1
flabel metal1 s 3214 1727 3248 1761 0 FreeSans 200 180 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 3214 2271 3248 2305 0 FreeSans 200 180 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel pwell s 3214 2271 3248 2305 0 FreeSans 200 180 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 3214 1727 3248 1761 0 FreeSans 200 180 0 0 VPB
port 6 nsew power bidirectional
flabel locali s 2938 1965 2972 1999 0 FreeSans 200 180 0 0 B
port 2 nsew signal input
flabel locali s 3030 2033 3064 2067 0 FreeSans 200 180 0 0 A
port 1 nsew signal input
flabel locali s 1830 1829 1864 1863 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 1830 1897 1864 1931 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 1830 1965 1864 1999 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 1830 2033 1864 2067 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 1830 2101 1864 2135 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 1830 2169 1864 2203 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 2198 1897 2232 1931 0 FreeSans 200 180 0 0 CIN
port 3 nsew signal input
flabel locali s 3214 2169 3248 2203 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 3214 1897 3248 1931 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 3214 1829 3248 1863 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
rlabel metal1 s 5492 1688 6964 1784 5 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 5492 2232 6964 2328 5 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 6612 1988 6670 1997 5 B
port 2 nsew signal input
rlabel metal1 s 5780 1960 6670 1988 5 B
port 2 nsew signal input
rlabel metal1 s 6612 1951 6670 1960 5 B
port 2 nsew signal input
rlabel metal1 s 6240 1988 6298 1997 5 B
port 2 nsew signal input
rlabel metal1 s 6240 1951 6298 1960 5 B
port 2 nsew signal input
rlabel metal1 s 5780 1988 5838 1997 5 B
port 2 nsew signal input
rlabel metal1 s 5780 1951 5838 1960 5 B
port 2 nsew signal input
rlabel locali s 5753 1927 5837 1991 5 B
port 2 nsew signal input
rlabel locali s 6252 1927 6324 1993 5 B
port 2 nsew signal input
rlabel metal1 s 6704 2056 6762 2065 5 A
port 1 nsew signal input
rlabel metal1 s 5688 2028 6762 2056 5 A
port 1 nsew signal input
rlabel metal1 s 6704 2019 6762 2028 5 A
port 1 nsew signal input
rlabel metal1 s 6428 2056 6486 2065 5 A
port 1 nsew signal input
rlabel metal1 s 6428 2019 6486 2028 5 A
port 1 nsew signal input
rlabel metal1 s 6056 2056 6114 2065 5 A
port 1 nsew signal input
rlabel metal1 s 6056 2019 6114 2028 5 A
port 1 nsew signal input
rlabel metal1 s 5688 2056 5746 2065 5 A
port 1 nsew signal input
rlabel metal1 s 5688 2019 5746 2028 5 A
port 1 nsew signal input
rlabel locali s 5699 2025 5787 2073 5 A
port 1 nsew signal input
rlabel locali s 6039 2025 6114 2089 5 A
port 1 nsew signal input
rlabel locali s 6440 2008 6518 2074 5 A
port 1 nsew signal input
rlabel comment s 6964 2280 6964 2280 8 fa_1
flabel metal1 s 6900 1719 6934 1753 0 FreeSans 200 180 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 6900 2263 6934 2297 0 FreeSans 200 180 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel pwell s 6900 2263 6934 2297 0 FreeSans 200 180 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 6900 1719 6934 1753 0 FreeSans 200 180 0 0 VPB
port 6 nsew power bidirectional
flabel locali s 6624 1957 6658 1991 0 FreeSans 200 180 0 0 B
port 2 nsew signal input
flabel locali s 6716 2025 6750 2059 0 FreeSans 200 180 0 0 A
port 1 nsew signal input
flabel locali s 5516 1821 5550 1855 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 5516 1889 5550 1923 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 5516 1957 5550 1991 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 5516 2025 5550 2059 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 5516 2093 5550 2127 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 5516 2161 5550 2195 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 5884 1889 5918 1923 0 FreeSans 200 180 0 0 CIN
port 3 nsew signal input
flabel locali s 6900 2161 6934 2195 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 6900 1889 6934 1923 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 6900 1821 6934 1855 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
rlabel metal1 s 7362 1684 8834 1780 5 VPWR
port 7 nsew power bidirectional abutment
rlabel metal1 s 7362 2228 8834 2324 5 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 8482 1984 8540 1993 5 B
port 2 nsew signal input
rlabel metal1 s 7650 1956 8540 1984 5 B
port 2 nsew signal input
rlabel metal1 s 8482 1947 8540 1956 5 B
port 2 nsew signal input
rlabel metal1 s 8110 1984 8168 1993 5 B
port 2 nsew signal input
rlabel metal1 s 8110 1947 8168 1956 5 B
port 2 nsew signal input
rlabel metal1 s 7650 1984 7708 1993 5 B
port 2 nsew signal input
rlabel metal1 s 7650 1947 7708 1956 5 B
port 2 nsew signal input
rlabel locali s 7623 1923 7707 1987 5 B
port 2 nsew signal input
rlabel locali s 8122 1923 8194 1989 5 B
port 2 nsew signal input
rlabel metal1 s 8574 2052 8632 2061 5 A
port 1 nsew signal input
rlabel metal1 s 7558 2024 8632 2052 5 A
port 1 nsew signal input
rlabel metal1 s 8574 2015 8632 2024 5 A
port 1 nsew signal input
rlabel metal1 s 8298 2052 8356 2061 5 A
port 1 nsew signal input
rlabel metal1 s 8298 2015 8356 2024 5 A
port 1 nsew signal input
rlabel metal1 s 7926 2052 7984 2061 5 A
port 1 nsew signal input
rlabel metal1 s 7926 2015 7984 2024 5 A
port 1 nsew signal input
rlabel metal1 s 7558 2052 7616 2061 5 A
port 1 nsew signal input
rlabel metal1 s 7558 2015 7616 2024 5 A
port 1 nsew signal input
rlabel locali s 7569 2021 7657 2069 5 A
port 1 nsew signal input
rlabel locali s 7909 2021 7984 2085 5 A
port 1 nsew signal input
rlabel locali s 8310 2004 8388 2070 5 A
port 1 nsew signal input
rlabel comment s 8834 2276 8834 2276 8 fa_1
flabel metal1 s 8770 1715 8804 1749 0 FreeSans 200 180 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 8770 2259 8804 2293 0 FreeSans 200 180 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel pwell s 8770 2259 8804 2293 0 FreeSans 200 180 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 8770 1715 8804 1749 0 FreeSans 200 180 0 0 VPB
port 6 nsew power bidirectional
flabel locali s 8494 1953 8528 1987 0 FreeSans 200 180 0 0 B
port 2 nsew signal input
flabel locali s 8586 2021 8620 2055 0 FreeSans 200 180 0 0 A
port 1 nsew signal input
flabel locali s 7386 1817 7420 1851 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 7386 1885 7420 1919 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 7386 1953 7420 1987 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 7386 2021 7420 2055 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 7386 2089 7420 2123 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 7386 2157 7420 2191 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 7754 1885 7788 1919 0 FreeSans 200 180 0 0 CIN
port 3 nsew signal input
flabel locali s 8770 2157 8804 2191 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 8770 1885 8804 1919 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 8770 1817 8804 1851 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 16140 1803 16174 1837 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 16140 1871 16174 1905 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 16140 2143 16174 2177 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 15124 1871 15158 1905 0 FreeSans 200 180 0 0 CIN
port 3 nsew signal input
flabel locali s 14756 2143 14790 2177 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 14756 2075 14790 2109 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 14756 2007 14790 2041 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 14756 1939 14790 1973 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 14756 1871 14790 1905 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 14756 1803 14790 1837 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 15956 2007 15990 2041 0 FreeSans 200 180 0 0 A
port 1 nsew signal input
flabel locali s 15864 1939 15898 1973 0 FreeSans 200 180 0 0 B
port 2 nsew signal input
flabel nwell s 16140 1701 16174 1735 0 FreeSans 200 180 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 16140 2245 16174 2279 0 FreeSans 200 180 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 16140 2245 16174 2279 0 FreeSans 200 180 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 16140 1701 16174 1735 0 FreeSans 200 180 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 16204 2262 16204 2262 8 fa_1
rlabel locali s 15680 1990 15758 2056 5 A
port 1 nsew signal input
rlabel locali s 15279 2007 15354 2071 5 A
port 1 nsew signal input
rlabel locali s 14939 2007 15027 2055 5 A
port 1 nsew signal input
rlabel metal1 s 14928 2001 14986 2010 5 A
port 1 nsew signal input
rlabel metal1 s 14928 2038 14986 2047 5 A
port 1 nsew signal input
rlabel metal1 s 15296 2001 15354 2010 5 A
port 1 nsew signal input
rlabel metal1 s 15296 2038 15354 2047 5 A
port 1 nsew signal input
rlabel metal1 s 15668 2001 15726 2010 5 A
port 1 nsew signal input
rlabel metal1 s 15668 2038 15726 2047 5 A
port 1 nsew signal input
rlabel metal1 s 15944 2001 16002 2010 5 A
port 1 nsew signal input
rlabel metal1 s 14928 2010 16002 2038 5 A
port 1 nsew signal input
rlabel metal1 s 15944 2038 16002 2047 5 A
port 1 nsew signal input
rlabel locali s 15492 1909 15564 1975 5 B
port 2 nsew signal input
rlabel locali s 14993 1909 15077 1973 5 B
port 2 nsew signal input
rlabel metal1 s 15020 1933 15078 1942 5 B
port 2 nsew signal input
rlabel metal1 s 15020 1970 15078 1979 5 B
port 2 nsew signal input
rlabel metal1 s 15480 1933 15538 1942 5 B
port 2 nsew signal input
rlabel metal1 s 15480 1970 15538 1979 5 B
port 2 nsew signal input
rlabel metal1 s 15852 1933 15910 1942 5 B
port 2 nsew signal input
rlabel metal1 s 15020 1942 15910 1970 5 B
port 2 nsew signal input
rlabel metal1 s 15852 1970 15910 1979 5 B
port 2 nsew signal input
rlabel metal1 s 14732 2214 16204 2310 5 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 14732 1670 16204 1766 5 VPWR
port 7 nsew power bidirectional abutment
flabel locali s 14270 1807 14304 1841 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 14270 1875 14304 1909 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 14270 2147 14304 2181 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 13254 1875 13288 1909 0 FreeSans 200 180 0 0 CIN
port 3 nsew signal input
flabel locali s 12886 2147 12920 2181 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 12886 2079 12920 2113 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 12886 2011 12920 2045 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 12886 1943 12920 1977 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 12886 1875 12920 1909 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 12886 1807 12920 1841 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 14086 2011 14120 2045 0 FreeSans 200 180 0 0 A
port 1 nsew signal input
flabel locali s 13994 1943 14028 1977 0 FreeSans 200 180 0 0 B
port 2 nsew signal input
flabel nwell s 14270 1705 14304 1739 0 FreeSans 200 180 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 14270 2249 14304 2283 0 FreeSans 200 180 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 14270 2249 14304 2283 0 FreeSans 200 180 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 14270 1705 14304 1739 0 FreeSans 200 180 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 14334 2266 14334 2266 8 fa_1
rlabel locali s 13810 1994 13888 2060 5 A
port 1 nsew signal input
rlabel locali s 13409 2011 13484 2075 5 A
port 1 nsew signal input
rlabel locali s 13069 2011 13157 2059 5 A
port 1 nsew signal input
rlabel metal1 s 13058 2005 13116 2014 5 A
port 1 nsew signal input
rlabel metal1 s 13058 2042 13116 2051 5 A
port 1 nsew signal input
rlabel metal1 s 13426 2005 13484 2014 5 A
port 1 nsew signal input
rlabel metal1 s 13426 2042 13484 2051 5 A
port 1 nsew signal input
rlabel metal1 s 13798 2005 13856 2014 5 A
port 1 nsew signal input
rlabel metal1 s 13798 2042 13856 2051 5 A
port 1 nsew signal input
rlabel metal1 s 14074 2005 14132 2014 5 A
port 1 nsew signal input
rlabel metal1 s 13058 2014 14132 2042 5 A
port 1 nsew signal input
rlabel metal1 s 14074 2042 14132 2051 5 A
port 1 nsew signal input
rlabel locali s 13622 1913 13694 1979 5 B
port 2 nsew signal input
rlabel locali s 13123 1913 13207 1977 5 B
port 2 nsew signal input
rlabel metal1 s 13150 1937 13208 1946 5 B
port 2 nsew signal input
rlabel metal1 s 13150 1974 13208 1983 5 B
port 2 nsew signal input
rlabel metal1 s 13610 1937 13668 1946 5 B
port 2 nsew signal input
rlabel metal1 s 13610 1974 13668 1983 5 B
port 2 nsew signal input
rlabel metal1 s 13982 1937 14040 1946 5 B
port 2 nsew signal input
rlabel metal1 s 13150 1946 14040 1974 5 B
port 2 nsew signal input
rlabel metal1 s 13982 1974 14040 1983 5 B
port 2 nsew signal input
rlabel metal1 s 12862 2218 14334 2314 5 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 12862 1674 14334 1770 5 VPWR
port 7 nsew power bidirectional abutment
flabel locali s 10584 1815 10618 1849 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 10584 1883 10618 1917 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 10584 2155 10618 2189 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 9568 1883 9602 1917 0 FreeSans 200 180 0 0 CIN
port 3 nsew signal input
flabel locali s 9200 2155 9234 2189 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 9200 2087 9234 2121 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 9200 2019 9234 2053 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 9200 1951 9234 1985 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 9200 1883 9234 1917 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 9200 1815 9234 1849 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 10400 2019 10434 2053 0 FreeSans 200 180 0 0 A
port 1 nsew signal input
flabel locali s 10308 1951 10342 1985 0 FreeSans 200 180 0 0 B
port 2 nsew signal input
flabel nwell s 10584 1713 10618 1747 0 FreeSans 200 180 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 10584 2257 10618 2291 0 FreeSans 200 180 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 10584 2257 10618 2291 0 FreeSans 200 180 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 10584 1713 10618 1747 0 FreeSans 200 180 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 10648 2274 10648 2274 8 fa_1
rlabel locali s 10124 2002 10202 2068 5 A
port 1 nsew signal input
rlabel locali s 9723 2019 9798 2083 5 A
port 1 nsew signal input
rlabel locali s 9383 2019 9471 2067 5 A
port 1 nsew signal input
rlabel metal1 s 9372 2013 9430 2022 5 A
port 1 nsew signal input
rlabel metal1 s 9372 2050 9430 2059 5 A
port 1 nsew signal input
rlabel metal1 s 9740 2013 9798 2022 5 A
port 1 nsew signal input
rlabel metal1 s 9740 2050 9798 2059 5 A
port 1 nsew signal input
rlabel metal1 s 10112 2013 10170 2022 5 A
port 1 nsew signal input
rlabel metal1 s 10112 2050 10170 2059 5 A
port 1 nsew signal input
rlabel metal1 s 10388 2013 10446 2022 5 A
port 1 nsew signal input
rlabel metal1 s 9372 2022 10446 2050 5 A
port 1 nsew signal input
rlabel metal1 s 10388 2050 10446 2059 5 A
port 1 nsew signal input
rlabel locali s 9936 1921 10008 1987 5 B
port 2 nsew signal input
rlabel locali s 9437 1921 9521 1985 5 B
port 2 nsew signal input
rlabel metal1 s 9464 1945 9522 1954 5 B
port 2 nsew signal input
rlabel metal1 s 9464 1982 9522 1991 5 B
port 2 nsew signal input
rlabel metal1 s 9924 1945 9982 1954 5 B
port 2 nsew signal input
rlabel metal1 s 9924 1982 9982 1991 5 B
port 2 nsew signal input
rlabel metal1 s 10296 1945 10354 1954 5 B
port 2 nsew signal input
rlabel metal1 s 9464 1954 10354 1982 5 B
port 2 nsew signal input
rlabel metal1 s 10296 1982 10354 1991 5 B
port 2 nsew signal input
rlabel metal1 s 9176 2226 10648 2322 5 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 9176 1682 10648 1778 5 VPWR
port 7 nsew power bidirectional abutment
flabel locali s 12454 1811 12488 1845 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 12454 1879 12488 1913 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 12454 2151 12488 2185 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 11438 1879 11472 1913 0 FreeSans 200 180 0 0 CIN
port 3 nsew signal input
flabel locali s 11070 2151 11104 2185 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 11070 2083 11104 2117 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 11070 2015 11104 2049 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 11070 1947 11104 1981 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 11070 1879 11104 1913 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 11070 1811 11104 1845 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 12270 2015 12304 2049 0 FreeSans 200 180 0 0 A
port 1 nsew signal input
flabel locali s 12178 1947 12212 1981 0 FreeSans 200 180 0 0 B
port 2 nsew signal input
flabel nwell s 12454 1709 12488 1743 0 FreeSans 200 180 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 12454 2253 12488 2287 0 FreeSans 200 180 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 12454 2253 12488 2287 0 FreeSans 200 180 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 12454 1709 12488 1743 0 FreeSans 200 180 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 12518 2270 12518 2270 8 fa_1
rlabel locali s 11994 1998 12072 2064 5 A
port 1 nsew signal input
rlabel locali s 11593 2015 11668 2079 5 A
port 1 nsew signal input
rlabel locali s 11253 2015 11341 2063 5 A
port 1 nsew signal input
rlabel metal1 s 11242 2009 11300 2018 5 A
port 1 nsew signal input
rlabel metal1 s 11242 2046 11300 2055 5 A
port 1 nsew signal input
rlabel metal1 s 11610 2009 11668 2018 5 A
port 1 nsew signal input
rlabel metal1 s 11610 2046 11668 2055 5 A
port 1 nsew signal input
rlabel metal1 s 11982 2009 12040 2018 5 A
port 1 nsew signal input
rlabel metal1 s 11982 2046 12040 2055 5 A
port 1 nsew signal input
rlabel metal1 s 12258 2009 12316 2018 5 A
port 1 nsew signal input
rlabel metal1 s 11242 2018 12316 2046 5 A
port 1 nsew signal input
rlabel metal1 s 12258 2046 12316 2055 5 A
port 1 nsew signal input
rlabel locali s 11806 1917 11878 1983 5 B
port 2 nsew signal input
rlabel locali s 11307 1917 11391 1981 5 B
port 2 nsew signal input
rlabel metal1 s 11334 1941 11392 1950 5 B
port 2 nsew signal input
rlabel metal1 s 11334 1978 11392 1987 5 B
port 2 nsew signal input
rlabel metal1 s 11794 1941 11852 1950 5 B
port 2 nsew signal input
rlabel metal1 s 11794 1978 11852 1987 5 B
port 2 nsew signal input
rlabel metal1 s 12166 1941 12224 1950 5 B
port 2 nsew signal input
rlabel metal1 s 11334 1950 12224 1978 5 B
port 2 nsew signal input
rlabel metal1 s 12166 1978 12224 1987 5 B
port 2 nsew signal input
rlabel metal1 s 11046 2222 12518 2318 5 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 11046 1678 12518 1774 5 VPWR
port 7 nsew power bidirectional abutment
flabel locali s 6190 6277 6224 6311 0 FreeSans 340 180 0 0 Y
port 6 nsew signal output
flabel locali s 6190 6345 6224 6379 0 FreeSans 340 180 0 0 Y
port 6 nsew signal output
flabel locali s 6282 6345 6316 6379 0 FreeSans 340 180 0 0 A
port 1 nsew signal input
flabel nwell s 6325 6039 6359 6073 0 FreeSans 200 180 0 0 VPB
port 4 nsew power bidirectional
flabel pwell s 6325 6583 6359 6617 0 FreeSans 200 180 0 0 VNB
port 3 nsew ground bidirectional
flabel metal1 s 6325 6583 6359 6617 0 FreeSans 200 180 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel metal1 s 6325 6039 6359 6073 0 FreeSans 200 180 0 0 VPWR
port 5 nsew power bidirectional abutment
rlabel comment s 6388 6600 6388 6600 8 inv_1
rlabel metal1 s 6112 6552 6388 6648 5 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 6112 6008 6388 6104 5 VPWR
port 5 nsew power bidirectional abutment
flabel locali s 8800 5077 8834 5111 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 8800 5145 8834 5179 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 8800 5417 8834 5451 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 7784 5145 7818 5179 0 FreeSans 200 180 0 0 CIN
port 3 nsew signal input
flabel locali s 7416 5417 7450 5451 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 7416 5349 7450 5383 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 7416 5281 7450 5315 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 7416 5213 7450 5247 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 7416 5145 7450 5179 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 7416 5077 7450 5111 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 8616 5281 8650 5315 0 FreeSans 200 180 0 0 A
port 1 nsew signal input
flabel locali s 8524 5213 8558 5247 0 FreeSans 200 180 0 0 B
port 2 nsew signal input
flabel nwell s 8800 4975 8834 5009 0 FreeSans 200 180 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 8800 5519 8834 5553 0 FreeSans 200 180 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 8800 5519 8834 5553 0 FreeSans 200 180 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 8800 4975 8834 5009 0 FreeSans 200 180 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 8864 5536 8864 5536 8 fa_1
rlabel locali s 8340 5264 8418 5330 5 A
port 1 nsew signal input
rlabel locali s 7939 5281 8014 5345 5 A
port 1 nsew signal input
rlabel locali s 7599 5281 7687 5329 5 A
port 1 nsew signal input
rlabel metal1 s 7588 5275 7646 5284 5 A
port 1 nsew signal input
rlabel metal1 s 7588 5312 7646 5321 5 A
port 1 nsew signal input
rlabel metal1 s 7956 5275 8014 5284 5 A
port 1 nsew signal input
rlabel metal1 s 7956 5312 8014 5321 5 A
port 1 nsew signal input
rlabel metal1 s 8328 5275 8386 5284 5 A
port 1 nsew signal input
rlabel metal1 s 8328 5312 8386 5321 5 A
port 1 nsew signal input
rlabel metal1 s 8604 5275 8662 5284 5 A
port 1 nsew signal input
rlabel metal1 s 7588 5284 8662 5312 5 A
port 1 nsew signal input
rlabel metal1 s 8604 5312 8662 5321 5 A
port 1 nsew signal input
rlabel locali s 8152 5183 8224 5249 5 B
port 2 nsew signal input
rlabel locali s 7653 5183 7737 5247 5 B
port 2 nsew signal input
rlabel metal1 s 7680 5207 7738 5216 5 B
port 2 nsew signal input
rlabel metal1 s 7680 5244 7738 5253 5 B
port 2 nsew signal input
rlabel metal1 s 8140 5207 8198 5216 5 B
port 2 nsew signal input
rlabel metal1 s 8140 5244 8198 5253 5 B
port 2 nsew signal input
rlabel metal1 s 8512 5207 8570 5216 5 B
port 2 nsew signal input
rlabel metal1 s 7680 5216 8570 5244 5 B
port 2 nsew signal input
rlabel metal1 s 8512 5244 8570 5253 5 B
port 2 nsew signal input
rlabel metal1 s 7392 5488 8864 5584 5 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 7392 4944 8864 5040 5 VPWR
port 7 nsew power bidirectional abutment
flabel locali s 6930 5081 6964 5115 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 6930 5149 6964 5183 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 6930 5421 6964 5455 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 5914 5149 5948 5183 0 FreeSans 200 180 0 0 CIN
port 3 nsew signal input
flabel locali s 5546 5421 5580 5455 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 5546 5353 5580 5387 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 5546 5285 5580 5319 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 5546 5217 5580 5251 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 5546 5149 5580 5183 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 5546 5081 5580 5115 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 6746 5285 6780 5319 0 FreeSans 200 180 0 0 A
port 1 nsew signal input
flabel locali s 6654 5217 6688 5251 0 FreeSans 200 180 0 0 B
port 2 nsew signal input
flabel nwell s 6930 4979 6964 5013 0 FreeSans 200 180 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 6930 5523 6964 5557 0 FreeSans 200 180 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 6930 5523 6964 5557 0 FreeSans 200 180 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 6930 4979 6964 5013 0 FreeSans 200 180 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 6994 5540 6994 5540 8 fa_1
rlabel locali s 6470 5268 6548 5334 5 A
port 1 nsew signal input
rlabel locali s 6069 5285 6144 5349 5 A
port 1 nsew signal input
rlabel locali s 5729 5285 5817 5333 5 A
port 1 nsew signal input
rlabel metal1 s 5718 5279 5776 5288 5 A
port 1 nsew signal input
rlabel metal1 s 5718 5316 5776 5325 5 A
port 1 nsew signal input
rlabel metal1 s 6086 5279 6144 5288 5 A
port 1 nsew signal input
rlabel metal1 s 6086 5316 6144 5325 5 A
port 1 nsew signal input
rlabel metal1 s 6458 5279 6516 5288 5 A
port 1 nsew signal input
rlabel metal1 s 6458 5316 6516 5325 5 A
port 1 nsew signal input
rlabel metal1 s 6734 5279 6792 5288 5 A
port 1 nsew signal input
rlabel metal1 s 5718 5288 6792 5316 5 A
port 1 nsew signal input
rlabel metal1 s 6734 5316 6792 5325 5 A
port 1 nsew signal input
rlabel locali s 6282 5187 6354 5253 5 B
port 2 nsew signal input
rlabel locali s 5783 5187 5867 5251 5 B
port 2 nsew signal input
rlabel metal1 s 5810 5211 5868 5220 5 B
port 2 nsew signal input
rlabel metal1 s 5810 5248 5868 5257 5 B
port 2 nsew signal input
rlabel metal1 s 6270 5211 6328 5220 5 B
port 2 nsew signal input
rlabel metal1 s 6270 5248 6328 5257 5 B
port 2 nsew signal input
rlabel metal1 s 6642 5211 6700 5220 5 B
port 2 nsew signal input
rlabel metal1 s 5810 5220 6700 5248 5 B
port 2 nsew signal input
rlabel metal1 s 6642 5248 6700 5257 5 B
port 2 nsew signal input
rlabel metal1 s 5522 5492 6994 5588 5 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 5522 4948 6994 5044 5 VPWR
port 7 nsew power bidirectional abutment
flabel locali s 3244 5089 3278 5123 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 3244 5157 3278 5191 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 3244 5429 3278 5463 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 2228 5157 2262 5191 0 FreeSans 200 180 0 0 CIN
port 3 nsew signal input
flabel locali s 1860 5429 1894 5463 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 1860 5361 1894 5395 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 1860 5293 1894 5327 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 1860 5225 1894 5259 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 1860 5157 1894 5191 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 1860 5089 1894 5123 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 3060 5293 3094 5327 0 FreeSans 200 180 0 0 A
port 1 nsew signal input
flabel locali s 2968 5225 3002 5259 0 FreeSans 200 180 0 0 B
port 2 nsew signal input
flabel nwell s 3244 4987 3278 5021 0 FreeSans 200 180 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 3244 5531 3278 5565 0 FreeSans 200 180 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 3244 5531 3278 5565 0 FreeSans 200 180 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 3244 4987 3278 5021 0 FreeSans 200 180 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 3308 5548 3308 5548 8 fa_1
rlabel locali s 2784 5276 2862 5342 5 A
port 1 nsew signal input
rlabel locali s 2383 5293 2458 5357 5 A
port 1 nsew signal input
rlabel locali s 2043 5293 2131 5341 5 A
port 1 nsew signal input
rlabel metal1 s 2032 5287 2090 5296 5 A
port 1 nsew signal input
rlabel metal1 s 2032 5324 2090 5333 5 A
port 1 nsew signal input
rlabel metal1 s 2400 5287 2458 5296 5 A
port 1 nsew signal input
rlabel metal1 s 2400 5324 2458 5333 5 A
port 1 nsew signal input
rlabel metal1 s 2772 5287 2830 5296 5 A
port 1 nsew signal input
rlabel metal1 s 2772 5324 2830 5333 5 A
port 1 nsew signal input
rlabel metal1 s 3048 5287 3106 5296 5 A
port 1 nsew signal input
rlabel metal1 s 2032 5296 3106 5324 5 A
port 1 nsew signal input
rlabel metal1 s 3048 5324 3106 5333 5 A
port 1 nsew signal input
rlabel locali s 2596 5195 2668 5261 5 B
port 2 nsew signal input
rlabel locali s 2097 5195 2181 5259 5 B
port 2 nsew signal input
rlabel metal1 s 2124 5219 2182 5228 5 B
port 2 nsew signal input
rlabel metal1 s 2124 5256 2182 5265 5 B
port 2 nsew signal input
rlabel metal1 s 2584 5219 2642 5228 5 B
port 2 nsew signal input
rlabel metal1 s 2584 5256 2642 5265 5 B
port 2 nsew signal input
rlabel metal1 s 2956 5219 3014 5228 5 B
port 2 nsew signal input
rlabel metal1 s 2124 5228 3014 5256 5 B
port 2 nsew signal input
rlabel metal1 s 2956 5256 3014 5265 5 B
port 2 nsew signal input
rlabel metal1 s 1836 5500 3308 5596 5 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1836 4956 3308 5052 5 VPWR
port 7 nsew power bidirectional abutment
flabel locali s 5114 5085 5148 5119 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 5114 5153 5148 5187 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 5114 5425 5148 5459 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 4098 5153 4132 5187 0 FreeSans 200 180 0 0 CIN
port 3 nsew signal input
flabel locali s 3730 5425 3764 5459 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 3730 5357 3764 5391 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 3730 5289 3764 5323 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 3730 5221 3764 5255 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 3730 5153 3764 5187 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 3730 5085 3764 5119 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 4930 5289 4964 5323 0 FreeSans 200 180 0 0 A
port 1 nsew signal input
flabel locali s 4838 5221 4872 5255 0 FreeSans 200 180 0 0 B
port 2 nsew signal input
flabel nwell s 5114 4983 5148 5017 0 FreeSans 200 180 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 5114 5527 5148 5561 0 FreeSans 200 180 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 5114 5527 5148 5561 0 FreeSans 200 180 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 5114 4983 5148 5017 0 FreeSans 200 180 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 5178 5544 5178 5544 8 fa_1
rlabel locali s 4654 5272 4732 5338 5 A
port 1 nsew signal input
rlabel locali s 4253 5289 4328 5353 5 A
port 1 nsew signal input
rlabel locali s 3913 5289 4001 5337 5 A
port 1 nsew signal input
rlabel metal1 s 3902 5283 3960 5292 5 A
port 1 nsew signal input
rlabel metal1 s 3902 5320 3960 5329 5 A
port 1 nsew signal input
rlabel metal1 s 4270 5283 4328 5292 5 A
port 1 nsew signal input
rlabel metal1 s 4270 5320 4328 5329 5 A
port 1 nsew signal input
rlabel metal1 s 4642 5283 4700 5292 5 A
port 1 nsew signal input
rlabel metal1 s 4642 5320 4700 5329 5 A
port 1 nsew signal input
rlabel metal1 s 4918 5283 4976 5292 5 A
port 1 nsew signal input
rlabel metal1 s 3902 5292 4976 5320 5 A
port 1 nsew signal input
rlabel metal1 s 4918 5320 4976 5329 5 A
port 1 nsew signal input
rlabel locali s 4466 5191 4538 5257 5 B
port 2 nsew signal input
rlabel locali s 3967 5191 4051 5255 5 B
port 2 nsew signal input
rlabel metal1 s 3994 5215 4052 5224 5 B
port 2 nsew signal input
rlabel metal1 s 3994 5252 4052 5261 5 B
port 2 nsew signal input
rlabel metal1 s 4454 5215 4512 5224 5 B
port 2 nsew signal input
rlabel metal1 s 4454 5252 4512 5261 5 B
port 2 nsew signal input
rlabel metal1 s 4826 5215 4884 5224 5 B
port 2 nsew signal input
rlabel metal1 s 3994 5224 4884 5252 5 B
port 2 nsew signal input
rlabel metal1 s 4826 5252 4884 5261 5 B
port 2 nsew signal input
rlabel metal1 s 3706 5496 5178 5592 5 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3706 4952 5178 5048 5 VPWR
port 7 nsew power bidirectional abutment
flabel locali s 14340 4627 14374 4661 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 14340 4695 14374 4729 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 14340 4967 14374 5001 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 13324 4695 13358 4729 0 FreeSans 200 180 0 0 CIN
port 3 nsew signal input
flabel locali s 12956 4967 12990 5001 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 12956 4899 12990 4933 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 12956 4831 12990 4865 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 12956 4763 12990 4797 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 12956 4695 12990 4729 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 12956 4627 12990 4661 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 14156 4831 14190 4865 0 FreeSans 200 180 0 0 A
port 1 nsew signal input
flabel locali s 14064 4763 14098 4797 0 FreeSans 200 180 0 0 B
port 2 nsew signal input
flabel nwell s 14340 4525 14374 4559 0 FreeSans 200 180 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 14340 5069 14374 5103 0 FreeSans 200 180 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 14340 5069 14374 5103 0 FreeSans 200 180 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 14340 4525 14374 4559 0 FreeSans 200 180 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 14404 5086 14404 5086 8 fa_1
rlabel locali s 13880 4814 13958 4880 5 A
port 1 nsew signal input
rlabel locali s 13479 4831 13554 4895 5 A
port 1 nsew signal input
rlabel locali s 13139 4831 13227 4879 5 A
port 1 nsew signal input
rlabel metal1 s 13128 4825 13186 4834 5 A
port 1 nsew signal input
rlabel metal1 s 13128 4862 13186 4871 5 A
port 1 nsew signal input
rlabel metal1 s 13496 4825 13554 4834 5 A
port 1 nsew signal input
rlabel metal1 s 13496 4862 13554 4871 5 A
port 1 nsew signal input
rlabel metal1 s 13868 4825 13926 4834 5 A
port 1 nsew signal input
rlabel metal1 s 13868 4862 13926 4871 5 A
port 1 nsew signal input
rlabel metal1 s 14144 4825 14202 4834 5 A
port 1 nsew signal input
rlabel metal1 s 13128 4834 14202 4862 5 A
port 1 nsew signal input
rlabel metal1 s 14144 4862 14202 4871 5 A
port 1 nsew signal input
rlabel locali s 13692 4733 13764 4799 5 B
port 2 nsew signal input
rlabel locali s 13193 4733 13277 4797 5 B
port 2 nsew signal input
rlabel metal1 s 13220 4757 13278 4766 5 B
port 2 nsew signal input
rlabel metal1 s 13220 4794 13278 4803 5 B
port 2 nsew signal input
rlabel metal1 s 13680 4757 13738 4766 5 B
port 2 nsew signal input
rlabel metal1 s 13680 4794 13738 4803 5 B
port 2 nsew signal input
rlabel metal1 s 14052 4757 14110 4766 5 B
port 2 nsew signal input
rlabel metal1 s 13220 4766 14110 4794 5 B
port 2 nsew signal input
rlabel metal1 s 14052 4794 14110 4803 5 B
port 2 nsew signal input
rlabel metal1 s 12932 5038 14404 5134 5 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 12932 4494 14404 4590 5 VPWR
port 7 nsew power bidirectional abutment
flabel locali s 10654 4635 10688 4669 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 10654 4703 10688 4737 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 10654 4975 10688 5009 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 9638 4703 9672 4737 0 FreeSans 200 180 0 0 CIN
port 3 nsew signal input
flabel locali s 9270 4975 9304 5009 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 9270 4907 9304 4941 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 9270 4839 9304 4873 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 9270 4771 9304 4805 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 9270 4703 9304 4737 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 9270 4635 9304 4669 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 10470 4839 10504 4873 0 FreeSans 200 180 0 0 A
port 1 nsew signal input
flabel locali s 10378 4771 10412 4805 0 FreeSans 200 180 0 0 B
port 2 nsew signal input
flabel nwell s 10654 4533 10688 4567 0 FreeSans 200 180 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 10654 5077 10688 5111 0 FreeSans 200 180 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 10654 5077 10688 5111 0 FreeSans 200 180 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 10654 4533 10688 4567 0 FreeSans 200 180 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 10718 5094 10718 5094 8 fa_1
rlabel locali s 10194 4822 10272 4888 5 A
port 1 nsew signal input
rlabel locali s 9793 4839 9868 4903 5 A
port 1 nsew signal input
rlabel locali s 9453 4839 9541 4887 5 A
port 1 nsew signal input
rlabel metal1 s 9442 4833 9500 4842 5 A
port 1 nsew signal input
rlabel metal1 s 9442 4870 9500 4879 5 A
port 1 nsew signal input
rlabel metal1 s 9810 4833 9868 4842 5 A
port 1 nsew signal input
rlabel metal1 s 9810 4870 9868 4879 5 A
port 1 nsew signal input
rlabel metal1 s 10182 4833 10240 4842 5 A
port 1 nsew signal input
rlabel metal1 s 10182 4870 10240 4879 5 A
port 1 nsew signal input
rlabel metal1 s 10458 4833 10516 4842 5 A
port 1 nsew signal input
rlabel metal1 s 9442 4842 10516 4870 5 A
port 1 nsew signal input
rlabel metal1 s 10458 4870 10516 4879 5 A
port 1 nsew signal input
rlabel locali s 10006 4741 10078 4807 5 B
port 2 nsew signal input
rlabel locali s 9507 4741 9591 4805 5 B
port 2 nsew signal input
rlabel metal1 s 9534 4765 9592 4774 5 B
port 2 nsew signal input
rlabel metal1 s 9534 4802 9592 4811 5 B
port 2 nsew signal input
rlabel metal1 s 9994 4765 10052 4774 5 B
port 2 nsew signal input
rlabel metal1 s 9994 4802 10052 4811 5 B
port 2 nsew signal input
rlabel metal1 s 10366 4765 10424 4774 5 B
port 2 nsew signal input
rlabel metal1 s 9534 4774 10424 4802 5 B
port 2 nsew signal input
rlabel metal1 s 10366 4802 10424 4811 5 B
port 2 nsew signal input
rlabel metal1 s 9246 5046 10718 5142 5 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 9246 4502 10718 4598 5 VPWR
port 7 nsew power bidirectional abutment
flabel locali s 12524 4631 12558 4665 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 12524 4699 12558 4733 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 12524 4971 12558 5005 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 11508 4699 11542 4733 0 FreeSans 200 180 0 0 CIN
port 3 nsew signal input
flabel locali s 11140 4971 11174 5005 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 11140 4903 11174 4937 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 11140 4835 11174 4869 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 11140 4767 11174 4801 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 11140 4699 11174 4733 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 11140 4631 11174 4665 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 12340 4835 12374 4869 0 FreeSans 200 180 0 0 A
port 1 nsew signal input
flabel locali s 12248 4767 12282 4801 0 FreeSans 200 180 0 0 B
port 2 nsew signal input
flabel nwell s 12524 4529 12558 4563 0 FreeSans 200 180 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 12524 5073 12558 5107 0 FreeSans 200 180 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 12524 5073 12558 5107 0 FreeSans 200 180 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 12524 4529 12558 4563 0 FreeSans 200 180 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 12588 5090 12588 5090 8 fa_1
rlabel locali s 12064 4818 12142 4884 5 A
port 1 nsew signal input
rlabel locali s 11663 4835 11738 4899 5 A
port 1 nsew signal input
rlabel locali s 11323 4835 11411 4883 5 A
port 1 nsew signal input
rlabel metal1 s 11312 4829 11370 4838 5 A
port 1 nsew signal input
rlabel metal1 s 11312 4866 11370 4875 5 A
port 1 nsew signal input
rlabel metal1 s 11680 4829 11738 4838 5 A
port 1 nsew signal input
rlabel metal1 s 11680 4866 11738 4875 5 A
port 1 nsew signal input
rlabel metal1 s 12052 4829 12110 4838 5 A
port 1 nsew signal input
rlabel metal1 s 12052 4866 12110 4875 5 A
port 1 nsew signal input
rlabel metal1 s 12328 4829 12386 4838 5 A
port 1 nsew signal input
rlabel metal1 s 11312 4838 12386 4866 5 A
port 1 nsew signal input
rlabel metal1 s 12328 4866 12386 4875 5 A
port 1 nsew signal input
rlabel locali s 11876 4737 11948 4803 5 B
port 2 nsew signal input
rlabel locali s 11377 4737 11461 4801 5 B
port 2 nsew signal input
rlabel metal1 s 11404 4761 11462 4770 5 B
port 2 nsew signal input
rlabel metal1 s 11404 4798 11462 4807 5 B
port 2 nsew signal input
rlabel metal1 s 11864 4761 11922 4770 5 B
port 2 nsew signal input
rlabel metal1 s 11864 4798 11922 4807 5 B
port 2 nsew signal input
rlabel metal1 s 12236 4761 12294 4770 5 B
port 2 nsew signal input
rlabel metal1 s 11404 4770 12294 4798 5 B
port 2 nsew signal input
rlabel metal1 s 12236 4798 12294 4807 5 B
port 2 nsew signal input
rlabel metal1 s 11116 5042 12588 5138 5 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 11116 4498 12588 4594 5 VPWR
port 7 nsew power bidirectional abutment
flabel locali s 14312 5501 14346 5535 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 14312 5569 14346 5603 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 14312 5841 14346 5875 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 13296 5569 13330 5603 0 FreeSans 200 180 0 0 CIN
port 3 nsew signal input
flabel locali s 12928 5841 12962 5875 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 12928 5773 12962 5807 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 12928 5705 12962 5739 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 12928 5637 12962 5671 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 12928 5569 12962 5603 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 12928 5501 12962 5535 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 14128 5705 14162 5739 0 FreeSans 200 180 0 0 A
port 1 nsew signal input
flabel locali s 14036 5637 14070 5671 0 FreeSans 200 180 0 0 B
port 2 nsew signal input
flabel nwell s 14312 5399 14346 5433 0 FreeSans 200 180 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 14312 5943 14346 5977 0 FreeSans 200 180 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 14312 5943 14346 5977 0 FreeSans 200 180 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 14312 5399 14346 5433 0 FreeSans 200 180 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 14376 5960 14376 5960 8 fa_1
rlabel locali s 13852 5688 13930 5754 5 A
port 1 nsew signal input
rlabel locali s 13451 5705 13526 5769 5 A
port 1 nsew signal input
rlabel locali s 13111 5705 13199 5753 5 A
port 1 nsew signal input
rlabel metal1 s 13100 5699 13158 5708 5 A
port 1 nsew signal input
rlabel metal1 s 13100 5736 13158 5745 5 A
port 1 nsew signal input
rlabel metal1 s 13468 5699 13526 5708 5 A
port 1 nsew signal input
rlabel metal1 s 13468 5736 13526 5745 5 A
port 1 nsew signal input
rlabel metal1 s 13840 5699 13898 5708 5 A
port 1 nsew signal input
rlabel metal1 s 13840 5736 13898 5745 5 A
port 1 nsew signal input
rlabel metal1 s 14116 5699 14174 5708 5 A
port 1 nsew signal input
rlabel metal1 s 13100 5708 14174 5736 5 A
port 1 nsew signal input
rlabel metal1 s 14116 5736 14174 5745 5 A
port 1 nsew signal input
rlabel locali s 13664 5607 13736 5673 5 B
port 2 nsew signal input
rlabel locali s 13165 5607 13249 5671 5 B
port 2 nsew signal input
rlabel metal1 s 13192 5631 13250 5640 5 B
port 2 nsew signal input
rlabel metal1 s 13192 5668 13250 5677 5 B
port 2 nsew signal input
rlabel metal1 s 13652 5631 13710 5640 5 B
port 2 nsew signal input
rlabel metal1 s 13652 5668 13710 5677 5 B
port 2 nsew signal input
rlabel metal1 s 14024 5631 14082 5640 5 B
port 2 nsew signal input
rlabel metal1 s 13192 5640 14082 5668 5 B
port 2 nsew signal input
rlabel metal1 s 14024 5668 14082 5677 5 B
port 2 nsew signal input
rlabel metal1 s 12904 5912 14376 6008 5 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 12904 5368 14376 5464 5 VPWR
port 7 nsew power bidirectional abutment
flabel locali s 10626 5509 10660 5543 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 10626 5577 10660 5611 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 10626 5849 10660 5883 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 9610 5577 9644 5611 0 FreeSans 200 180 0 0 CIN
port 3 nsew signal input
flabel locali s 9242 5849 9276 5883 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 9242 5781 9276 5815 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 9242 5713 9276 5747 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 9242 5645 9276 5679 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 9242 5577 9276 5611 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 9242 5509 9276 5543 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 10442 5713 10476 5747 0 FreeSans 200 180 0 0 A
port 1 nsew signal input
flabel locali s 10350 5645 10384 5679 0 FreeSans 200 180 0 0 B
port 2 nsew signal input
flabel nwell s 10626 5407 10660 5441 0 FreeSans 200 180 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 10626 5951 10660 5985 0 FreeSans 200 180 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 10626 5951 10660 5985 0 FreeSans 200 180 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 10626 5407 10660 5441 0 FreeSans 200 180 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 10690 5968 10690 5968 8 fa_1
rlabel locali s 10166 5696 10244 5762 5 A
port 1 nsew signal input
rlabel locali s 9765 5713 9840 5777 5 A
port 1 nsew signal input
rlabel locali s 9425 5713 9513 5761 5 A
port 1 nsew signal input
rlabel metal1 s 9414 5707 9472 5716 5 A
port 1 nsew signal input
rlabel metal1 s 9414 5744 9472 5753 5 A
port 1 nsew signal input
rlabel metal1 s 9782 5707 9840 5716 5 A
port 1 nsew signal input
rlabel metal1 s 9782 5744 9840 5753 5 A
port 1 nsew signal input
rlabel metal1 s 10154 5707 10212 5716 5 A
port 1 nsew signal input
rlabel metal1 s 10154 5744 10212 5753 5 A
port 1 nsew signal input
rlabel metal1 s 10430 5707 10488 5716 5 A
port 1 nsew signal input
rlabel metal1 s 9414 5716 10488 5744 5 A
port 1 nsew signal input
rlabel metal1 s 10430 5744 10488 5753 5 A
port 1 nsew signal input
rlabel locali s 9978 5615 10050 5681 5 B
port 2 nsew signal input
rlabel locali s 9479 5615 9563 5679 5 B
port 2 nsew signal input
rlabel metal1 s 9506 5639 9564 5648 5 B
port 2 nsew signal input
rlabel metal1 s 9506 5676 9564 5685 5 B
port 2 nsew signal input
rlabel metal1 s 9966 5639 10024 5648 5 B
port 2 nsew signal input
rlabel metal1 s 9966 5676 10024 5685 5 B
port 2 nsew signal input
rlabel metal1 s 10338 5639 10396 5648 5 B
port 2 nsew signal input
rlabel metal1 s 9506 5648 10396 5676 5 B
port 2 nsew signal input
rlabel metal1 s 10338 5676 10396 5685 5 B
port 2 nsew signal input
rlabel metal1 s 9218 5920 10690 6016 5 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 9218 5376 10690 5472 5 VPWR
port 7 nsew power bidirectional abutment
flabel locali s 12496 5505 12530 5539 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 12496 5573 12530 5607 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 12496 5845 12530 5879 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 11480 5573 11514 5607 0 FreeSans 200 180 0 0 CIN
port 3 nsew signal input
flabel locali s 11112 5845 11146 5879 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 11112 5777 11146 5811 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 11112 5709 11146 5743 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 11112 5641 11146 5675 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 11112 5573 11146 5607 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 11112 5505 11146 5539 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 12312 5709 12346 5743 0 FreeSans 200 180 0 0 A
port 1 nsew signal input
flabel locali s 12220 5641 12254 5675 0 FreeSans 200 180 0 0 B
port 2 nsew signal input
flabel nwell s 12496 5403 12530 5437 0 FreeSans 200 180 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 12496 5947 12530 5981 0 FreeSans 200 180 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 12496 5947 12530 5981 0 FreeSans 200 180 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 12496 5403 12530 5437 0 FreeSans 200 180 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 12560 5964 12560 5964 8 fa_1
rlabel locali s 12036 5692 12114 5758 5 A
port 1 nsew signal input
rlabel locali s 11635 5709 11710 5773 5 A
port 1 nsew signal input
rlabel locali s 11295 5709 11383 5757 5 A
port 1 nsew signal input
rlabel metal1 s 11284 5703 11342 5712 5 A
port 1 nsew signal input
rlabel metal1 s 11284 5740 11342 5749 5 A
port 1 nsew signal input
rlabel metal1 s 11652 5703 11710 5712 5 A
port 1 nsew signal input
rlabel metal1 s 11652 5740 11710 5749 5 A
port 1 nsew signal input
rlabel metal1 s 12024 5703 12082 5712 5 A
port 1 nsew signal input
rlabel metal1 s 12024 5740 12082 5749 5 A
port 1 nsew signal input
rlabel metal1 s 12300 5703 12358 5712 5 A
port 1 nsew signal input
rlabel metal1 s 11284 5712 12358 5740 5 A
port 1 nsew signal input
rlabel metal1 s 12300 5740 12358 5749 5 A
port 1 nsew signal input
rlabel locali s 11848 5611 11920 5677 5 B
port 2 nsew signal input
rlabel locali s 11349 5611 11433 5675 5 B
port 2 nsew signal input
rlabel metal1 s 11376 5635 11434 5644 5 B
port 2 nsew signal input
rlabel metal1 s 11376 5672 11434 5681 5 B
port 2 nsew signal input
rlabel metal1 s 11836 5635 11894 5644 5 B
port 2 nsew signal input
rlabel metal1 s 11836 5672 11894 5681 5 B
port 2 nsew signal input
rlabel metal1 s 12208 5635 12266 5644 5 B
port 2 nsew signal input
rlabel metal1 s 11376 5644 12266 5672 5 B
port 2 nsew signal input
rlabel metal1 s 12208 5672 12266 5681 5 B
port 2 nsew signal input
rlabel metal1 s 11088 5916 12560 6012 5 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 11088 5372 12560 5468 5 VPWR
port 7 nsew power bidirectional abutment
flabel locali s 16210 4623 16244 4657 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 16210 4691 16244 4725 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 16210 4963 16244 4997 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 15194 4691 15228 4725 0 FreeSans 200 180 0 0 CIN
port 3 nsew signal input
flabel locali s 14826 4963 14860 4997 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 14826 4895 14860 4929 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 14826 4827 14860 4861 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 14826 4759 14860 4793 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 14826 4691 14860 4725 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 14826 4623 14860 4657 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 16026 4827 16060 4861 0 FreeSans 200 180 0 0 A
port 1 nsew signal input
flabel locali s 15934 4759 15968 4793 0 FreeSans 200 180 0 0 B
port 2 nsew signal input
flabel nwell s 16210 4521 16244 4555 0 FreeSans 200 180 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 16210 5065 16244 5099 0 FreeSans 200 180 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 16210 5065 16244 5099 0 FreeSans 200 180 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 16210 4521 16244 4555 0 FreeSans 200 180 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 16274 5082 16274 5082 8 fa_1
rlabel locali s 15750 4810 15828 4876 5 A
port 1 nsew signal input
rlabel locali s 15349 4827 15424 4891 5 A
port 1 nsew signal input
rlabel locali s 15009 4827 15097 4875 5 A
port 1 nsew signal input
rlabel metal1 s 14998 4821 15056 4830 5 A
port 1 nsew signal input
rlabel metal1 s 14998 4858 15056 4867 5 A
port 1 nsew signal input
rlabel metal1 s 15366 4821 15424 4830 5 A
port 1 nsew signal input
rlabel metal1 s 15366 4858 15424 4867 5 A
port 1 nsew signal input
rlabel metal1 s 15738 4821 15796 4830 5 A
port 1 nsew signal input
rlabel metal1 s 15738 4858 15796 4867 5 A
port 1 nsew signal input
rlabel metal1 s 16014 4821 16072 4830 5 A
port 1 nsew signal input
rlabel metal1 s 14998 4830 16072 4858 5 A
port 1 nsew signal input
rlabel metal1 s 16014 4858 16072 4867 5 A
port 1 nsew signal input
rlabel locali s 15562 4729 15634 4795 5 B
port 2 nsew signal input
rlabel locali s 15063 4729 15147 4793 5 B
port 2 nsew signal input
rlabel metal1 s 15090 4753 15148 4762 5 B
port 2 nsew signal input
rlabel metal1 s 15090 4790 15148 4799 5 B
port 2 nsew signal input
rlabel metal1 s 15550 4753 15608 4762 5 B
port 2 nsew signal input
rlabel metal1 s 15550 4790 15608 4799 5 B
port 2 nsew signal input
rlabel metal1 s 15922 4753 15980 4762 5 B
port 2 nsew signal input
rlabel metal1 s 15090 4762 15980 4790 5 B
port 2 nsew signal input
rlabel metal1 s 15922 4790 15980 4799 5 B
port 2 nsew signal input
rlabel metal1 s 14802 5034 16274 5130 5 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 14802 4490 16274 4586 5 VPWR
port 7 nsew power bidirectional abutment
flabel locali s 16182 5497 16216 5531 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 16182 5565 16216 5599 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 16182 5837 16216 5871 0 FreeSans 200 180 0 0 COUT
port 8 nsew signal output
flabel locali s 15166 5565 15200 5599 0 FreeSans 200 180 0 0 CIN
port 3 nsew signal input
flabel locali s 14798 5837 14832 5871 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 14798 5769 14832 5803 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 14798 5701 14832 5735 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 14798 5633 14832 5667 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 14798 5565 14832 5599 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 14798 5497 14832 5531 0 FreeSans 200 180 0 0 SUM
port 9 nsew signal output
flabel locali s 15998 5701 16032 5735 0 FreeSans 200 180 0 0 A
port 1 nsew signal input
flabel locali s 15906 5633 15940 5667 0 FreeSans 200 180 0 0 B
port 2 nsew signal input
flabel nwell s 16182 5395 16216 5429 0 FreeSans 200 180 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 16182 5939 16216 5973 0 FreeSans 200 180 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 16182 5939 16216 5973 0 FreeSans 200 180 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 16182 5395 16216 5429 0 FreeSans 200 180 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 16246 5956 16246 5956 8 fa_1
rlabel locali s 15722 5684 15800 5750 5 A
port 1 nsew signal input
rlabel locali s 15321 5701 15396 5765 5 A
port 1 nsew signal input
rlabel locali s 14981 5701 15069 5749 5 A
port 1 nsew signal input
rlabel metal1 s 14970 5695 15028 5704 5 A
port 1 nsew signal input
rlabel metal1 s 14970 5732 15028 5741 5 A
port 1 nsew signal input
rlabel metal1 s 15338 5695 15396 5704 5 A
port 1 nsew signal input
rlabel metal1 s 15338 5732 15396 5741 5 A
port 1 nsew signal input
rlabel metal1 s 15710 5695 15768 5704 5 A
port 1 nsew signal input
rlabel metal1 s 15710 5732 15768 5741 5 A
port 1 nsew signal input
rlabel metal1 s 15986 5695 16044 5704 5 A
port 1 nsew signal input
rlabel metal1 s 14970 5704 16044 5732 5 A
port 1 nsew signal input
rlabel metal1 s 15986 5732 16044 5741 5 A
port 1 nsew signal input
rlabel locali s 15534 5603 15606 5669 5 B
port 2 nsew signal input
rlabel locali s 15035 5603 15119 5667 5 B
port 2 nsew signal input
rlabel metal1 s 15062 5627 15120 5636 5 B
port 2 nsew signal input
rlabel metal1 s 15062 5664 15120 5673 5 B
port 2 nsew signal input
rlabel metal1 s 15522 5627 15580 5636 5 B
port 2 nsew signal input
rlabel metal1 s 15522 5664 15580 5673 5 B
port 2 nsew signal input
rlabel metal1 s 15894 5627 15952 5636 5 B
port 2 nsew signal input
rlabel metal1 s 15062 5636 15952 5664 5 B
port 2 nsew signal input
rlabel metal1 s 15894 5664 15952 5673 5 B
port 2 nsew signal input
rlabel metal1 s 14774 5908 16246 6004 5 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 14774 5364 16246 5460 5 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 9569 11013 9603 11047 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 9569 10469 9603 10503 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel locali s 9937 10639 9971 10673 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 9937 10571 9971 10605 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 9937 10707 9971 10741 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 9937 10775 9971 10809 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 9937 10843 9971 10877 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 9937 10911 9971 10945 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 9753 10707 9787 10741 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 9661 10707 9695 10741 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 9569 10707 9603 10741 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel nwell s 9569 11013 9603 11047 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 9569 10469 9603 10503 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
rlabel comment s 9540 10486 9540 10486 4 and2_1
rlabel metal1 s 9540 10438 10000 10534 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 9540 10982 10000 11078 1 VPWR
port 6 nsew power bidirectional abutment
flabel locali s 9563 11519 9597 11553 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 10023 11519 10057 11553 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 9655 11451 9689 11485 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel pwell s 9471 11213 9505 11247 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 9471 11757 9505 11791 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 9471 11757 9505 11791 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 9471 11213 9505 11247 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel comment s 9442 11230 9442 11230 4 xor2_1
rlabel metal1 s 9442 11182 10086 11278 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 9442 11726 10086 11822 1 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 9559 12577 9593 12611 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 9559 12033 9593 12067 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel locali s 9927 12203 9961 12237 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 9927 12135 9961 12169 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 9927 12271 9961 12305 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 9927 12339 9961 12373 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 9927 12407 9961 12441 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 9927 12475 9961 12509 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 9743 12271 9777 12305 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 9651 12271 9685 12305 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 9559 12271 9593 12305 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel nwell s 9559 12577 9593 12611 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 9559 12033 9593 12067 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
rlabel comment s 9530 12050 9530 12050 4 and2_1
rlabel metal1 s 9530 12002 9990 12098 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 9530 12546 9990 12642 1 VPWR
port 6 nsew power bidirectional abutment
flabel locali s 9553 13083 9587 13117 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 10013 13083 10047 13117 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 9645 13015 9679 13049 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel pwell s 9461 12777 9495 12811 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 9461 13321 9495 13355 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 9461 13321 9495 13355 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 9461 12777 9495 12811 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel comment s 9432 12794 9432 12794 4 xor2_1
rlabel metal1 s 9432 12746 10076 12842 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 9432 13290 10076 13386 1 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 10935 12371 10969 12405 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 10935 11827 10969 11861 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel locali s 11303 11997 11337 12031 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 11303 11929 11337 11963 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 11303 12065 11337 12099 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 11303 12133 11337 12167 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 11303 12201 11337 12235 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 11303 12269 11337 12303 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 11119 12065 11153 12099 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 11027 12065 11061 12099 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 10935 12065 10969 12099 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel nwell s 10935 12371 10969 12405 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 10935 11827 10969 11861 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
rlabel comment s 10906 11844 10906 11844 4 and2_1
rlabel metal1 s 10906 11796 11366 11892 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 10906 12340 11366 12436 1 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 10939 12847 10973 12881 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 10939 13391 10973 13425 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel locali s 11307 13289 11341 13323 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 11307 12949 11341 12983 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 11123 13289 11157 13323 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 10939 13017 10973 13051 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 11145 13017 11179 13051 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel nwell s 10939 13391 10973 13425 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 10939 12847 10973 12881 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
rlabel comment s 10910 12864 10910 12864 4 and3_1
rlabel metal1 s 10910 12816 11370 12912 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 10910 13360 11370 13456 1 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 9567 14245 9601 14279 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 9567 13701 9601 13735 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel locali s 9935 13871 9969 13905 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 9935 13803 9969 13837 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 9935 13939 9969 13973 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 9935 14007 9969 14041 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 9935 14075 9969 14109 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 9935 14143 9969 14177 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 9751 13939 9785 13973 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 9659 13939 9693 13973 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 9567 13939 9601 13973 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel nwell s 9567 14245 9601 14279 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 9567 13701 9601 13735 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
rlabel comment s 9538 13718 9538 13718 4 and2_1
rlabel metal1 s 9538 13670 9998 13766 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 9538 14214 9998 14310 1 VPWR
port 6 nsew power bidirectional abutment
flabel locali s 11367 14131 11401 14165 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 11091 13791 11125 13825 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 11091 13859 11125 13893 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 10815 13927 10849 13961 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 11091 13927 11125 13961 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 10999 13791 11033 13825 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 10999 13859 11033 13893 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 11183 13927 11217 13961 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel locali s 11367 13791 11401 13825 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 11367 13859 11401 13893 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 11367 13927 11401 13961 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 11367 13995 11401 14029 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 11367 14063 11401 14097 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel metal1 s 10815 13689 10849 13723 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 10815 14233 10849 14267 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel nwell s 10815 14233 10849 14267 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 10815 13689 10849 13723 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
rlabel comment s 10786 13706 10786 13706 4 and4_1
rlabel metal1 s 10786 13658 11430 13754 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 10786 14202 11430 14298 1 VPWR
port 8 nsew power bidirectional abutment
flabel locali s 11969 13553 12003 13587 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 12153 13689 12187 13723 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 11785 13553 11819 13587 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel nwell s 11785 13859 11819 13893 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 11785 13315 11819 13349 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 11785 13315 11819 13349 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 11785 13859 11819 13893 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
rlabel comment s 11756 13332 11756 13332 4 or2_1
rlabel metal1 s 11756 13284 12216 13380 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 11756 13828 12216 13924 1 VPWR
port 6 nsew power bidirectional abutment
flabel locali s 12818 13911 12852 13945 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 12910 13911 12944 13945 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 13094 14047 13128 14081 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 12726 13911 12760 13945 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 12818 14115 12852 14149 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 12726 14115 12760 14149 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 12726 13979 12760 14013 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 12634 14115 12668 14149 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 12818 13979 12852 14013 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 12634 13911 12668 13945 0 FreeSans 400 0 0 0 D
port 4 nsew signal input
flabel locali s 12634 13843 12668 13877 0 FreeSans 400 0 0 0 D
port 4 nsew signal input
flabel metal1 s 12634 14217 12668 14251 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel metal1 s 12634 13673 12668 13707 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel nwell s 12634 14217 12668 14251 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 12634 13673 12668 13707 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
rlabel comment s 12604 13690 12604 13690 4 or4_1
rlabel metal1 s 12604 13642 13156 13738 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 12604 14186 13156 14282 1 VPWR
port 8 nsew power bidirectional abutment
flabel metal1 s 9557 15809 9591 15843 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 9557 15265 9591 15299 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel locali s 9925 15435 9959 15469 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 9925 15367 9959 15401 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 9925 15503 9959 15537 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 9925 15571 9959 15605 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 9925 15639 9959 15673 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 9925 15707 9959 15741 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 9741 15503 9775 15537 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 9649 15503 9683 15537 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 9557 15503 9591 15537 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel nwell s 9557 15809 9591 15843 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 9557 15265 9591 15299 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
rlabel comment s 9528 15282 9528 15282 4 and2_1
rlabel metal1 s 9528 15234 9988 15330 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 9528 15778 9988 15874 1 VPWR
port 6 nsew power bidirectional abutment
flabel locali s 9561 14751 9595 14785 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 10021 14751 10055 14785 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 9653 14683 9687 14717 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel pwell s 9469 14445 9503 14479 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 9469 14989 9503 15023 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 9469 14989 9503 15023 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 9469 14445 9503 14479 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel comment s 9440 14462 9440 14462 4 xor2_1
rlabel metal1 s 9440 14414 10084 14510 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 9440 14958 10084 15054 1 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 10741 15199 10775 15233 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 10741 14655 10775 14689 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel locali s 11109 14825 11143 14859 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 11109 14757 11143 14791 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 11109 14893 11143 14927 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 11109 14961 11143 14995 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 11109 15029 11143 15063 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 11109 15097 11143 15131 0 FreeSans 250 0 0 0 X
port 7 nsew signal output
flabel locali s 10925 14893 10959 14927 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel locali s 10833 14893 10867 14927 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 10741 14893 10775 14927 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel nwell s 10741 15199 10775 15233 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 10741 14655 10775 14689 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
rlabel comment s 10712 14672 10712 14672 4 and2_1
rlabel metal1 s 10712 14624 11172 14720 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 10712 15168 11172 15264 1 VPWR
port 6 nsew power bidirectional abutment
flabel locali s 12151 15597 12185 15631 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 11875 15257 11909 15291 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 11875 15325 11909 15359 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 11599 15393 11633 15427 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 11875 15393 11909 15427 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 11783 15257 11817 15291 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 11783 15325 11817 15359 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 11967 15393 12001 15427 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel locali s 12151 15257 12185 15291 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 12151 15325 12185 15359 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 12151 15393 12185 15427 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 12151 15461 12185 15495 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 12151 15529 12185 15563 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel metal1 s 11599 15155 11633 15189 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 11599 15699 11633 15733 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel nwell s 11599 15699 11633 15733 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 11599 15155 11633 15189 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
rlabel comment s 11570 15172 11570 15172 4 and4_1
rlabel metal1 s 11570 15124 12214 15220 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 11570 15668 12214 15764 1 VPWR
port 8 nsew power bidirectional abutment
flabel locali s 9551 16315 9585 16349 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 10011 16315 10045 16349 0 FreeSans 200 0 0 0 X
port 7 nsew signal output
flabel locali s 9643 16247 9677 16281 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel pwell s 9459 16009 9493 16043 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 9459 16553 9493 16587 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 9459 16553 9493 16587 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 9459 16009 9493 16043 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel comment s 9430 16026 9430 16026 4 xor2_1
rlabel metal1 s 9430 15978 10074 16074 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 9430 16522 10074 16618 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
