magic
tech sky130A
magscale 1 2
timestamp 1754942322
<< nwell >>
rect 9296 16307 10016 16628
rect 9394 15563 9930 15884
rect 11436 15453 12156 15774
rect 9306 14743 10026 15064
rect 10578 14953 11114 15274
rect 9404 13999 9940 14320
rect 10652 13987 11372 14308
rect 12550 13971 13178 14292
rect 11622 13613 12158 13934
rect 9298 13075 10018 13396
rect 10776 13145 11312 13466
rect 9396 12331 9932 12652
rect 10772 12125 11308 12446
rect 9308 11511 10028 11832
rect 9406 10767 9942 11088
rect 6074 6018 6426 6339
rect 9980 5386 11528 5707
rect 12042 5374 13588 5695
rect 14000 5382 15546 5703
rect 15994 5388 17542 5709
rect 1798 4966 3346 5287
rect 3932 4958 5480 5279
rect 5884 4958 7432 5279
rect 7886 4964 9434 5285
rect 10008 4512 11556 4833
rect 12278 4468 13826 4789
rect 14280 4462 15828 4783
rect 16302 4444 17850 4765
rect 1768 1706 3316 2027
rect 3838 1702 5386 2023
rect 5790 1702 7338 2023
rect 7792 1708 9340 2029
rect 9744 1708 11292 2029
rect 11736 1708 13284 2029
rect 13688 1708 15236 2029
rect 15752 1708 17300 2029
<< pwell >>
rect 9343 16067 9977 16249
rect 9363 16029 9397 16067
rect 9661 15487 9851 15505
rect 9465 15323 9851 15487
rect 11890 15349 12117 15395
rect 9465 15319 9495 15323
rect 9461 15285 9495 15319
rect 11475 15213 12117 15349
rect 11503 15175 11537 15213
rect 10845 14877 11035 14895
rect 10649 14713 11035 14877
rect 10649 14709 10679 14713
rect 9353 14503 9987 14685
rect 10645 14675 10679 14709
rect 9373 14465 9407 14503
rect 9671 13923 9861 13941
rect 9475 13759 9861 13923
rect 11106 13883 11333 13929
rect 9475 13755 9505 13759
rect 9471 13721 9505 13755
rect 10691 13747 11333 13883
rect 10719 13709 10753 13747
rect 12950 13873 13139 13913
rect 12589 13737 13139 13873
rect 12618 13693 12652 13737
rect 12950 13731 13139 13737
rect 11871 13509 12057 13555
rect 11690 13373 12057 13509
rect 11690 13369 11723 13373
rect 11689 13335 11723 13369
rect 11089 13041 11273 13087
rect 9345 12835 9979 13017
rect 10815 12905 11273 13041
rect 10843 12867 10877 12905
rect 9365 12797 9399 12835
rect 9663 12255 9853 12273
rect 9467 12091 9853 12255
rect 9467 12087 9497 12091
rect 9463 12053 9497 12087
rect 11039 12049 11229 12067
rect 10843 11885 11229 12049
rect 10843 11881 10873 11885
rect 10839 11847 10873 11881
rect 9355 11271 9989 11453
rect 9375 11233 9409 11271
rect 9673 10691 9863 10709
rect 9477 10527 9863 10691
rect 9477 10523 9507 10527
rect 9473 10489 9507 10523
rect 6325 6583 6359 6617
rect 6325 6579 6346 6583
rect 6160 6397 6346 6579
rect 11426 5947 11460 5985
rect 10054 5811 11489 5947
rect 13488 5935 13522 5973
rect 15446 5943 15480 5981
rect 17440 5949 17474 5987
rect 10054 5765 10240 5811
rect 11303 5765 11489 5811
rect 12116 5799 13551 5935
rect 12116 5753 12302 5799
rect 13365 5753 13551 5799
rect 14074 5807 15509 5943
rect 14074 5761 14260 5807
rect 15323 5761 15509 5807
rect 16068 5813 17503 5949
rect 16068 5767 16254 5813
rect 17317 5767 17503 5813
rect 3244 5527 3278 5565
rect 1872 5391 3307 5527
rect 5378 5519 5412 5557
rect 7330 5519 7364 5557
rect 9332 5525 9366 5563
rect 1872 5345 2058 5391
rect 3121 5345 3307 5391
rect 4006 5383 5441 5519
rect 4006 5337 4192 5383
rect 5255 5337 5441 5383
rect 5958 5383 7393 5519
rect 5958 5337 6144 5383
rect 7207 5337 7393 5383
rect 7960 5389 9395 5525
rect 7960 5343 8146 5389
rect 9209 5343 9395 5389
rect 11454 5073 11488 5111
rect 10082 4937 11517 5073
rect 13724 5029 13758 5067
rect 10082 4891 10268 4937
rect 11331 4891 11517 4937
rect 12352 4893 13787 5029
rect 15726 5023 15760 5061
rect 12352 4847 12538 4893
rect 13601 4847 13787 4893
rect 14354 4887 15789 5023
rect 17748 5005 17782 5043
rect 14354 4841 14540 4887
rect 15603 4841 15789 4887
rect 16376 4869 17811 5005
rect 16376 4823 16562 4869
rect 17625 4823 17811 4869
rect 3214 2267 3248 2305
rect 1842 2131 3277 2267
rect 5284 2263 5318 2301
rect 7236 2263 7270 2301
rect 9238 2269 9272 2307
rect 11190 2269 11224 2307
rect 13182 2269 13216 2307
rect 15134 2269 15168 2307
rect 17198 2269 17232 2307
rect 1842 2085 2028 2131
rect 3091 2085 3277 2131
rect 3912 2127 5347 2263
rect 3912 2081 4098 2127
rect 5161 2081 5347 2127
rect 5864 2127 7299 2263
rect 5864 2081 6050 2127
rect 7113 2081 7299 2127
rect 7866 2133 9301 2269
rect 7866 2087 8052 2133
rect 9115 2087 9301 2133
rect 9818 2133 11253 2269
rect 9818 2087 10004 2133
rect 11067 2087 11253 2133
rect 11810 2133 13245 2269
rect 11810 2087 11996 2133
rect 13059 2087 13245 2133
rect 13762 2133 15197 2269
rect 13762 2087 13948 2133
rect 15011 2087 15197 2133
rect 15826 2133 17261 2269
rect 15826 2087 16012 2133
rect 17075 2087 17261 2133
<< ndiff >>
rect 9369 16141 9421 16223
rect 9369 16107 9377 16141
rect 9411 16107 9421 16141
rect 9369 16093 9421 16107
rect 9451 16163 9505 16223
rect 9451 16129 9461 16163
rect 9495 16129 9505 16163
rect 9451 16093 9505 16129
rect 9535 16141 9589 16223
rect 9535 16107 9545 16141
rect 9579 16107 9589 16141
rect 9535 16093 9589 16107
rect 9619 16093 9673 16223
rect 9703 16143 9857 16223
rect 9703 16109 9713 16143
rect 9747 16109 9813 16143
rect 9847 16109 9857 16143
rect 9703 16093 9857 16109
rect 9887 16214 9951 16223
rect 9887 16180 9903 16214
rect 9937 16180 9951 16214
rect 9887 16146 9951 16180
rect 9887 16112 9903 16146
rect 9937 16112 9951 16146
rect 9887 16093 9951 16112
rect 9687 15461 9739 15479
rect 9491 15423 9547 15461
rect 9491 15389 9503 15423
rect 9537 15389 9547 15423
rect 9491 15377 9547 15389
rect 9577 15377 9631 15461
rect 9661 15395 9739 15461
rect 9661 15377 9695 15395
rect 9687 15361 9695 15377
rect 9729 15361 9739 15395
rect 9687 15349 9739 15361
rect 9769 15395 9825 15479
rect 9769 15361 9779 15395
rect 9813 15361 9825 15395
rect 9769 15349 9825 15361
rect 11916 15353 12009 15369
rect 11916 15323 11950 15353
rect 11501 15293 11553 15323
rect 11501 15259 11509 15293
rect 11543 15259 11553 15293
rect 11501 15239 11553 15259
rect 11583 15239 11641 15323
rect 11671 15239 11747 15323
rect 11777 15239 11843 15323
rect 11873 15319 11950 15323
rect 11984 15319 12009 15353
rect 11873 15285 12009 15319
rect 11873 15251 11950 15285
rect 11984 15251 12009 15285
rect 11873 15239 12009 15251
rect 12039 15353 12091 15369
rect 12039 15319 12049 15353
rect 12083 15319 12091 15353
rect 12039 15285 12091 15319
rect 12039 15251 12049 15285
rect 12083 15251 12091 15285
rect 12039 15239 12091 15251
rect 10871 14851 10923 14869
rect 10675 14813 10731 14851
rect 10675 14779 10687 14813
rect 10721 14779 10731 14813
rect 10675 14767 10731 14779
rect 10761 14767 10815 14851
rect 10845 14785 10923 14851
rect 10845 14767 10879 14785
rect 10871 14751 10879 14767
rect 10913 14751 10923 14785
rect 10871 14739 10923 14751
rect 10953 14785 11009 14869
rect 10953 14751 10963 14785
rect 10997 14751 11009 14785
rect 10953 14739 11009 14751
rect 9379 14577 9431 14659
rect 9379 14543 9387 14577
rect 9421 14543 9431 14577
rect 9379 14529 9431 14543
rect 9461 14599 9515 14659
rect 9461 14565 9471 14599
rect 9505 14565 9515 14599
rect 9461 14529 9515 14565
rect 9545 14577 9599 14659
rect 9545 14543 9555 14577
rect 9589 14543 9599 14577
rect 9545 14529 9599 14543
rect 9629 14529 9683 14659
rect 9713 14579 9867 14659
rect 9713 14545 9723 14579
rect 9757 14545 9823 14579
rect 9857 14545 9867 14579
rect 9713 14529 9867 14545
rect 9897 14650 9961 14659
rect 9897 14616 9913 14650
rect 9947 14616 9961 14650
rect 9897 14582 9961 14616
rect 9897 14548 9913 14582
rect 9947 14548 9961 14582
rect 9897 14529 9961 14548
rect 9697 13897 9749 13915
rect 9501 13859 9557 13897
rect 9501 13825 9513 13859
rect 9547 13825 9557 13859
rect 9501 13813 9557 13825
rect 9587 13813 9641 13897
rect 9671 13831 9749 13897
rect 9671 13813 9705 13831
rect 9697 13797 9705 13813
rect 9739 13797 9749 13831
rect 9697 13785 9749 13797
rect 9779 13831 9835 13915
rect 11132 13887 11225 13903
rect 11132 13857 11166 13887
rect 9779 13797 9789 13831
rect 9823 13797 9835 13831
rect 9779 13785 9835 13797
rect 10717 13827 10769 13857
rect 10717 13793 10725 13827
rect 10759 13793 10769 13827
rect 10717 13773 10769 13793
rect 10799 13773 10857 13857
rect 10887 13773 10963 13857
rect 10993 13773 11059 13857
rect 11089 13853 11166 13857
rect 11200 13853 11225 13887
rect 11089 13819 11225 13853
rect 11089 13785 11166 13819
rect 11200 13785 11225 13819
rect 11089 13773 11225 13785
rect 11255 13887 11307 13903
rect 11255 13853 11265 13887
rect 11299 13853 11307 13887
rect 11255 13819 11307 13853
rect 11255 13785 11265 13819
rect 11299 13785 11307 13819
rect 11255 13773 11307 13785
rect 12976 13847 13029 13887
rect 12615 13827 12667 13847
rect 12615 13793 12623 13827
rect 12657 13793 12667 13827
rect 12615 13763 12667 13793
rect 12697 13821 12763 13847
rect 12697 13787 12713 13821
rect 12747 13787 12763 13821
rect 12697 13763 12763 13787
rect 12793 13807 12847 13847
rect 12793 13773 12803 13807
rect 12837 13773 12847 13807
rect 12793 13763 12847 13773
rect 12877 13821 12931 13847
rect 12877 13787 12887 13821
rect 12921 13787 12931 13821
rect 12877 13763 12931 13787
rect 12961 13807 13029 13847
rect 12961 13773 12981 13807
rect 13015 13773 13029 13807
rect 12961 13763 13029 13773
rect 12976 13757 13029 13763
rect 13059 13845 13113 13887
rect 13059 13811 13069 13845
rect 13103 13811 13113 13845
rect 13059 13757 13113 13811
rect 11897 13483 11949 13529
rect 11716 13455 11768 13483
rect 11716 13421 11724 13455
rect 11758 13421 11768 13455
rect 11716 13399 11768 13421
rect 11798 13455 11852 13483
rect 11798 13421 11808 13455
rect 11842 13421 11852 13455
rect 11798 13399 11852 13421
rect 11882 13455 11949 13483
rect 11882 13421 11904 13455
rect 11938 13421 11949 13455
rect 11882 13399 11949 13421
rect 11979 13515 12031 13529
rect 11979 13481 11989 13515
rect 12023 13481 12031 13515
rect 11979 13447 12031 13481
rect 11979 13413 11989 13447
rect 12023 13413 12031 13447
rect 11979 13399 12031 13413
rect 11115 13015 11165 13061
rect 9371 12909 9423 12991
rect 9371 12875 9379 12909
rect 9413 12875 9423 12909
rect 9371 12861 9423 12875
rect 9453 12931 9507 12991
rect 9453 12897 9463 12931
rect 9497 12897 9507 12931
rect 9453 12861 9507 12897
rect 9537 12909 9591 12991
rect 9537 12875 9547 12909
rect 9581 12875 9591 12909
rect 9537 12861 9591 12875
rect 9621 12861 9675 12991
rect 9705 12911 9859 12991
rect 9705 12877 9715 12911
rect 9749 12877 9815 12911
rect 9849 12877 9859 12911
rect 9705 12861 9859 12877
rect 9889 12982 9953 12991
rect 9889 12948 9905 12982
rect 9939 12948 9953 12982
rect 9889 12914 9953 12948
rect 10841 12977 10893 13015
rect 10841 12943 10849 12977
rect 10883 12943 10893 12977
rect 10841 12931 10893 12943
rect 10923 12931 10965 13015
rect 10995 12931 11037 13015
rect 11067 12993 11165 13015
rect 11067 12959 11121 12993
rect 11155 12959 11165 12993
rect 11067 12931 11165 12959
rect 11195 13003 11247 13061
rect 11195 12969 11205 13003
rect 11239 12969 11247 13003
rect 11195 12931 11247 12969
rect 9889 12880 9905 12914
rect 9939 12880 9953 12914
rect 9889 12861 9953 12880
rect 9689 12229 9741 12247
rect 9493 12191 9549 12229
rect 9493 12157 9505 12191
rect 9539 12157 9549 12191
rect 9493 12145 9549 12157
rect 9579 12145 9633 12229
rect 9663 12163 9741 12229
rect 9663 12145 9697 12163
rect 9689 12129 9697 12145
rect 9731 12129 9741 12163
rect 9689 12117 9741 12129
rect 9771 12163 9827 12247
rect 9771 12129 9781 12163
rect 9815 12129 9827 12163
rect 9771 12117 9827 12129
rect 11065 12023 11117 12041
rect 10869 11985 10925 12023
rect 10869 11951 10881 11985
rect 10915 11951 10925 11985
rect 10869 11939 10925 11951
rect 10955 11939 11009 12023
rect 11039 11957 11117 12023
rect 11039 11939 11073 11957
rect 11065 11923 11073 11939
rect 11107 11923 11117 11957
rect 11065 11911 11117 11923
rect 11147 11957 11203 12041
rect 11147 11923 11157 11957
rect 11191 11923 11203 11957
rect 11147 11911 11203 11923
rect 9381 11345 9433 11427
rect 9381 11311 9389 11345
rect 9423 11311 9433 11345
rect 9381 11297 9433 11311
rect 9463 11367 9517 11427
rect 9463 11333 9473 11367
rect 9507 11333 9517 11367
rect 9463 11297 9517 11333
rect 9547 11345 9601 11427
rect 9547 11311 9557 11345
rect 9591 11311 9601 11345
rect 9547 11297 9601 11311
rect 9631 11297 9685 11427
rect 9715 11347 9869 11427
rect 9715 11313 9725 11347
rect 9759 11313 9825 11347
rect 9859 11313 9869 11347
rect 9715 11297 9869 11313
rect 9899 11418 9963 11427
rect 9899 11384 9915 11418
rect 9949 11384 9963 11418
rect 9899 11350 9963 11384
rect 9899 11316 9915 11350
rect 9949 11316 9963 11350
rect 9899 11297 9963 11316
rect 9699 10665 9751 10683
rect 9503 10627 9559 10665
rect 9503 10593 9515 10627
rect 9549 10593 9559 10627
rect 9503 10581 9559 10593
rect 9589 10581 9643 10665
rect 9673 10599 9751 10665
rect 9673 10581 9707 10599
rect 9699 10565 9707 10581
rect 9741 10565 9751 10599
rect 9699 10553 9751 10565
rect 9781 10599 9837 10683
rect 9781 10565 9791 10599
rect 9825 10565 9837 10599
rect 9781 10553 9837 10565
rect 6186 6537 6238 6553
rect 6186 6503 6194 6537
rect 6228 6503 6238 6537
rect 6186 6469 6238 6503
rect 6186 6435 6194 6469
rect 6228 6435 6238 6469
rect 6186 6423 6238 6435
rect 6268 6537 6320 6553
rect 6268 6503 6278 6537
rect 6312 6503 6320 6537
rect 6268 6469 6320 6503
rect 6268 6435 6278 6469
rect 6312 6435 6320 6469
rect 6268 6423 6320 6435
rect 10080 5873 10132 5921
rect 10080 5839 10088 5873
rect 10122 5839 10132 5873
rect 10080 5791 10132 5839
rect 10162 5913 10231 5921
rect 10162 5879 10187 5913
rect 10221 5879 10231 5913
rect 10162 5837 10231 5879
rect 10261 5837 10327 5921
rect 10357 5837 10399 5921
rect 10429 5901 10495 5921
rect 10429 5867 10439 5901
rect 10473 5867 10495 5901
rect 10429 5837 10495 5867
rect 10525 5896 10584 5921
rect 10525 5862 10540 5896
rect 10574 5862 10584 5896
rect 10525 5837 10584 5862
rect 10614 5913 10668 5921
rect 10614 5879 10624 5913
rect 10658 5879 10668 5913
rect 10614 5837 10668 5879
rect 10698 5896 10752 5921
rect 10698 5862 10708 5896
rect 10742 5862 10752 5896
rect 10698 5837 10752 5862
rect 10782 5904 10834 5921
rect 10782 5870 10792 5904
rect 10826 5870 10834 5904
rect 10782 5837 10834 5870
rect 10888 5896 10940 5921
rect 10888 5862 10896 5896
rect 10930 5862 10940 5896
rect 10888 5837 10940 5862
rect 10970 5913 11024 5921
rect 10970 5879 10980 5913
rect 11014 5879 11024 5913
rect 10970 5837 11024 5879
rect 11054 5896 11108 5921
rect 11054 5862 11064 5896
rect 11098 5862 11108 5896
rect 11054 5837 11108 5862
rect 11138 5896 11192 5921
rect 11138 5862 11148 5896
rect 11182 5862 11192 5896
rect 11138 5837 11192 5862
rect 11222 5837 11282 5921
rect 11312 5909 11381 5921
rect 11312 5875 11337 5909
rect 11371 5875 11381 5909
rect 11312 5837 11381 5875
rect 10162 5791 10214 5837
rect 1898 5453 1950 5501
rect 1898 5419 1906 5453
rect 1940 5419 1950 5453
rect 1898 5371 1950 5419
rect 1980 5493 2049 5501
rect 1980 5459 2005 5493
rect 2039 5459 2049 5493
rect 1980 5417 2049 5459
rect 2079 5417 2145 5501
rect 2175 5417 2217 5501
rect 2247 5481 2313 5501
rect 2247 5447 2257 5481
rect 2291 5447 2313 5481
rect 2247 5417 2313 5447
rect 2343 5476 2402 5501
rect 2343 5442 2358 5476
rect 2392 5442 2402 5476
rect 2343 5417 2402 5442
rect 2432 5493 2486 5501
rect 2432 5459 2442 5493
rect 2476 5459 2486 5493
rect 2432 5417 2486 5459
rect 2516 5476 2570 5501
rect 2516 5442 2526 5476
rect 2560 5442 2570 5476
rect 2516 5417 2570 5442
rect 2600 5484 2652 5501
rect 2600 5450 2610 5484
rect 2644 5450 2652 5484
rect 2600 5417 2652 5450
rect 2706 5476 2758 5501
rect 2706 5442 2714 5476
rect 2748 5442 2758 5476
rect 2706 5417 2758 5442
rect 2788 5493 2842 5501
rect 2788 5459 2798 5493
rect 2832 5459 2842 5493
rect 2788 5417 2842 5459
rect 2872 5476 2926 5501
rect 2872 5442 2882 5476
rect 2916 5442 2926 5476
rect 2872 5417 2926 5442
rect 2956 5476 3010 5501
rect 2956 5442 2966 5476
rect 3000 5442 3010 5476
rect 2956 5417 3010 5442
rect 3040 5417 3100 5501
rect 3130 5489 3199 5501
rect 3130 5455 3155 5489
rect 3189 5455 3199 5489
rect 3130 5417 3199 5455
rect 1980 5371 2032 5417
rect 3147 5371 3199 5417
rect 3229 5453 3281 5501
rect 3229 5419 3239 5453
rect 3273 5419 3281 5453
rect 3229 5371 3281 5419
rect 4032 5445 4084 5493
rect 4032 5411 4040 5445
rect 4074 5411 4084 5445
rect 4032 5363 4084 5411
rect 4114 5485 4183 5493
rect 4114 5451 4139 5485
rect 4173 5451 4183 5485
rect 4114 5409 4183 5451
rect 4213 5409 4279 5493
rect 4309 5409 4351 5493
rect 4381 5473 4447 5493
rect 4381 5439 4391 5473
rect 4425 5439 4447 5473
rect 4381 5409 4447 5439
rect 4477 5468 4536 5493
rect 4477 5434 4492 5468
rect 4526 5434 4536 5468
rect 4477 5409 4536 5434
rect 4566 5485 4620 5493
rect 4566 5451 4576 5485
rect 4610 5451 4620 5485
rect 4566 5409 4620 5451
rect 4650 5468 4704 5493
rect 4650 5434 4660 5468
rect 4694 5434 4704 5468
rect 4650 5409 4704 5434
rect 4734 5476 4786 5493
rect 4734 5442 4744 5476
rect 4778 5442 4786 5476
rect 4734 5409 4786 5442
rect 4840 5468 4892 5493
rect 4840 5434 4848 5468
rect 4882 5434 4892 5468
rect 4840 5409 4892 5434
rect 4922 5485 4976 5493
rect 4922 5451 4932 5485
rect 4966 5451 4976 5485
rect 4922 5409 4976 5451
rect 5006 5468 5060 5493
rect 5006 5434 5016 5468
rect 5050 5434 5060 5468
rect 5006 5409 5060 5434
rect 5090 5468 5144 5493
rect 5090 5434 5100 5468
rect 5134 5434 5144 5468
rect 5090 5409 5144 5434
rect 5174 5409 5234 5493
rect 5264 5481 5333 5493
rect 5264 5447 5289 5481
rect 5323 5447 5333 5481
rect 5264 5409 5333 5447
rect 4114 5363 4166 5409
rect 5281 5363 5333 5409
rect 5363 5445 5415 5493
rect 5363 5411 5373 5445
rect 5407 5411 5415 5445
rect 5363 5363 5415 5411
rect 5984 5445 6036 5493
rect 5984 5411 5992 5445
rect 6026 5411 6036 5445
rect 5984 5363 6036 5411
rect 6066 5485 6135 5493
rect 6066 5451 6091 5485
rect 6125 5451 6135 5485
rect 6066 5409 6135 5451
rect 6165 5409 6231 5493
rect 6261 5409 6303 5493
rect 6333 5473 6399 5493
rect 6333 5439 6343 5473
rect 6377 5439 6399 5473
rect 6333 5409 6399 5439
rect 6429 5468 6488 5493
rect 6429 5434 6444 5468
rect 6478 5434 6488 5468
rect 6429 5409 6488 5434
rect 6518 5485 6572 5493
rect 6518 5451 6528 5485
rect 6562 5451 6572 5485
rect 6518 5409 6572 5451
rect 6602 5468 6656 5493
rect 6602 5434 6612 5468
rect 6646 5434 6656 5468
rect 6602 5409 6656 5434
rect 6686 5476 6738 5493
rect 6686 5442 6696 5476
rect 6730 5442 6738 5476
rect 6686 5409 6738 5442
rect 6792 5468 6844 5493
rect 6792 5434 6800 5468
rect 6834 5434 6844 5468
rect 6792 5409 6844 5434
rect 6874 5485 6928 5493
rect 6874 5451 6884 5485
rect 6918 5451 6928 5485
rect 6874 5409 6928 5451
rect 6958 5468 7012 5493
rect 6958 5434 6968 5468
rect 7002 5434 7012 5468
rect 6958 5409 7012 5434
rect 7042 5468 7096 5493
rect 7042 5434 7052 5468
rect 7086 5434 7096 5468
rect 7042 5409 7096 5434
rect 7126 5409 7186 5493
rect 7216 5481 7285 5493
rect 7216 5447 7241 5481
rect 7275 5447 7285 5481
rect 7216 5409 7285 5447
rect 6066 5363 6118 5409
rect 7233 5363 7285 5409
rect 7315 5445 7367 5493
rect 7315 5411 7325 5445
rect 7359 5411 7367 5445
rect 7315 5363 7367 5411
rect 7986 5451 8038 5499
rect 7986 5417 7994 5451
rect 8028 5417 8038 5451
rect 7986 5369 8038 5417
rect 8068 5491 8137 5499
rect 8068 5457 8093 5491
rect 8127 5457 8137 5491
rect 8068 5415 8137 5457
rect 8167 5415 8233 5499
rect 8263 5415 8305 5499
rect 8335 5479 8401 5499
rect 8335 5445 8345 5479
rect 8379 5445 8401 5479
rect 8335 5415 8401 5445
rect 8431 5474 8490 5499
rect 8431 5440 8446 5474
rect 8480 5440 8490 5474
rect 8431 5415 8490 5440
rect 8520 5491 8574 5499
rect 8520 5457 8530 5491
rect 8564 5457 8574 5491
rect 8520 5415 8574 5457
rect 8604 5474 8658 5499
rect 8604 5440 8614 5474
rect 8648 5440 8658 5474
rect 8604 5415 8658 5440
rect 8688 5482 8740 5499
rect 8688 5448 8698 5482
rect 8732 5448 8740 5482
rect 8688 5415 8740 5448
rect 8794 5474 8846 5499
rect 8794 5440 8802 5474
rect 8836 5440 8846 5474
rect 8794 5415 8846 5440
rect 8876 5491 8930 5499
rect 8876 5457 8886 5491
rect 8920 5457 8930 5491
rect 8876 5415 8930 5457
rect 8960 5474 9014 5499
rect 8960 5440 8970 5474
rect 9004 5440 9014 5474
rect 8960 5415 9014 5440
rect 9044 5474 9098 5499
rect 9044 5440 9054 5474
rect 9088 5440 9098 5474
rect 9044 5415 9098 5440
rect 9128 5415 9188 5499
rect 9218 5487 9287 5499
rect 9218 5453 9243 5487
rect 9277 5453 9287 5487
rect 9218 5415 9287 5453
rect 8068 5369 8120 5415
rect 9235 5369 9287 5415
rect 9317 5451 9369 5499
rect 11329 5791 11381 5837
rect 11411 5873 11463 5921
rect 11411 5839 11421 5873
rect 11455 5839 11463 5873
rect 11411 5791 11463 5839
rect 12142 5861 12194 5909
rect 12142 5827 12150 5861
rect 12184 5827 12194 5861
rect 12142 5779 12194 5827
rect 12224 5901 12293 5909
rect 12224 5867 12249 5901
rect 12283 5867 12293 5901
rect 12224 5825 12293 5867
rect 12323 5825 12389 5909
rect 12419 5825 12461 5909
rect 12491 5889 12557 5909
rect 12491 5855 12501 5889
rect 12535 5855 12557 5889
rect 12491 5825 12557 5855
rect 12587 5884 12646 5909
rect 12587 5850 12602 5884
rect 12636 5850 12646 5884
rect 12587 5825 12646 5850
rect 12676 5901 12730 5909
rect 12676 5867 12686 5901
rect 12720 5867 12730 5901
rect 12676 5825 12730 5867
rect 12760 5884 12814 5909
rect 12760 5850 12770 5884
rect 12804 5850 12814 5884
rect 12760 5825 12814 5850
rect 12844 5892 12896 5909
rect 12844 5858 12854 5892
rect 12888 5858 12896 5892
rect 12844 5825 12896 5858
rect 12950 5884 13002 5909
rect 12950 5850 12958 5884
rect 12992 5850 13002 5884
rect 12950 5825 13002 5850
rect 13032 5901 13086 5909
rect 13032 5867 13042 5901
rect 13076 5867 13086 5901
rect 13032 5825 13086 5867
rect 13116 5884 13170 5909
rect 13116 5850 13126 5884
rect 13160 5850 13170 5884
rect 13116 5825 13170 5850
rect 13200 5884 13254 5909
rect 13200 5850 13210 5884
rect 13244 5850 13254 5884
rect 13200 5825 13254 5850
rect 13284 5825 13344 5909
rect 13374 5897 13443 5909
rect 13374 5863 13399 5897
rect 13433 5863 13443 5897
rect 13374 5825 13443 5863
rect 12224 5779 12276 5825
rect 9317 5417 9327 5451
rect 9361 5417 9369 5451
rect 13391 5779 13443 5825
rect 13473 5861 13525 5909
rect 13473 5827 13483 5861
rect 13517 5827 13525 5861
rect 13473 5779 13525 5827
rect 14100 5869 14152 5917
rect 14100 5835 14108 5869
rect 14142 5835 14152 5869
rect 14100 5787 14152 5835
rect 14182 5909 14251 5917
rect 14182 5875 14207 5909
rect 14241 5875 14251 5909
rect 14182 5833 14251 5875
rect 14281 5833 14347 5917
rect 14377 5833 14419 5917
rect 14449 5897 14515 5917
rect 14449 5863 14459 5897
rect 14493 5863 14515 5897
rect 14449 5833 14515 5863
rect 14545 5892 14604 5917
rect 14545 5858 14560 5892
rect 14594 5858 14604 5892
rect 14545 5833 14604 5858
rect 14634 5909 14688 5917
rect 14634 5875 14644 5909
rect 14678 5875 14688 5909
rect 14634 5833 14688 5875
rect 14718 5892 14772 5917
rect 14718 5858 14728 5892
rect 14762 5858 14772 5892
rect 14718 5833 14772 5858
rect 14802 5900 14854 5917
rect 14802 5866 14812 5900
rect 14846 5866 14854 5900
rect 14802 5833 14854 5866
rect 14908 5892 14960 5917
rect 14908 5858 14916 5892
rect 14950 5858 14960 5892
rect 14908 5833 14960 5858
rect 14990 5909 15044 5917
rect 14990 5875 15000 5909
rect 15034 5875 15044 5909
rect 14990 5833 15044 5875
rect 15074 5892 15128 5917
rect 15074 5858 15084 5892
rect 15118 5858 15128 5892
rect 15074 5833 15128 5858
rect 15158 5892 15212 5917
rect 15158 5858 15168 5892
rect 15202 5858 15212 5892
rect 15158 5833 15212 5858
rect 15242 5833 15302 5917
rect 15332 5905 15401 5917
rect 15332 5871 15357 5905
rect 15391 5871 15401 5905
rect 15332 5833 15401 5871
rect 14182 5787 14234 5833
rect 15349 5787 15401 5833
rect 15431 5869 15483 5917
rect 15431 5835 15441 5869
rect 15475 5835 15483 5869
rect 15431 5787 15483 5835
rect 16094 5875 16146 5923
rect 16094 5841 16102 5875
rect 16136 5841 16146 5875
rect 16094 5793 16146 5841
rect 16176 5915 16245 5923
rect 16176 5881 16201 5915
rect 16235 5881 16245 5915
rect 16176 5839 16245 5881
rect 16275 5839 16341 5923
rect 16371 5839 16413 5923
rect 16443 5903 16509 5923
rect 16443 5869 16453 5903
rect 16487 5869 16509 5903
rect 16443 5839 16509 5869
rect 16539 5898 16598 5923
rect 16539 5864 16554 5898
rect 16588 5864 16598 5898
rect 16539 5839 16598 5864
rect 16628 5915 16682 5923
rect 16628 5881 16638 5915
rect 16672 5881 16682 5915
rect 16628 5839 16682 5881
rect 16712 5898 16766 5923
rect 16712 5864 16722 5898
rect 16756 5864 16766 5898
rect 16712 5839 16766 5864
rect 16796 5906 16848 5923
rect 16796 5872 16806 5906
rect 16840 5872 16848 5906
rect 16796 5839 16848 5872
rect 16902 5898 16954 5923
rect 16902 5864 16910 5898
rect 16944 5864 16954 5898
rect 16902 5839 16954 5864
rect 16984 5915 17038 5923
rect 16984 5881 16994 5915
rect 17028 5881 17038 5915
rect 16984 5839 17038 5881
rect 17068 5898 17122 5923
rect 17068 5864 17078 5898
rect 17112 5864 17122 5898
rect 17068 5839 17122 5864
rect 17152 5898 17206 5923
rect 17152 5864 17162 5898
rect 17196 5864 17206 5898
rect 17152 5839 17206 5864
rect 17236 5839 17296 5923
rect 17326 5911 17395 5923
rect 17326 5877 17351 5911
rect 17385 5877 17395 5911
rect 17326 5839 17395 5877
rect 16176 5793 16228 5839
rect 17343 5793 17395 5839
rect 17425 5875 17477 5923
rect 17425 5841 17435 5875
rect 17469 5841 17477 5875
rect 17425 5793 17477 5841
rect 9317 5369 9369 5417
rect 10108 4999 10160 5047
rect 10108 4965 10116 4999
rect 10150 4965 10160 4999
rect 10108 4917 10160 4965
rect 10190 5039 10259 5047
rect 10190 5005 10215 5039
rect 10249 5005 10259 5039
rect 10190 4963 10259 5005
rect 10289 4963 10355 5047
rect 10385 4963 10427 5047
rect 10457 5027 10523 5047
rect 10457 4993 10467 5027
rect 10501 4993 10523 5027
rect 10457 4963 10523 4993
rect 10553 5022 10612 5047
rect 10553 4988 10568 5022
rect 10602 4988 10612 5022
rect 10553 4963 10612 4988
rect 10642 5039 10696 5047
rect 10642 5005 10652 5039
rect 10686 5005 10696 5039
rect 10642 4963 10696 5005
rect 10726 5022 10780 5047
rect 10726 4988 10736 5022
rect 10770 4988 10780 5022
rect 10726 4963 10780 4988
rect 10810 5030 10862 5047
rect 10810 4996 10820 5030
rect 10854 4996 10862 5030
rect 10810 4963 10862 4996
rect 10916 5022 10968 5047
rect 10916 4988 10924 5022
rect 10958 4988 10968 5022
rect 10916 4963 10968 4988
rect 10998 5039 11052 5047
rect 10998 5005 11008 5039
rect 11042 5005 11052 5039
rect 10998 4963 11052 5005
rect 11082 5022 11136 5047
rect 11082 4988 11092 5022
rect 11126 4988 11136 5022
rect 11082 4963 11136 4988
rect 11166 5022 11220 5047
rect 11166 4988 11176 5022
rect 11210 4988 11220 5022
rect 11166 4963 11220 4988
rect 11250 4963 11310 5047
rect 11340 5035 11409 5047
rect 11340 5001 11365 5035
rect 11399 5001 11409 5035
rect 11340 4963 11409 5001
rect 10190 4917 10242 4963
rect 11357 4917 11409 4963
rect 11439 4999 11491 5047
rect 11439 4965 11449 4999
rect 11483 4965 11491 4999
rect 11439 4917 11491 4965
rect 12378 4955 12430 5003
rect 12378 4921 12386 4955
rect 12420 4921 12430 4955
rect 12378 4873 12430 4921
rect 12460 4995 12529 5003
rect 12460 4961 12485 4995
rect 12519 4961 12529 4995
rect 12460 4919 12529 4961
rect 12559 4919 12625 5003
rect 12655 4919 12697 5003
rect 12727 4983 12793 5003
rect 12727 4949 12737 4983
rect 12771 4949 12793 4983
rect 12727 4919 12793 4949
rect 12823 4978 12882 5003
rect 12823 4944 12838 4978
rect 12872 4944 12882 4978
rect 12823 4919 12882 4944
rect 12912 4995 12966 5003
rect 12912 4961 12922 4995
rect 12956 4961 12966 4995
rect 12912 4919 12966 4961
rect 12996 4978 13050 5003
rect 12996 4944 13006 4978
rect 13040 4944 13050 4978
rect 12996 4919 13050 4944
rect 13080 4986 13132 5003
rect 13080 4952 13090 4986
rect 13124 4952 13132 4986
rect 13080 4919 13132 4952
rect 13186 4978 13238 5003
rect 13186 4944 13194 4978
rect 13228 4944 13238 4978
rect 13186 4919 13238 4944
rect 13268 4995 13322 5003
rect 13268 4961 13278 4995
rect 13312 4961 13322 4995
rect 13268 4919 13322 4961
rect 13352 4978 13406 5003
rect 13352 4944 13362 4978
rect 13396 4944 13406 4978
rect 13352 4919 13406 4944
rect 13436 4978 13490 5003
rect 13436 4944 13446 4978
rect 13480 4944 13490 4978
rect 13436 4919 13490 4944
rect 13520 4919 13580 5003
rect 13610 4991 13679 5003
rect 13610 4957 13635 4991
rect 13669 4957 13679 4991
rect 13610 4919 13679 4957
rect 12460 4873 12512 4919
rect 13627 4873 13679 4919
rect 13709 4955 13761 5003
rect 13709 4921 13719 4955
rect 13753 4921 13761 4955
rect 13709 4873 13761 4921
rect 14380 4949 14432 4997
rect 14380 4915 14388 4949
rect 14422 4915 14432 4949
rect 14380 4867 14432 4915
rect 14462 4989 14531 4997
rect 14462 4955 14487 4989
rect 14521 4955 14531 4989
rect 14462 4913 14531 4955
rect 14561 4913 14627 4997
rect 14657 4913 14699 4997
rect 14729 4977 14795 4997
rect 14729 4943 14739 4977
rect 14773 4943 14795 4977
rect 14729 4913 14795 4943
rect 14825 4972 14884 4997
rect 14825 4938 14840 4972
rect 14874 4938 14884 4972
rect 14825 4913 14884 4938
rect 14914 4989 14968 4997
rect 14914 4955 14924 4989
rect 14958 4955 14968 4989
rect 14914 4913 14968 4955
rect 14998 4972 15052 4997
rect 14998 4938 15008 4972
rect 15042 4938 15052 4972
rect 14998 4913 15052 4938
rect 15082 4980 15134 4997
rect 15082 4946 15092 4980
rect 15126 4946 15134 4980
rect 15082 4913 15134 4946
rect 15188 4972 15240 4997
rect 15188 4938 15196 4972
rect 15230 4938 15240 4972
rect 15188 4913 15240 4938
rect 15270 4989 15324 4997
rect 15270 4955 15280 4989
rect 15314 4955 15324 4989
rect 15270 4913 15324 4955
rect 15354 4972 15408 4997
rect 15354 4938 15364 4972
rect 15398 4938 15408 4972
rect 15354 4913 15408 4938
rect 15438 4972 15492 4997
rect 15438 4938 15448 4972
rect 15482 4938 15492 4972
rect 15438 4913 15492 4938
rect 15522 4913 15582 4997
rect 15612 4985 15681 4997
rect 15612 4951 15637 4985
rect 15671 4951 15681 4985
rect 15612 4913 15681 4951
rect 14462 4867 14514 4913
rect 15629 4867 15681 4913
rect 15711 4949 15763 4997
rect 15711 4915 15721 4949
rect 15755 4915 15763 4949
rect 15711 4867 15763 4915
rect 16402 4931 16454 4979
rect 16402 4897 16410 4931
rect 16444 4897 16454 4931
rect 16402 4849 16454 4897
rect 16484 4971 16553 4979
rect 16484 4937 16509 4971
rect 16543 4937 16553 4971
rect 16484 4895 16553 4937
rect 16583 4895 16649 4979
rect 16679 4895 16721 4979
rect 16751 4959 16817 4979
rect 16751 4925 16761 4959
rect 16795 4925 16817 4959
rect 16751 4895 16817 4925
rect 16847 4954 16906 4979
rect 16847 4920 16862 4954
rect 16896 4920 16906 4954
rect 16847 4895 16906 4920
rect 16936 4971 16990 4979
rect 16936 4937 16946 4971
rect 16980 4937 16990 4971
rect 16936 4895 16990 4937
rect 17020 4954 17074 4979
rect 17020 4920 17030 4954
rect 17064 4920 17074 4954
rect 17020 4895 17074 4920
rect 17104 4962 17156 4979
rect 17104 4928 17114 4962
rect 17148 4928 17156 4962
rect 17104 4895 17156 4928
rect 17210 4954 17262 4979
rect 17210 4920 17218 4954
rect 17252 4920 17262 4954
rect 17210 4895 17262 4920
rect 17292 4971 17346 4979
rect 17292 4937 17302 4971
rect 17336 4937 17346 4971
rect 17292 4895 17346 4937
rect 17376 4954 17430 4979
rect 17376 4920 17386 4954
rect 17420 4920 17430 4954
rect 17376 4895 17430 4920
rect 17460 4954 17514 4979
rect 17460 4920 17470 4954
rect 17504 4920 17514 4954
rect 17460 4895 17514 4920
rect 17544 4895 17604 4979
rect 17634 4967 17703 4979
rect 17634 4933 17659 4967
rect 17693 4933 17703 4967
rect 17634 4895 17703 4933
rect 16484 4849 16536 4895
rect 17651 4849 17703 4895
rect 17733 4931 17785 4979
rect 17733 4897 17743 4931
rect 17777 4897 17785 4931
rect 17733 4849 17785 4897
rect 1868 2193 1920 2241
rect 1868 2159 1876 2193
rect 1910 2159 1920 2193
rect 1868 2111 1920 2159
rect 1950 2233 2019 2241
rect 1950 2199 1975 2233
rect 2009 2199 2019 2233
rect 1950 2157 2019 2199
rect 2049 2157 2115 2241
rect 2145 2157 2187 2241
rect 2217 2221 2283 2241
rect 2217 2187 2227 2221
rect 2261 2187 2283 2221
rect 2217 2157 2283 2187
rect 2313 2216 2372 2241
rect 2313 2182 2328 2216
rect 2362 2182 2372 2216
rect 2313 2157 2372 2182
rect 2402 2233 2456 2241
rect 2402 2199 2412 2233
rect 2446 2199 2456 2233
rect 2402 2157 2456 2199
rect 2486 2216 2540 2241
rect 2486 2182 2496 2216
rect 2530 2182 2540 2216
rect 2486 2157 2540 2182
rect 2570 2224 2622 2241
rect 2570 2190 2580 2224
rect 2614 2190 2622 2224
rect 2570 2157 2622 2190
rect 2676 2216 2728 2241
rect 2676 2182 2684 2216
rect 2718 2182 2728 2216
rect 2676 2157 2728 2182
rect 2758 2233 2812 2241
rect 2758 2199 2768 2233
rect 2802 2199 2812 2233
rect 2758 2157 2812 2199
rect 2842 2216 2896 2241
rect 2842 2182 2852 2216
rect 2886 2182 2896 2216
rect 2842 2157 2896 2182
rect 2926 2216 2980 2241
rect 2926 2182 2936 2216
rect 2970 2182 2980 2216
rect 2926 2157 2980 2182
rect 3010 2157 3070 2241
rect 3100 2229 3169 2241
rect 3100 2195 3125 2229
rect 3159 2195 3169 2229
rect 3100 2157 3169 2195
rect 1950 2111 2002 2157
rect 3117 2111 3169 2157
rect 3199 2193 3251 2241
rect 3199 2159 3209 2193
rect 3243 2159 3251 2193
rect 3199 2111 3251 2159
rect 3938 2189 3990 2237
rect 3938 2155 3946 2189
rect 3980 2155 3990 2189
rect 3938 2107 3990 2155
rect 4020 2229 4089 2237
rect 4020 2195 4045 2229
rect 4079 2195 4089 2229
rect 4020 2153 4089 2195
rect 4119 2153 4185 2237
rect 4215 2153 4257 2237
rect 4287 2217 4353 2237
rect 4287 2183 4297 2217
rect 4331 2183 4353 2217
rect 4287 2153 4353 2183
rect 4383 2212 4442 2237
rect 4383 2178 4398 2212
rect 4432 2178 4442 2212
rect 4383 2153 4442 2178
rect 4472 2229 4526 2237
rect 4472 2195 4482 2229
rect 4516 2195 4526 2229
rect 4472 2153 4526 2195
rect 4556 2212 4610 2237
rect 4556 2178 4566 2212
rect 4600 2178 4610 2212
rect 4556 2153 4610 2178
rect 4640 2220 4692 2237
rect 4640 2186 4650 2220
rect 4684 2186 4692 2220
rect 4640 2153 4692 2186
rect 4746 2212 4798 2237
rect 4746 2178 4754 2212
rect 4788 2178 4798 2212
rect 4746 2153 4798 2178
rect 4828 2229 4882 2237
rect 4828 2195 4838 2229
rect 4872 2195 4882 2229
rect 4828 2153 4882 2195
rect 4912 2212 4966 2237
rect 4912 2178 4922 2212
rect 4956 2178 4966 2212
rect 4912 2153 4966 2178
rect 4996 2212 5050 2237
rect 4996 2178 5006 2212
rect 5040 2178 5050 2212
rect 4996 2153 5050 2178
rect 5080 2153 5140 2237
rect 5170 2225 5239 2237
rect 5170 2191 5195 2225
rect 5229 2191 5239 2225
rect 5170 2153 5239 2191
rect 4020 2107 4072 2153
rect 5187 2107 5239 2153
rect 5269 2189 5321 2237
rect 5269 2155 5279 2189
rect 5313 2155 5321 2189
rect 5269 2107 5321 2155
rect 5890 2189 5942 2237
rect 5890 2155 5898 2189
rect 5932 2155 5942 2189
rect 5890 2107 5942 2155
rect 5972 2229 6041 2237
rect 5972 2195 5997 2229
rect 6031 2195 6041 2229
rect 5972 2153 6041 2195
rect 6071 2153 6137 2237
rect 6167 2153 6209 2237
rect 6239 2217 6305 2237
rect 6239 2183 6249 2217
rect 6283 2183 6305 2217
rect 6239 2153 6305 2183
rect 6335 2212 6394 2237
rect 6335 2178 6350 2212
rect 6384 2178 6394 2212
rect 6335 2153 6394 2178
rect 6424 2229 6478 2237
rect 6424 2195 6434 2229
rect 6468 2195 6478 2229
rect 6424 2153 6478 2195
rect 6508 2212 6562 2237
rect 6508 2178 6518 2212
rect 6552 2178 6562 2212
rect 6508 2153 6562 2178
rect 6592 2220 6644 2237
rect 6592 2186 6602 2220
rect 6636 2186 6644 2220
rect 6592 2153 6644 2186
rect 6698 2212 6750 2237
rect 6698 2178 6706 2212
rect 6740 2178 6750 2212
rect 6698 2153 6750 2178
rect 6780 2229 6834 2237
rect 6780 2195 6790 2229
rect 6824 2195 6834 2229
rect 6780 2153 6834 2195
rect 6864 2212 6918 2237
rect 6864 2178 6874 2212
rect 6908 2178 6918 2212
rect 6864 2153 6918 2178
rect 6948 2212 7002 2237
rect 6948 2178 6958 2212
rect 6992 2178 7002 2212
rect 6948 2153 7002 2178
rect 7032 2153 7092 2237
rect 7122 2225 7191 2237
rect 7122 2191 7147 2225
rect 7181 2191 7191 2225
rect 7122 2153 7191 2191
rect 5972 2107 6024 2153
rect 7139 2107 7191 2153
rect 7221 2189 7273 2237
rect 7221 2155 7231 2189
rect 7265 2155 7273 2189
rect 7221 2107 7273 2155
rect 7892 2195 7944 2243
rect 7892 2161 7900 2195
rect 7934 2161 7944 2195
rect 7892 2113 7944 2161
rect 7974 2235 8043 2243
rect 7974 2201 7999 2235
rect 8033 2201 8043 2235
rect 7974 2159 8043 2201
rect 8073 2159 8139 2243
rect 8169 2159 8211 2243
rect 8241 2223 8307 2243
rect 8241 2189 8251 2223
rect 8285 2189 8307 2223
rect 8241 2159 8307 2189
rect 8337 2218 8396 2243
rect 8337 2184 8352 2218
rect 8386 2184 8396 2218
rect 8337 2159 8396 2184
rect 8426 2235 8480 2243
rect 8426 2201 8436 2235
rect 8470 2201 8480 2235
rect 8426 2159 8480 2201
rect 8510 2218 8564 2243
rect 8510 2184 8520 2218
rect 8554 2184 8564 2218
rect 8510 2159 8564 2184
rect 8594 2226 8646 2243
rect 8594 2192 8604 2226
rect 8638 2192 8646 2226
rect 8594 2159 8646 2192
rect 8700 2218 8752 2243
rect 8700 2184 8708 2218
rect 8742 2184 8752 2218
rect 8700 2159 8752 2184
rect 8782 2235 8836 2243
rect 8782 2201 8792 2235
rect 8826 2201 8836 2235
rect 8782 2159 8836 2201
rect 8866 2218 8920 2243
rect 8866 2184 8876 2218
rect 8910 2184 8920 2218
rect 8866 2159 8920 2184
rect 8950 2218 9004 2243
rect 8950 2184 8960 2218
rect 8994 2184 9004 2218
rect 8950 2159 9004 2184
rect 9034 2159 9094 2243
rect 9124 2231 9193 2243
rect 9124 2197 9149 2231
rect 9183 2197 9193 2231
rect 9124 2159 9193 2197
rect 7974 2113 8026 2159
rect 9141 2113 9193 2159
rect 9223 2195 9275 2243
rect 9223 2161 9233 2195
rect 9267 2161 9275 2195
rect 9223 2113 9275 2161
rect 9844 2195 9896 2243
rect 9844 2161 9852 2195
rect 9886 2161 9896 2195
rect 9844 2113 9896 2161
rect 9926 2235 9995 2243
rect 9926 2201 9951 2235
rect 9985 2201 9995 2235
rect 9926 2159 9995 2201
rect 10025 2159 10091 2243
rect 10121 2159 10163 2243
rect 10193 2223 10259 2243
rect 10193 2189 10203 2223
rect 10237 2189 10259 2223
rect 10193 2159 10259 2189
rect 10289 2218 10348 2243
rect 10289 2184 10304 2218
rect 10338 2184 10348 2218
rect 10289 2159 10348 2184
rect 10378 2235 10432 2243
rect 10378 2201 10388 2235
rect 10422 2201 10432 2235
rect 10378 2159 10432 2201
rect 10462 2218 10516 2243
rect 10462 2184 10472 2218
rect 10506 2184 10516 2218
rect 10462 2159 10516 2184
rect 10546 2226 10598 2243
rect 10546 2192 10556 2226
rect 10590 2192 10598 2226
rect 10546 2159 10598 2192
rect 10652 2218 10704 2243
rect 10652 2184 10660 2218
rect 10694 2184 10704 2218
rect 10652 2159 10704 2184
rect 10734 2235 10788 2243
rect 10734 2201 10744 2235
rect 10778 2201 10788 2235
rect 10734 2159 10788 2201
rect 10818 2218 10872 2243
rect 10818 2184 10828 2218
rect 10862 2184 10872 2218
rect 10818 2159 10872 2184
rect 10902 2218 10956 2243
rect 10902 2184 10912 2218
rect 10946 2184 10956 2218
rect 10902 2159 10956 2184
rect 10986 2159 11046 2243
rect 11076 2231 11145 2243
rect 11076 2197 11101 2231
rect 11135 2197 11145 2231
rect 11076 2159 11145 2197
rect 9926 2113 9978 2159
rect 11093 2113 11145 2159
rect 11175 2195 11227 2243
rect 11175 2161 11185 2195
rect 11219 2161 11227 2195
rect 11175 2113 11227 2161
rect 11836 2195 11888 2243
rect 11836 2161 11844 2195
rect 11878 2161 11888 2195
rect 11836 2113 11888 2161
rect 11918 2235 11987 2243
rect 11918 2201 11943 2235
rect 11977 2201 11987 2235
rect 11918 2159 11987 2201
rect 12017 2159 12083 2243
rect 12113 2159 12155 2243
rect 12185 2223 12251 2243
rect 12185 2189 12195 2223
rect 12229 2189 12251 2223
rect 12185 2159 12251 2189
rect 12281 2218 12340 2243
rect 12281 2184 12296 2218
rect 12330 2184 12340 2218
rect 12281 2159 12340 2184
rect 12370 2235 12424 2243
rect 12370 2201 12380 2235
rect 12414 2201 12424 2235
rect 12370 2159 12424 2201
rect 12454 2218 12508 2243
rect 12454 2184 12464 2218
rect 12498 2184 12508 2218
rect 12454 2159 12508 2184
rect 12538 2226 12590 2243
rect 12538 2192 12548 2226
rect 12582 2192 12590 2226
rect 12538 2159 12590 2192
rect 12644 2218 12696 2243
rect 12644 2184 12652 2218
rect 12686 2184 12696 2218
rect 12644 2159 12696 2184
rect 12726 2235 12780 2243
rect 12726 2201 12736 2235
rect 12770 2201 12780 2235
rect 12726 2159 12780 2201
rect 12810 2218 12864 2243
rect 12810 2184 12820 2218
rect 12854 2184 12864 2218
rect 12810 2159 12864 2184
rect 12894 2218 12948 2243
rect 12894 2184 12904 2218
rect 12938 2184 12948 2218
rect 12894 2159 12948 2184
rect 12978 2159 13038 2243
rect 13068 2231 13137 2243
rect 13068 2197 13093 2231
rect 13127 2197 13137 2231
rect 13068 2159 13137 2197
rect 11918 2113 11970 2159
rect 13085 2113 13137 2159
rect 13167 2195 13219 2243
rect 13167 2161 13177 2195
rect 13211 2161 13219 2195
rect 13167 2113 13219 2161
rect 13788 2195 13840 2243
rect 13788 2161 13796 2195
rect 13830 2161 13840 2195
rect 13788 2113 13840 2161
rect 13870 2235 13939 2243
rect 13870 2201 13895 2235
rect 13929 2201 13939 2235
rect 13870 2159 13939 2201
rect 13969 2159 14035 2243
rect 14065 2159 14107 2243
rect 14137 2223 14203 2243
rect 14137 2189 14147 2223
rect 14181 2189 14203 2223
rect 14137 2159 14203 2189
rect 14233 2218 14292 2243
rect 14233 2184 14248 2218
rect 14282 2184 14292 2218
rect 14233 2159 14292 2184
rect 14322 2235 14376 2243
rect 14322 2201 14332 2235
rect 14366 2201 14376 2235
rect 14322 2159 14376 2201
rect 14406 2218 14460 2243
rect 14406 2184 14416 2218
rect 14450 2184 14460 2218
rect 14406 2159 14460 2184
rect 14490 2226 14542 2243
rect 14490 2192 14500 2226
rect 14534 2192 14542 2226
rect 14490 2159 14542 2192
rect 14596 2218 14648 2243
rect 14596 2184 14604 2218
rect 14638 2184 14648 2218
rect 14596 2159 14648 2184
rect 14678 2235 14732 2243
rect 14678 2201 14688 2235
rect 14722 2201 14732 2235
rect 14678 2159 14732 2201
rect 14762 2218 14816 2243
rect 14762 2184 14772 2218
rect 14806 2184 14816 2218
rect 14762 2159 14816 2184
rect 14846 2218 14900 2243
rect 14846 2184 14856 2218
rect 14890 2184 14900 2218
rect 14846 2159 14900 2184
rect 14930 2159 14990 2243
rect 15020 2231 15089 2243
rect 15020 2197 15045 2231
rect 15079 2197 15089 2231
rect 15020 2159 15089 2197
rect 13870 2113 13922 2159
rect 15037 2113 15089 2159
rect 15119 2195 15171 2243
rect 15119 2161 15129 2195
rect 15163 2161 15171 2195
rect 15119 2113 15171 2161
rect 15852 2195 15904 2243
rect 15852 2161 15860 2195
rect 15894 2161 15904 2195
rect 15852 2113 15904 2161
rect 15934 2235 16003 2243
rect 15934 2201 15959 2235
rect 15993 2201 16003 2235
rect 15934 2159 16003 2201
rect 16033 2159 16099 2243
rect 16129 2159 16171 2243
rect 16201 2223 16267 2243
rect 16201 2189 16211 2223
rect 16245 2189 16267 2223
rect 16201 2159 16267 2189
rect 16297 2218 16356 2243
rect 16297 2184 16312 2218
rect 16346 2184 16356 2218
rect 16297 2159 16356 2184
rect 16386 2235 16440 2243
rect 16386 2201 16396 2235
rect 16430 2201 16440 2235
rect 16386 2159 16440 2201
rect 16470 2218 16524 2243
rect 16470 2184 16480 2218
rect 16514 2184 16524 2218
rect 16470 2159 16524 2184
rect 16554 2226 16606 2243
rect 16554 2192 16564 2226
rect 16598 2192 16606 2226
rect 16554 2159 16606 2192
rect 16660 2218 16712 2243
rect 16660 2184 16668 2218
rect 16702 2184 16712 2218
rect 16660 2159 16712 2184
rect 16742 2235 16796 2243
rect 16742 2201 16752 2235
rect 16786 2201 16796 2235
rect 16742 2159 16796 2201
rect 16826 2218 16880 2243
rect 16826 2184 16836 2218
rect 16870 2184 16880 2218
rect 16826 2159 16880 2184
rect 16910 2218 16964 2243
rect 16910 2184 16920 2218
rect 16954 2184 16964 2218
rect 16910 2159 16964 2184
rect 16994 2159 17054 2243
rect 17084 2231 17153 2243
rect 17084 2197 17109 2231
rect 17143 2197 17153 2231
rect 17084 2159 17153 2197
rect 15934 2113 15986 2159
rect 17101 2113 17153 2159
rect 17183 2195 17235 2243
rect 17183 2161 17193 2195
rect 17227 2161 17235 2195
rect 17183 2113 17235 2161
<< pdiff >>
rect 9369 16531 9421 16543
rect 9369 16497 9377 16531
rect 9411 16497 9421 16531
rect 9369 16463 9421 16497
rect 9369 16429 9377 16463
rect 9411 16429 9421 16463
rect 9369 16343 9421 16429
rect 9451 16343 9505 16543
rect 9535 16521 9589 16543
rect 9535 16487 9545 16521
rect 9579 16487 9589 16521
rect 9535 16453 9589 16487
rect 9535 16419 9545 16453
rect 9579 16419 9589 16453
rect 9535 16343 9589 16419
rect 9619 16521 9673 16543
rect 9619 16487 9629 16521
rect 9663 16487 9673 16521
rect 9619 16453 9673 16487
rect 9619 16419 9629 16453
rect 9663 16419 9673 16453
rect 9619 16343 9673 16419
rect 9703 16521 9755 16543
rect 9703 16487 9713 16521
rect 9747 16487 9755 16521
rect 9703 16343 9755 16487
rect 9809 16521 9861 16543
rect 9809 16487 9817 16521
rect 9851 16487 9861 16521
rect 9809 16453 9861 16487
rect 9809 16419 9817 16453
rect 9851 16419 9861 16453
rect 9809 16343 9861 16419
rect 9891 16523 9951 16543
rect 9891 16489 9901 16523
rect 9935 16489 9951 16523
rect 9891 16455 9951 16489
rect 9891 16421 9901 16455
rect 9935 16421 9951 16455
rect 9891 16387 9951 16421
rect 9891 16353 9901 16387
rect 9935 16353 9951 16387
rect 9891 16343 9951 16353
rect 9687 15787 9739 15799
rect 9687 15757 9695 15787
rect 9491 15745 9547 15757
rect 9491 15711 9503 15745
rect 9537 15711 9547 15745
rect 9491 15673 9547 15711
rect 9577 15745 9631 15757
rect 9577 15711 9587 15745
rect 9621 15711 9631 15745
rect 9577 15673 9631 15711
rect 9661 15753 9695 15757
rect 9729 15753 9739 15787
rect 9661 15719 9739 15753
rect 9661 15685 9695 15719
rect 9729 15685 9739 15719
rect 9661 15673 9739 15685
rect 9677 15599 9739 15673
rect 9769 15787 9864 15799
rect 9769 15753 9799 15787
rect 9833 15753 9864 15787
rect 9769 15719 9864 15753
rect 9769 15685 9799 15719
rect 9833 15685 9864 15719
rect 9769 15599 9864 15685
rect 11501 15677 11553 15689
rect 11501 15643 11509 15677
rect 11543 15643 11553 15677
rect 11501 15605 11553 15643
rect 11583 15669 11653 15689
rect 11583 15635 11601 15669
rect 11635 15635 11653 15669
rect 11583 15605 11653 15635
rect 11683 15677 11757 15689
rect 11683 15643 11703 15677
rect 11737 15643 11757 15677
rect 11683 15605 11757 15643
rect 11787 15669 11843 15689
rect 11787 15635 11798 15669
rect 11832 15635 11843 15669
rect 11787 15605 11843 15635
rect 11873 15677 12009 15689
rect 11873 15643 11949 15677
rect 11983 15643 12009 15677
rect 11873 15609 12009 15643
rect 11873 15605 11949 15609
rect 11892 15575 11949 15605
rect 11983 15575 12009 15609
rect 11892 15489 12009 15575
rect 12039 15677 12091 15689
rect 12039 15643 12049 15677
rect 12083 15643 12091 15677
rect 12039 15609 12091 15643
rect 12039 15575 12049 15609
rect 12083 15575 12091 15609
rect 12039 15541 12091 15575
rect 12039 15507 12049 15541
rect 12083 15507 12091 15541
rect 12039 15489 12091 15507
rect 10871 15177 10923 15189
rect 10871 15147 10879 15177
rect 10675 15135 10731 15147
rect 10675 15101 10687 15135
rect 10721 15101 10731 15135
rect 10675 15063 10731 15101
rect 10761 15135 10815 15147
rect 10761 15101 10771 15135
rect 10805 15101 10815 15135
rect 10761 15063 10815 15101
rect 10845 15143 10879 15147
rect 10913 15143 10923 15177
rect 10845 15109 10923 15143
rect 10845 15075 10879 15109
rect 10913 15075 10923 15109
rect 10845 15063 10923 15075
rect 9379 14967 9431 14979
rect 9379 14933 9387 14967
rect 9421 14933 9431 14967
rect 9379 14899 9431 14933
rect 9379 14865 9387 14899
rect 9421 14865 9431 14899
rect 9379 14779 9431 14865
rect 9461 14779 9515 14979
rect 9545 14957 9599 14979
rect 9545 14923 9555 14957
rect 9589 14923 9599 14957
rect 9545 14889 9599 14923
rect 9545 14855 9555 14889
rect 9589 14855 9599 14889
rect 9545 14779 9599 14855
rect 9629 14957 9683 14979
rect 9629 14923 9639 14957
rect 9673 14923 9683 14957
rect 9629 14889 9683 14923
rect 9629 14855 9639 14889
rect 9673 14855 9683 14889
rect 9629 14779 9683 14855
rect 9713 14957 9765 14979
rect 9713 14923 9723 14957
rect 9757 14923 9765 14957
rect 9713 14779 9765 14923
rect 9819 14957 9871 14979
rect 9819 14923 9827 14957
rect 9861 14923 9871 14957
rect 9819 14889 9871 14923
rect 9819 14855 9827 14889
rect 9861 14855 9871 14889
rect 9819 14779 9871 14855
rect 9901 14959 9961 14979
rect 9901 14925 9911 14959
rect 9945 14925 9961 14959
rect 9901 14891 9961 14925
rect 9901 14857 9911 14891
rect 9945 14857 9961 14891
rect 9901 14823 9961 14857
rect 10861 14989 10923 15063
rect 10953 15177 11048 15189
rect 10953 15143 10983 15177
rect 11017 15143 11048 15177
rect 10953 15109 11048 15143
rect 10953 15075 10983 15109
rect 11017 15075 11048 15109
rect 10953 14989 11048 15075
rect 9901 14789 9911 14823
rect 9945 14789 9961 14823
rect 9901 14779 9961 14789
rect 9697 14223 9749 14235
rect 9697 14193 9705 14223
rect 9501 14181 9557 14193
rect 9501 14147 9513 14181
rect 9547 14147 9557 14181
rect 9501 14109 9557 14147
rect 9587 14181 9641 14193
rect 9587 14147 9597 14181
rect 9631 14147 9641 14181
rect 9587 14109 9641 14147
rect 9671 14189 9705 14193
rect 9739 14189 9749 14223
rect 9671 14155 9749 14189
rect 9671 14121 9705 14155
rect 9739 14121 9749 14155
rect 9671 14109 9749 14121
rect 9687 14035 9749 14109
rect 9779 14223 9874 14235
rect 9779 14189 9809 14223
rect 9843 14189 9874 14223
rect 9779 14155 9874 14189
rect 9779 14121 9809 14155
rect 9843 14121 9874 14155
rect 10717 14211 10769 14223
rect 10717 14177 10725 14211
rect 10759 14177 10769 14211
rect 10717 14139 10769 14177
rect 10799 14203 10869 14223
rect 10799 14169 10817 14203
rect 10851 14169 10869 14203
rect 10799 14139 10869 14169
rect 10899 14211 10973 14223
rect 10899 14177 10919 14211
rect 10953 14177 10973 14211
rect 10899 14139 10973 14177
rect 11003 14203 11059 14223
rect 11003 14169 11014 14203
rect 11048 14169 11059 14203
rect 11003 14139 11059 14169
rect 11089 14211 11225 14223
rect 11089 14177 11165 14211
rect 11199 14177 11225 14211
rect 11089 14143 11225 14177
rect 11089 14139 11165 14143
rect 9779 14035 9874 14121
rect 11108 14109 11165 14139
rect 11199 14109 11225 14143
rect 11108 14023 11225 14109
rect 11255 14211 11307 14223
rect 11255 14177 11265 14211
rect 11299 14177 11307 14211
rect 12976 14195 13029 14207
rect 11255 14143 11307 14177
rect 11255 14109 11265 14143
rect 11299 14109 11307 14143
rect 12976 14161 12984 14195
rect 13018 14161 13029 14195
rect 11255 14075 11307 14109
rect 12976 14127 13029 14161
rect 12976 14093 12984 14127
rect 13018 14093 13029 14127
rect 12976 14091 13029 14093
rect 11255 14041 11265 14075
rect 11299 14041 11307 14075
rect 11255 14023 11307 14041
rect 12615 14064 12667 14091
rect 12615 14030 12623 14064
rect 12657 14030 12667 14064
rect 12615 14007 12667 14030
rect 12697 14007 12763 14091
rect 12793 14007 12835 14091
rect 12865 14007 12931 14091
rect 12961 14007 13029 14091
rect 13059 14164 13113 14207
rect 13059 14130 13069 14164
rect 13103 14130 13113 14164
rect 13059 14096 13113 14130
rect 13059 14062 13069 14096
rect 13103 14062 13113 14096
rect 13059 14007 13113 14062
rect 11897 13821 11949 13849
rect 11897 13787 11905 13821
rect 11939 13787 11949 13821
rect 11897 13753 11949 13787
rect 11897 13733 11905 13753
rect 11728 13701 11780 13733
rect 11728 13667 11736 13701
rect 11770 13667 11780 13701
rect 11728 13649 11780 13667
rect 11810 13649 11852 13733
rect 11882 13719 11905 13733
rect 11939 13719 11949 13753
rect 11882 13649 11949 13719
rect 11979 13837 12047 13849
rect 11979 13803 12005 13837
rect 12039 13803 12047 13837
rect 11979 13769 12047 13803
rect 11979 13735 12005 13769
rect 12039 13735 12047 13769
rect 11979 13649 12047 13735
rect 9371 13299 9423 13311
rect 9371 13265 9379 13299
rect 9413 13265 9423 13299
rect 9371 13231 9423 13265
rect 9371 13197 9379 13231
rect 9413 13197 9423 13231
rect 9371 13111 9423 13197
rect 9453 13111 9507 13311
rect 9537 13289 9591 13311
rect 9537 13255 9547 13289
rect 9581 13255 9591 13289
rect 9537 13221 9591 13255
rect 9537 13187 9547 13221
rect 9581 13187 9591 13221
rect 9537 13111 9591 13187
rect 9621 13289 9675 13311
rect 9621 13255 9631 13289
rect 9665 13255 9675 13289
rect 9621 13221 9675 13255
rect 9621 13187 9631 13221
rect 9665 13187 9675 13221
rect 9621 13111 9675 13187
rect 9705 13289 9757 13311
rect 9705 13255 9715 13289
rect 9749 13255 9757 13289
rect 9705 13111 9757 13255
rect 9811 13289 9863 13311
rect 9811 13255 9819 13289
rect 9853 13255 9863 13289
rect 9811 13221 9863 13255
rect 9811 13187 9819 13221
rect 9853 13187 9863 13221
rect 9811 13111 9863 13187
rect 9893 13291 9953 13311
rect 11113 13369 11165 13381
rect 11113 13335 11121 13369
rect 11155 13335 11165 13369
rect 11113 13322 11165 13335
rect 9893 13257 9903 13291
rect 9937 13257 9953 13291
rect 11115 13268 11165 13322
rect 9893 13223 9953 13257
rect 9893 13189 9903 13223
rect 9937 13189 9953 13223
rect 9893 13155 9953 13189
rect 10841 13230 10893 13268
rect 10841 13196 10849 13230
rect 10883 13196 10893 13230
rect 10841 13184 10893 13196
rect 10923 13260 10977 13268
rect 10923 13226 10933 13260
rect 10967 13226 10977 13260
rect 10923 13184 10977 13226
rect 11007 13241 11070 13268
rect 11007 13207 11026 13241
rect 11060 13207 11070 13241
rect 11007 13184 11070 13207
rect 11100 13184 11165 13268
rect 9893 13121 9903 13155
rect 9937 13121 9953 13155
rect 9893 13111 9953 13121
rect 11115 13181 11165 13184
rect 11195 13355 11247 13381
rect 11195 13321 11205 13355
rect 11239 13321 11247 13355
rect 11195 13287 11247 13321
rect 11195 13253 11205 13287
rect 11239 13253 11247 13287
rect 11195 13181 11247 13253
rect 9689 12555 9741 12567
rect 9689 12525 9697 12555
rect 9493 12513 9549 12525
rect 9493 12479 9505 12513
rect 9539 12479 9549 12513
rect 9493 12441 9549 12479
rect 9579 12513 9633 12525
rect 9579 12479 9589 12513
rect 9623 12479 9633 12513
rect 9579 12441 9633 12479
rect 9663 12521 9697 12525
rect 9731 12521 9741 12555
rect 9663 12487 9741 12521
rect 9663 12453 9697 12487
rect 9731 12453 9741 12487
rect 9663 12441 9741 12453
rect 9679 12367 9741 12441
rect 9771 12555 9866 12567
rect 9771 12521 9801 12555
rect 9835 12521 9866 12555
rect 9771 12487 9866 12521
rect 9771 12453 9801 12487
rect 9835 12453 9866 12487
rect 9771 12367 9866 12453
rect 11065 12349 11117 12361
rect 11065 12319 11073 12349
rect 10869 12307 10925 12319
rect 10869 12273 10881 12307
rect 10915 12273 10925 12307
rect 10869 12235 10925 12273
rect 10955 12307 11009 12319
rect 10955 12273 10965 12307
rect 10999 12273 11009 12307
rect 10955 12235 11009 12273
rect 11039 12315 11073 12319
rect 11107 12315 11117 12349
rect 11039 12281 11117 12315
rect 11039 12247 11073 12281
rect 11107 12247 11117 12281
rect 11039 12235 11117 12247
rect 11055 12161 11117 12235
rect 11147 12349 11242 12361
rect 11147 12315 11177 12349
rect 11211 12315 11242 12349
rect 11147 12281 11242 12315
rect 11147 12247 11177 12281
rect 11211 12247 11242 12281
rect 11147 12161 11242 12247
rect 9381 11735 9433 11747
rect 9381 11701 9389 11735
rect 9423 11701 9433 11735
rect 9381 11667 9433 11701
rect 9381 11633 9389 11667
rect 9423 11633 9433 11667
rect 9381 11547 9433 11633
rect 9463 11547 9517 11747
rect 9547 11725 9601 11747
rect 9547 11691 9557 11725
rect 9591 11691 9601 11725
rect 9547 11657 9601 11691
rect 9547 11623 9557 11657
rect 9591 11623 9601 11657
rect 9547 11547 9601 11623
rect 9631 11725 9685 11747
rect 9631 11691 9641 11725
rect 9675 11691 9685 11725
rect 9631 11657 9685 11691
rect 9631 11623 9641 11657
rect 9675 11623 9685 11657
rect 9631 11547 9685 11623
rect 9715 11725 9767 11747
rect 9715 11691 9725 11725
rect 9759 11691 9767 11725
rect 9715 11547 9767 11691
rect 9821 11725 9873 11747
rect 9821 11691 9829 11725
rect 9863 11691 9873 11725
rect 9821 11657 9873 11691
rect 9821 11623 9829 11657
rect 9863 11623 9873 11657
rect 9821 11547 9873 11623
rect 9903 11727 9963 11747
rect 9903 11693 9913 11727
rect 9947 11693 9963 11727
rect 9903 11659 9963 11693
rect 9903 11625 9913 11659
rect 9947 11625 9963 11659
rect 9903 11591 9963 11625
rect 9903 11557 9913 11591
rect 9947 11557 9963 11591
rect 9903 11547 9963 11557
rect 9699 10991 9751 11003
rect 9699 10961 9707 10991
rect 9503 10949 9559 10961
rect 9503 10915 9515 10949
rect 9549 10915 9559 10949
rect 9503 10877 9559 10915
rect 9589 10949 9643 10961
rect 9589 10915 9599 10949
rect 9633 10915 9643 10949
rect 9589 10877 9643 10915
rect 9673 10957 9707 10961
rect 9741 10957 9751 10991
rect 9673 10923 9751 10957
rect 9673 10889 9707 10923
rect 9741 10889 9751 10923
rect 9673 10877 9751 10889
rect 9689 10803 9751 10877
rect 9781 10991 9876 11003
rect 9781 10957 9811 10991
rect 9845 10957 9876 10991
rect 9781 10923 9876 10957
rect 9781 10889 9811 10923
rect 9845 10889 9876 10923
rect 9781 10803 9876 10889
rect 6186 6285 6238 6303
rect 6186 6251 6194 6285
rect 6228 6251 6238 6285
rect 6186 6217 6238 6251
rect 6186 6183 6194 6217
rect 6228 6183 6238 6217
rect 6186 6149 6238 6183
rect 6186 6115 6194 6149
rect 6228 6115 6238 6149
rect 6186 6103 6238 6115
rect 6268 6285 6320 6303
rect 6268 6251 6278 6285
rect 6312 6251 6320 6285
rect 6268 6217 6320 6251
rect 6268 6183 6278 6217
rect 6312 6183 6320 6217
rect 6268 6149 6320 6183
rect 6268 6115 6278 6149
rect 6312 6115 6320 6149
rect 6268 6103 6320 6115
rect 10080 5633 10132 5671
rect 10080 5599 10088 5633
rect 10122 5599 10132 5633
rect 10080 5543 10132 5599
rect 1898 5213 1950 5251
rect 1898 5179 1906 5213
rect 1940 5179 1950 5213
rect 1898 5123 1950 5179
rect 1898 5089 1906 5123
rect 1940 5089 1950 5123
rect 1898 5051 1950 5089
rect 1980 5135 2032 5251
rect 10080 5509 10088 5543
rect 10122 5509 10132 5543
rect 3147 5135 3199 5251
rect 1980 5093 2049 5135
rect 1980 5059 1990 5093
rect 2024 5059 2049 5093
rect 1980 5051 2049 5059
rect 2079 5051 2145 5135
rect 2175 5051 2217 5135
rect 2247 5105 2313 5135
rect 2247 5071 2257 5105
rect 2291 5071 2313 5105
rect 2247 5051 2313 5071
rect 2343 5110 2402 5135
rect 2343 5076 2358 5110
rect 2392 5076 2402 5110
rect 2343 5051 2402 5076
rect 2432 5093 2486 5135
rect 2432 5059 2442 5093
rect 2476 5059 2486 5093
rect 2432 5051 2486 5059
rect 2516 5110 2570 5135
rect 2516 5076 2526 5110
rect 2560 5076 2570 5110
rect 2516 5051 2570 5076
rect 2600 5097 2652 5135
rect 2600 5063 2610 5097
rect 2644 5063 2652 5097
rect 2600 5051 2652 5063
rect 2706 5110 2758 5135
rect 2706 5076 2714 5110
rect 2748 5076 2758 5110
rect 2706 5051 2758 5076
rect 2788 5093 2842 5135
rect 2788 5059 2798 5093
rect 2832 5059 2842 5093
rect 2788 5051 2842 5059
rect 2872 5110 2926 5135
rect 2872 5076 2882 5110
rect 2916 5076 2926 5110
rect 2872 5051 2926 5076
rect 2956 5110 3010 5135
rect 2956 5076 2966 5110
rect 3000 5076 3010 5110
rect 2956 5051 3010 5076
rect 3040 5051 3100 5135
rect 3130 5101 3199 5135
rect 3130 5067 3155 5101
rect 3189 5067 3199 5101
rect 3130 5051 3199 5067
rect 3229 5210 3281 5251
rect 3229 5176 3239 5210
rect 3273 5176 3281 5210
rect 3229 5116 3281 5176
rect 3229 5082 3239 5116
rect 3273 5082 3281 5116
rect 3229 5051 3281 5082
rect 4032 5205 4084 5243
rect 4032 5171 4040 5205
rect 4074 5171 4084 5205
rect 4032 5115 4084 5171
rect 4032 5081 4040 5115
rect 4074 5081 4084 5115
rect 4032 5043 4084 5081
rect 4114 5127 4166 5243
rect 5281 5127 5333 5243
rect 4114 5085 4183 5127
rect 4114 5051 4124 5085
rect 4158 5051 4183 5085
rect 4114 5043 4183 5051
rect 4213 5043 4279 5127
rect 4309 5043 4351 5127
rect 4381 5097 4447 5127
rect 4381 5063 4391 5097
rect 4425 5063 4447 5097
rect 4381 5043 4447 5063
rect 4477 5102 4536 5127
rect 4477 5068 4492 5102
rect 4526 5068 4536 5102
rect 4477 5043 4536 5068
rect 4566 5085 4620 5127
rect 4566 5051 4576 5085
rect 4610 5051 4620 5085
rect 4566 5043 4620 5051
rect 4650 5102 4704 5127
rect 4650 5068 4660 5102
rect 4694 5068 4704 5102
rect 4650 5043 4704 5068
rect 4734 5089 4786 5127
rect 4734 5055 4744 5089
rect 4778 5055 4786 5089
rect 4734 5043 4786 5055
rect 4840 5102 4892 5127
rect 4840 5068 4848 5102
rect 4882 5068 4892 5102
rect 4840 5043 4892 5068
rect 4922 5085 4976 5127
rect 4922 5051 4932 5085
rect 4966 5051 4976 5085
rect 4922 5043 4976 5051
rect 5006 5102 5060 5127
rect 5006 5068 5016 5102
rect 5050 5068 5060 5102
rect 5006 5043 5060 5068
rect 5090 5102 5144 5127
rect 5090 5068 5100 5102
rect 5134 5068 5144 5102
rect 5090 5043 5144 5068
rect 5174 5043 5234 5127
rect 5264 5093 5333 5127
rect 5264 5059 5289 5093
rect 5323 5059 5333 5093
rect 5264 5043 5333 5059
rect 5363 5202 5415 5243
rect 5363 5168 5373 5202
rect 5407 5168 5415 5202
rect 5363 5108 5415 5168
rect 5363 5074 5373 5108
rect 5407 5074 5415 5108
rect 5363 5043 5415 5074
rect 5984 5205 6036 5243
rect 5984 5171 5992 5205
rect 6026 5171 6036 5205
rect 5984 5115 6036 5171
rect 5984 5081 5992 5115
rect 6026 5081 6036 5115
rect 5984 5043 6036 5081
rect 6066 5127 6118 5243
rect 7233 5127 7285 5243
rect 6066 5085 6135 5127
rect 6066 5051 6076 5085
rect 6110 5051 6135 5085
rect 6066 5043 6135 5051
rect 6165 5043 6231 5127
rect 6261 5043 6303 5127
rect 6333 5097 6399 5127
rect 6333 5063 6343 5097
rect 6377 5063 6399 5097
rect 6333 5043 6399 5063
rect 6429 5102 6488 5127
rect 6429 5068 6444 5102
rect 6478 5068 6488 5102
rect 6429 5043 6488 5068
rect 6518 5085 6572 5127
rect 6518 5051 6528 5085
rect 6562 5051 6572 5085
rect 6518 5043 6572 5051
rect 6602 5102 6656 5127
rect 6602 5068 6612 5102
rect 6646 5068 6656 5102
rect 6602 5043 6656 5068
rect 6686 5089 6738 5127
rect 6686 5055 6696 5089
rect 6730 5055 6738 5089
rect 6686 5043 6738 5055
rect 6792 5102 6844 5127
rect 6792 5068 6800 5102
rect 6834 5068 6844 5102
rect 6792 5043 6844 5068
rect 6874 5085 6928 5127
rect 6874 5051 6884 5085
rect 6918 5051 6928 5085
rect 6874 5043 6928 5051
rect 6958 5102 7012 5127
rect 6958 5068 6968 5102
rect 7002 5068 7012 5102
rect 6958 5043 7012 5068
rect 7042 5102 7096 5127
rect 7042 5068 7052 5102
rect 7086 5068 7096 5102
rect 7042 5043 7096 5068
rect 7126 5043 7186 5127
rect 7216 5093 7285 5127
rect 7216 5059 7241 5093
rect 7275 5059 7285 5093
rect 7216 5043 7285 5059
rect 7315 5202 7367 5243
rect 7315 5168 7325 5202
rect 7359 5168 7367 5202
rect 7315 5108 7367 5168
rect 7315 5074 7325 5108
rect 7359 5074 7367 5108
rect 7315 5043 7367 5074
rect 7986 5211 8038 5249
rect 7986 5177 7994 5211
rect 8028 5177 8038 5211
rect 7986 5121 8038 5177
rect 7986 5087 7994 5121
rect 8028 5087 8038 5121
rect 7986 5049 8038 5087
rect 8068 5133 8120 5249
rect 10080 5471 10132 5509
rect 10162 5555 10214 5671
rect 11329 5555 11381 5671
rect 10162 5513 10231 5555
rect 10162 5479 10172 5513
rect 10206 5479 10231 5513
rect 10162 5471 10231 5479
rect 10261 5471 10327 5555
rect 10357 5471 10399 5555
rect 10429 5525 10495 5555
rect 10429 5491 10439 5525
rect 10473 5491 10495 5525
rect 10429 5471 10495 5491
rect 10525 5530 10584 5555
rect 10525 5496 10540 5530
rect 10574 5496 10584 5530
rect 10525 5471 10584 5496
rect 10614 5513 10668 5555
rect 10614 5479 10624 5513
rect 10658 5479 10668 5513
rect 10614 5471 10668 5479
rect 10698 5530 10752 5555
rect 10698 5496 10708 5530
rect 10742 5496 10752 5530
rect 10698 5471 10752 5496
rect 10782 5517 10834 5555
rect 10782 5483 10792 5517
rect 10826 5483 10834 5517
rect 10782 5471 10834 5483
rect 10888 5530 10940 5555
rect 10888 5496 10896 5530
rect 10930 5496 10940 5530
rect 10888 5471 10940 5496
rect 10970 5513 11024 5555
rect 10970 5479 10980 5513
rect 11014 5479 11024 5513
rect 10970 5471 11024 5479
rect 11054 5530 11108 5555
rect 11054 5496 11064 5530
rect 11098 5496 11108 5530
rect 11054 5471 11108 5496
rect 11138 5530 11192 5555
rect 11138 5496 11148 5530
rect 11182 5496 11192 5530
rect 11138 5471 11192 5496
rect 11222 5471 11282 5555
rect 11312 5521 11381 5555
rect 11312 5487 11337 5521
rect 11371 5487 11381 5521
rect 11312 5471 11381 5487
rect 11411 5630 11463 5671
rect 11411 5596 11421 5630
rect 11455 5596 11463 5630
rect 11411 5536 11463 5596
rect 11411 5502 11421 5536
rect 11455 5502 11463 5536
rect 11411 5471 11463 5502
rect 12142 5621 12194 5659
rect 12142 5587 12150 5621
rect 12184 5587 12194 5621
rect 12142 5531 12194 5587
rect 12142 5497 12150 5531
rect 12184 5497 12194 5531
rect 12142 5459 12194 5497
rect 12224 5543 12276 5659
rect 13391 5543 13443 5659
rect 12224 5501 12293 5543
rect 12224 5467 12234 5501
rect 12268 5467 12293 5501
rect 12224 5459 12293 5467
rect 12323 5459 12389 5543
rect 12419 5459 12461 5543
rect 12491 5513 12557 5543
rect 12491 5479 12501 5513
rect 12535 5479 12557 5513
rect 12491 5459 12557 5479
rect 12587 5518 12646 5543
rect 12587 5484 12602 5518
rect 12636 5484 12646 5518
rect 12587 5459 12646 5484
rect 12676 5501 12730 5543
rect 12676 5467 12686 5501
rect 12720 5467 12730 5501
rect 12676 5459 12730 5467
rect 12760 5518 12814 5543
rect 12760 5484 12770 5518
rect 12804 5484 12814 5518
rect 12760 5459 12814 5484
rect 12844 5505 12896 5543
rect 12844 5471 12854 5505
rect 12888 5471 12896 5505
rect 12844 5459 12896 5471
rect 12950 5518 13002 5543
rect 12950 5484 12958 5518
rect 12992 5484 13002 5518
rect 12950 5459 13002 5484
rect 13032 5501 13086 5543
rect 13032 5467 13042 5501
rect 13076 5467 13086 5501
rect 13032 5459 13086 5467
rect 13116 5518 13170 5543
rect 13116 5484 13126 5518
rect 13160 5484 13170 5518
rect 13116 5459 13170 5484
rect 13200 5518 13254 5543
rect 13200 5484 13210 5518
rect 13244 5484 13254 5518
rect 13200 5459 13254 5484
rect 13284 5459 13344 5543
rect 13374 5509 13443 5543
rect 13374 5475 13399 5509
rect 13433 5475 13443 5509
rect 13374 5459 13443 5475
rect 13473 5618 13525 5659
rect 13473 5584 13483 5618
rect 13517 5584 13525 5618
rect 13473 5524 13525 5584
rect 13473 5490 13483 5524
rect 13517 5490 13525 5524
rect 13473 5459 13525 5490
rect 14100 5629 14152 5667
rect 14100 5595 14108 5629
rect 14142 5595 14152 5629
rect 14100 5539 14152 5595
rect 14100 5505 14108 5539
rect 14142 5505 14152 5539
rect 14100 5467 14152 5505
rect 14182 5551 14234 5667
rect 15349 5551 15401 5667
rect 14182 5509 14251 5551
rect 14182 5475 14192 5509
rect 14226 5475 14251 5509
rect 14182 5467 14251 5475
rect 14281 5467 14347 5551
rect 14377 5467 14419 5551
rect 14449 5521 14515 5551
rect 14449 5487 14459 5521
rect 14493 5487 14515 5521
rect 14449 5467 14515 5487
rect 14545 5526 14604 5551
rect 14545 5492 14560 5526
rect 14594 5492 14604 5526
rect 14545 5467 14604 5492
rect 14634 5509 14688 5551
rect 14634 5475 14644 5509
rect 14678 5475 14688 5509
rect 14634 5467 14688 5475
rect 14718 5526 14772 5551
rect 14718 5492 14728 5526
rect 14762 5492 14772 5526
rect 14718 5467 14772 5492
rect 14802 5513 14854 5551
rect 14802 5479 14812 5513
rect 14846 5479 14854 5513
rect 14802 5467 14854 5479
rect 14908 5526 14960 5551
rect 14908 5492 14916 5526
rect 14950 5492 14960 5526
rect 14908 5467 14960 5492
rect 14990 5509 15044 5551
rect 14990 5475 15000 5509
rect 15034 5475 15044 5509
rect 14990 5467 15044 5475
rect 15074 5526 15128 5551
rect 15074 5492 15084 5526
rect 15118 5492 15128 5526
rect 15074 5467 15128 5492
rect 15158 5526 15212 5551
rect 15158 5492 15168 5526
rect 15202 5492 15212 5526
rect 15158 5467 15212 5492
rect 15242 5467 15302 5551
rect 15332 5517 15401 5551
rect 15332 5483 15357 5517
rect 15391 5483 15401 5517
rect 15332 5467 15401 5483
rect 15431 5626 15483 5667
rect 15431 5592 15441 5626
rect 15475 5592 15483 5626
rect 15431 5532 15483 5592
rect 15431 5498 15441 5532
rect 15475 5498 15483 5532
rect 15431 5467 15483 5498
rect 16094 5635 16146 5673
rect 16094 5601 16102 5635
rect 16136 5601 16146 5635
rect 16094 5545 16146 5601
rect 16094 5511 16102 5545
rect 16136 5511 16146 5545
rect 16094 5473 16146 5511
rect 16176 5557 16228 5673
rect 17343 5557 17395 5673
rect 16176 5515 16245 5557
rect 16176 5481 16186 5515
rect 16220 5481 16245 5515
rect 16176 5473 16245 5481
rect 16275 5473 16341 5557
rect 16371 5473 16413 5557
rect 16443 5527 16509 5557
rect 16443 5493 16453 5527
rect 16487 5493 16509 5527
rect 16443 5473 16509 5493
rect 16539 5532 16598 5557
rect 16539 5498 16554 5532
rect 16588 5498 16598 5532
rect 16539 5473 16598 5498
rect 16628 5515 16682 5557
rect 16628 5481 16638 5515
rect 16672 5481 16682 5515
rect 16628 5473 16682 5481
rect 16712 5532 16766 5557
rect 16712 5498 16722 5532
rect 16756 5498 16766 5532
rect 16712 5473 16766 5498
rect 16796 5519 16848 5557
rect 16796 5485 16806 5519
rect 16840 5485 16848 5519
rect 16796 5473 16848 5485
rect 16902 5532 16954 5557
rect 16902 5498 16910 5532
rect 16944 5498 16954 5532
rect 16902 5473 16954 5498
rect 16984 5515 17038 5557
rect 16984 5481 16994 5515
rect 17028 5481 17038 5515
rect 16984 5473 17038 5481
rect 17068 5532 17122 5557
rect 17068 5498 17078 5532
rect 17112 5498 17122 5532
rect 17068 5473 17122 5498
rect 17152 5532 17206 5557
rect 17152 5498 17162 5532
rect 17196 5498 17206 5532
rect 17152 5473 17206 5498
rect 17236 5473 17296 5557
rect 17326 5523 17395 5557
rect 17326 5489 17351 5523
rect 17385 5489 17395 5523
rect 17326 5473 17395 5489
rect 17425 5632 17477 5673
rect 17425 5598 17435 5632
rect 17469 5598 17477 5632
rect 17425 5538 17477 5598
rect 17425 5504 17435 5538
rect 17469 5504 17477 5538
rect 17425 5473 17477 5504
rect 9235 5133 9287 5249
rect 8068 5091 8137 5133
rect 8068 5057 8078 5091
rect 8112 5057 8137 5091
rect 8068 5049 8137 5057
rect 8167 5049 8233 5133
rect 8263 5049 8305 5133
rect 8335 5103 8401 5133
rect 8335 5069 8345 5103
rect 8379 5069 8401 5103
rect 8335 5049 8401 5069
rect 8431 5108 8490 5133
rect 8431 5074 8446 5108
rect 8480 5074 8490 5108
rect 8431 5049 8490 5074
rect 8520 5091 8574 5133
rect 8520 5057 8530 5091
rect 8564 5057 8574 5091
rect 8520 5049 8574 5057
rect 8604 5108 8658 5133
rect 8604 5074 8614 5108
rect 8648 5074 8658 5108
rect 8604 5049 8658 5074
rect 8688 5095 8740 5133
rect 8688 5061 8698 5095
rect 8732 5061 8740 5095
rect 8688 5049 8740 5061
rect 8794 5108 8846 5133
rect 8794 5074 8802 5108
rect 8836 5074 8846 5108
rect 8794 5049 8846 5074
rect 8876 5091 8930 5133
rect 8876 5057 8886 5091
rect 8920 5057 8930 5091
rect 8876 5049 8930 5057
rect 8960 5108 9014 5133
rect 8960 5074 8970 5108
rect 9004 5074 9014 5108
rect 8960 5049 9014 5074
rect 9044 5108 9098 5133
rect 9044 5074 9054 5108
rect 9088 5074 9098 5108
rect 9044 5049 9098 5074
rect 9128 5049 9188 5133
rect 9218 5099 9287 5133
rect 9218 5065 9243 5099
rect 9277 5065 9287 5099
rect 9218 5049 9287 5065
rect 9317 5208 9369 5249
rect 9317 5174 9327 5208
rect 9361 5174 9369 5208
rect 9317 5114 9369 5174
rect 9317 5080 9327 5114
rect 9361 5080 9369 5114
rect 9317 5049 9369 5080
rect 10108 4759 10160 4797
rect 10108 4725 10116 4759
rect 10150 4725 10160 4759
rect 10108 4669 10160 4725
rect 10108 4635 10116 4669
rect 10150 4635 10160 4669
rect 10108 4597 10160 4635
rect 10190 4681 10242 4797
rect 11357 4681 11409 4797
rect 10190 4639 10259 4681
rect 10190 4605 10200 4639
rect 10234 4605 10259 4639
rect 10190 4597 10259 4605
rect 10289 4597 10355 4681
rect 10385 4597 10427 4681
rect 10457 4651 10523 4681
rect 10457 4617 10467 4651
rect 10501 4617 10523 4651
rect 10457 4597 10523 4617
rect 10553 4656 10612 4681
rect 10553 4622 10568 4656
rect 10602 4622 10612 4656
rect 10553 4597 10612 4622
rect 10642 4639 10696 4681
rect 10642 4605 10652 4639
rect 10686 4605 10696 4639
rect 10642 4597 10696 4605
rect 10726 4656 10780 4681
rect 10726 4622 10736 4656
rect 10770 4622 10780 4656
rect 10726 4597 10780 4622
rect 10810 4643 10862 4681
rect 10810 4609 10820 4643
rect 10854 4609 10862 4643
rect 10810 4597 10862 4609
rect 10916 4656 10968 4681
rect 10916 4622 10924 4656
rect 10958 4622 10968 4656
rect 10916 4597 10968 4622
rect 10998 4639 11052 4681
rect 10998 4605 11008 4639
rect 11042 4605 11052 4639
rect 10998 4597 11052 4605
rect 11082 4656 11136 4681
rect 11082 4622 11092 4656
rect 11126 4622 11136 4656
rect 11082 4597 11136 4622
rect 11166 4656 11220 4681
rect 11166 4622 11176 4656
rect 11210 4622 11220 4656
rect 11166 4597 11220 4622
rect 11250 4597 11310 4681
rect 11340 4647 11409 4681
rect 11340 4613 11365 4647
rect 11399 4613 11409 4647
rect 11340 4597 11409 4613
rect 11439 4756 11491 4797
rect 11439 4722 11449 4756
rect 11483 4722 11491 4756
rect 11439 4662 11491 4722
rect 11439 4628 11449 4662
rect 11483 4628 11491 4662
rect 11439 4597 11491 4628
rect 12378 4715 12430 4753
rect 12378 4681 12386 4715
rect 12420 4681 12430 4715
rect 12378 4625 12430 4681
rect 12378 4591 12386 4625
rect 12420 4591 12430 4625
rect 12378 4553 12430 4591
rect 12460 4637 12512 4753
rect 13627 4637 13679 4753
rect 12460 4595 12529 4637
rect 12460 4561 12470 4595
rect 12504 4561 12529 4595
rect 12460 4553 12529 4561
rect 12559 4553 12625 4637
rect 12655 4553 12697 4637
rect 12727 4607 12793 4637
rect 12727 4573 12737 4607
rect 12771 4573 12793 4607
rect 12727 4553 12793 4573
rect 12823 4612 12882 4637
rect 12823 4578 12838 4612
rect 12872 4578 12882 4612
rect 12823 4553 12882 4578
rect 12912 4595 12966 4637
rect 12912 4561 12922 4595
rect 12956 4561 12966 4595
rect 12912 4553 12966 4561
rect 12996 4612 13050 4637
rect 12996 4578 13006 4612
rect 13040 4578 13050 4612
rect 12996 4553 13050 4578
rect 13080 4599 13132 4637
rect 13080 4565 13090 4599
rect 13124 4565 13132 4599
rect 13080 4553 13132 4565
rect 13186 4612 13238 4637
rect 13186 4578 13194 4612
rect 13228 4578 13238 4612
rect 13186 4553 13238 4578
rect 13268 4595 13322 4637
rect 13268 4561 13278 4595
rect 13312 4561 13322 4595
rect 13268 4553 13322 4561
rect 13352 4612 13406 4637
rect 13352 4578 13362 4612
rect 13396 4578 13406 4612
rect 13352 4553 13406 4578
rect 13436 4612 13490 4637
rect 13436 4578 13446 4612
rect 13480 4578 13490 4612
rect 13436 4553 13490 4578
rect 13520 4553 13580 4637
rect 13610 4603 13679 4637
rect 13610 4569 13635 4603
rect 13669 4569 13679 4603
rect 13610 4553 13679 4569
rect 13709 4712 13761 4753
rect 13709 4678 13719 4712
rect 13753 4678 13761 4712
rect 13709 4618 13761 4678
rect 13709 4584 13719 4618
rect 13753 4584 13761 4618
rect 13709 4553 13761 4584
rect 14380 4709 14432 4747
rect 14380 4675 14388 4709
rect 14422 4675 14432 4709
rect 14380 4619 14432 4675
rect 14380 4585 14388 4619
rect 14422 4585 14432 4619
rect 14380 4547 14432 4585
rect 14462 4631 14514 4747
rect 15629 4631 15681 4747
rect 14462 4589 14531 4631
rect 14462 4555 14472 4589
rect 14506 4555 14531 4589
rect 14462 4547 14531 4555
rect 14561 4547 14627 4631
rect 14657 4547 14699 4631
rect 14729 4601 14795 4631
rect 14729 4567 14739 4601
rect 14773 4567 14795 4601
rect 14729 4547 14795 4567
rect 14825 4606 14884 4631
rect 14825 4572 14840 4606
rect 14874 4572 14884 4606
rect 14825 4547 14884 4572
rect 14914 4589 14968 4631
rect 14914 4555 14924 4589
rect 14958 4555 14968 4589
rect 14914 4547 14968 4555
rect 14998 4606 15052 4631
rect 14998 4572 15008 4606
rect 15042 4572 15052 4606
rect 14998 4547 15052 4572
rect 15082 4593 15134 4631
rect 15082 4559 15092 4593
rect 15126 4559 15134 4593
rect 15082 4547 15134 4559
rect 15188 4606 15240 4631
rect 15188 4572 15196 4606
rect 15230 4572 15240 4606
rect 15188 4547 15240 4572
rect 15270 4589 15324 4631
rect 15270 4555 15280 4589
rect 15314 4555 15324 4589
rect 15270 4547 15324 4555
rect 15354 4606 15408 4631
rect 15354 4572 15364 4606
rect 15398 4572 15408 4606
rect 15354 4547 15408 4572
rect 15438 4606 15492 4631
rect 15438 4572 15448 4606
rect 15482 4572 15492 4606
rect 15438 4547 15492 4572
rect 15522 4547 15582 4631
rect 15612 4597 15681 4631
rect 15612 4563 15637 4597
rect 15671 4563 15681 4597
rect 15612 4547 15681 4563
rect 15711 4706 15763 4747
rect 15711 4672 15721 4706
rect 15755 4672 15763 4706
rect 15711 4612 15763 4672
rect 15711 4578 15721 4612
rect 15755 4578 15763 4612
rect 15711 4547 15763 4578
rect 16402 4691 16454 4729
rect 16402 4657 16410 4691
rect 16444 4657 16454 4691
rect 16402 4601 16454 4657
rect 16402 4567 16410 4601
rect 16444 4567 16454 4601
rect 16402 4529 16454 4567
rect 16484 4613 16536 4729
rect 17651 4613 17703 4729
rect 16484 4571 16553 4613
rect 16484 4537 16494 4571
rect 16528 4537 16553 4571
rect 16484 4529 16553 4537
rect 16583 4529 16649 4613
rect 16679 4529 16721 4613
rect 16751 4583 16817 4613
rect 16751 4549 16761 4583
rect 16795 4549 16817 4583
rect 16751 4529 16817 4549
rect 16847 4588 16906 4613
rect 16847 4554 16862 4588
rect 16896 4554 16906 4588
rect 16847 4529 16906 4554
rect 16936 4571 16990 4613
rect 16936 4537 16946 4571
rect 16980 4537 16990 4571
rect 16936 4529 16990 4537
rect 17020 4588 17074 4613
rect 17020 4554 17030 4588
rect 17064 4554 17074 4588
rect 17020 4529 17074 4554
rect 17104 4575 17156 4613
rect 17104 4541 17114 4575
rect 17148 4541 17156 4575
rect 17104 4529 17156 4541
rect 17210 4588 17262 4613
rect 17210 4554 17218 4588
rect 17252 4554 17262 4588
rect 17210 4529 17262 4554
rect 17292 4571 17346 4613
rect 17292 4537 17302 4571
rect 17336 4537 17346 4571
rect 17292 4529 17346 4537
rect 17376 4588 17430 4613
rect 17376 4554 17386 4588
rect 17420 4554 17430 4588
rect 17376 4529 17430 4554
rect 17460 4588 17514 4613
rect 17460 4554 17470 4588
rect 17504 4554 17514 4588
rect 17460 4529 17514 4554
rect 17544 4529 17604 4613
rect 17634 4579 17703 4613
rect 17634 4545 17659 4579
rect 17693 4545 17703 4579
rect 17634 4529 17703 4545
rect 17733 4688 17785 4729
rect 17733 4654 17743 4688
rect 17777 4654 17785 4688
rect 17733 4594 17785 4654
rect 17733 4560 17743 4594
rect 17777 4560 17785 4594
rect 17733 4529 17785 4560
rect 1868 1953 1920 1991
rect 1868 1919 1876 1953
rect 1910 1919 1920 1953
rect 1868 1863 1920 1919
rect 1868 1829 1876 1863
rect 1910 1829 1920 1863
rect 1868 1791 1920 1829
rect 1950 1875 2002 1991
rect 3117 1875 3169 1991
rect 1950 1833 2019 1875
rect 1950 1799 1960 1833
rect 1994 1799 2019 1833
rect 1950 1791 2019 1799
rect 2049 1791 2115 1875
rect 2145 1791 2187 1875
rect 2217 1845 2283 1875
rect 2217 1811 2227 1845
rect 2261 1811 2283 1845
rect 2217 1791 2283 1811
rect 2313 1850 2372 1875
rect 2313 1816 2328 1850
rect 2362 1816 2372 1850
rect 2313 1791 2372 1816
rect 2402 1833 2456 1875
rect 2402 1799 2412 1833
rect 2446 1799 2456 1833
rect 2402 1791 2456 1799
rect 2486 1850 2540 1875
rect 2486 1816 2496 1850
rect 2530 1816 2540 1850
rect 2486 1791 2540 1816
rect 2570 1837 2622 1875
rect 2570 1803 2580 1837
rect 2614 1803 2622 1837
rect 2570 1791 2622 1803
rect 2676 1850 2728 1875
rect 2676 1816 2684 1850
rect 2718 1816 2728 1850
rect 2676 1791 2728 1816
rect 2758 1833 2812 1875
rect 2758 1799 2768 1833
rect 2802 1799 2812 1833
rect 2758 1791 2812 1799
rect 2842 1850 2896 1875
rect 2842 1816 2852 1850
rect 2886 1816 2896 1850
rect 2842 1791 2896 1816
rect 2926 1850 2980 1875
rect 2926 1816 2936 1850
rect 2970 1816 2980 1850
rect 2926 1791 2980 1816
rect 3010 1791 3070 1875
rect 3100 1841 3169 1875
rect 3100 1807 3125 1841
rect 3159 1807 3169 1841
rect 3100 1791 3169 1807
rect 3199 1950 3251 1991
rect 3199 1916 3209 1950
rect 3243 1916 3251 1950
rect 3199 1856 3251 1916
rect 3199 1822 3209 1856
rect 3243 1822 3251 1856
rect 3199 1791 3251 1822
rect 3938 1949 3990 1987
rect 3938 1915 3946 1949
rect 3980 1915 3990 1949
rect 3938 1859 3990 1915
rect 3938 1825 3946 1859
rect 3980 1825 3990 1859
rect 3938 1787 3990 1825
rect 4020 1871 4072 1987
rect 5187 1871 5239 1987
rect 4020 1829 4089 1871
rect 4020 1795 4030 1829
rect 4064 1795 4089 1829
rect 4020 1787 4089 1795
rect 4119 1787 4185 1871
rect 4215 1787 4257 1871
rect 4287 1841 4353 1871
rect 4287 1807 4297 1841
rect 4331 1807 4353 1841
rect 4287 1787 4353 1807
rect 4383 1846 4442 1871
rect 4383 1812 4398 1846
rect 4432 1812 4442 1846
rect 4383 1787 4442 1812
rect 4472 1829 4526 1871
rect 4472 1795 4482 1829
rect 4516 1795 4526 1829
rect 4472 1787 4526 1795
rect 4556 1846 4610 1871
rect 4556 1812 4566 1846
rect 4600 1812 4610 1846
rect 4556 1787 4610 1812
rect 4640 1833 4692 1871
rect 4640 1799 4650 1833
rect 4684 1799 4692 1833
rect 4640 1787 4692 1799
rect 4746 1846 4798 1871
rect 4746 1812 4754 1846
rect 4788 1812 4798 1846
rect 4746 1787 4798 1812
rect 4828 1829 4882 1871
rect 4828 1795 4838 1829
rect 4872 1795 4882 1829
rect 4828 1787 4882 1795
rect 4912 1846 4966 1871
rect 4912 1812 4922 1846
rect 4956 1812 4966 1846
rect 4912 1787 4966 1812
rect 4996 1846 5050 1871
rect 4996 1812 5006 1846
rect 5040 1812 5050 1846
rect 4996 1787 5050 1812
rect 5080 1787 5140 1871
rect 5170 1837 5239 1871
rect 5170 1803 5195 1837
rect 5229 1803 5239 1837
rect 5170 1787 5239 1803
rect 5269 1946 5321 1987
rect 5269 1912 5279 1946
rect 5313 1912 5321 1946
rect 5269 1852 5321 1912
rect 5269 1818 5279 1852
rect 5313 1818 5321 1852
rect 5269 1787 5321 1818
rect 5890 1949 5942 1987
rect 5890 1915 5898 1949
rect 5932 1915 5942 1949
rect 5890 1859 5942 1915
rect 5890 1825 5898 1859
rect 5932 1825 5942 1859
rect 5890 1787 5942 1825
rect 5972 1871 6024 1987
rect 7139 1871 7191 1987
rect 5972 1829 6041 1871
rect 5972 1795 5982 1829
rect 6016 1795 6041 1829
rect 5972 1787 6041 1795
rect 6071 1787 6137 1871
rect 6167 1787 6209 1871
rect 6239 1841 6305 1871
rect 6239 1807 6249 1841
rect 6283 1807 6305 1841
rect 6239 1787 6305 1807
rect 6335 1846 6394 1871
rect 6335 1812 6350 1846
rect 6384 1812 6394 1846
rect 6335 1787 6394 1812
rect 6424 1829 6478 1871
rect 6424 1795 6434 1829
rect 6468 1795 6478 1829
rect 6424 1787 6478 1795
rect 6508 1846 6562 1871
rect 6508 1812 6518 1846
rect 6552 1812 6562 1846
rect 6508 1787 6562 1812
rect 6592 1833 6644 1871
rect 6592 1799 6602 1833
rect 6636 1799 6644 1833
rect 6592 1787 6644 1799
rect 6698 1846 6750 1871
rect 6698 1812 6706 1846
rect 6740 1812 6750 1846
rect 6698 1787 6750 1812
rect 6780 1829 6834 1871
rect 6780 1795 6790 1829
rect 6824 1795 6834 1829
rect 6780 1787 6834 1795
rect 6864 1846 6918 1871
rect 6864 1812 6874 1846
rect 6908 1812 6918 1846
rect 6864 1787 6918 1812
rect 6948 1846 7002 1871
rect 6948 1812 6958 1846
rect 6992 1812 7002 1846
rect 6948 1787 7002 1812
rect 7032 1787 7092 1871
rect 7122 1837 7191 1871
rect 7122 1803 7147 1837
rect 7181 1803 7191 1837
rect 7122 1787 7191 1803
rect 7221 1946 7273 1987
rect 7221 1912 7231 1946
rect 7265 1912 7273 1946
rect 7221 1852 7273 1912
rect 7221 1818 7231 1852
rect 7265 1818 7273 1852
rect 7221 1787 7273 1818
rect 7892 1955 7944 1993
rect 7892 1921 7900 1955
rect 7934 1921 7944 1955
rect 7892 1865 7944 1921
rect 7892 1831 7900 1865
rect 7934 1831 7944 1865
rect 7892 1793 7944 1831
rect 7974 1877 8026 1993
rect 9141 1877 9193 1993
rect 7974 1835 8043 1877
rect 7974 1801 7984 1835
rect 8018 1801 8043 1835
rect 7974 1793 8043 1801
rect 8073 1793 8139 1877
rect 8169 1793 8211 1877
rect 8241 1847 8307 1877
rect 8241 1813 8251 1847
rect 8285 1813 8307 1847
rect 8241 1793 8307 1813
rect 8337 1852 8396 1877
rect 8337 1818 8352 1852
rect 8386 1818 8396 1852
rect 8337 1793 8396 1818
rect 8426 1835 8480 1877
rect 8426 1801 8436 1835
rect 8470 1801 8480 1835
rect 8426 1793 8480 1801
rect 8510 1852 8564 1877
rect 8510 1818 8520 1852
rect 8554 1818 8564 1852
rect 8510 1793 8564 1818
rect 8594 1839 8646 1877
rect 8594 1805 8604 1839
rect 8638 1805 8646 1839
rect 8594 1793 8646 1805
rect 8700 1852 8752 1877
rect 8700 1818 8708 1852
rect 8742 1818 8752 1852
rect 8700 1793 8752 1818
rect 8782 1835 8836 1877
rect 8782 1801 8792 1835
rect 8826 1801 8836 1835
rect 8782 1793 8836 1801
rect 8866 1852 8920 1877
rect 8866 1818 8876 1852
rect 8910 1818 8920 1852
rect 8866 1793 8920 1818
rect 8950 1852 9004 1877
rect 8950 1818 8960 1852
rect 8994 1818 9004 1852
rect 8950 1793 9004 1818
rect 9034 1793 9094 1877
rect 9124 1843 9193 1877
rect 9124 1809 9149 1843
rect 9183 1809 9193 1843
rect 9124 1793 9193 1809
rect 9223 1952 9275 1993
rect 9223 1918 9233 1952
rect 9267 1918 9275 1952
rect 9223 1858 9275 1918
rect 9223 1824 9233 1858
rect 9267 1824 9275 1858
rect 9223 1793 9275 1824
rect 9844 1955 9896 1993
rect 9844 1921 9852 1955
rect 9886 1921 9896 1955
rect 9844 1865 9896 1921
rect 9844 1831 9852 1865
rect 9886 1831 9896 1865
rect 9844 1793 9896 1831
rect 9926 1877 9978 1993
rect 11093 1877 11145 1993
rect 9926 1835 9995 1877
rect 9926 1801 9936 1835
rect 9970 1801 9995 1835
rect 9926 1793 9995 1801
rect 10025 1793 10091 1877
rect 10121 1793 10163 1877
rect 10193 1847 10259 1877
rect 10193 1813 10203 1847
rect 10237 1813 10259 1847
rect 10193 1793 10259 1813
rect 10289 1852 10348 1877
rect 10289 1818 10304 1852
rect 10338 1818 10348 1852
rect 10289 1793 10348 1818
rect 10378 1835 10432 1877
rect 10378 1801 10388 1835
rect 10422 1801 10432 1835
rect 10378 1793 10432 1801
rect 10462 1852 10516 1877
rect 10462 1818 10472 1852
rect 10506 1818 10516 1852
rect 10462 1793 10516 1818
rect 10546 1839 10598 1877
rect 10546 1805 10556 1839
rect 10590 1805 10598 1839
rect 10546 1793 10598 1805
rect 10652 1852 10704 1877
rect 10652 1818 10660 1852
rect 10694 1818 10704 1852
rect 10652 1793 10704 1818
rect 10734 1835 10788 1877
rect 10734 1801 10744 1835
rect 10778 1801 10788 1835
rect 10734 1793 10788 1801
rect 10818 1852 10872 1877
rect 10818 1818 10828 1852
rect 10862 1818 10872 1852
rect 10818 1793 10872 1818
rect 10902 1852 10956 1877
rect 10902 1818 10912 1852
rect 10946 1818 10956 1852
rect 10902 1793 10956 1818
rect 10986 1793 11046 1877
rect 11076 1843 11145 1877
rect 11076 1809 11101 1843
rect 11135 1809 11145 1843
rect 11076 1793 11145 1809
rect 11175 1952 11227 1993
rect 11175 1918 11185 1952
rect 11219 1918 11227 1952
rect 11175 1858 11227 1918
rect 11175 1824 11185 1858
rect 11219 1824 11227 1858
rect 11175 1793 11227 1824
rect 11836 1955 11888 1993
rect 11836 1921 11844 1955
rect 11878 1921 11888 1955
rect 11836 1865 11888 1921
rect 11836 1831 11844 1865
rect 11878 1831 11888 1865
rect 11836 1793 11888 1831
rect 11918 1877 11970 1993
rect 13085 1877 13137 1993
rect 11918 1835 11987 1877
rect 11918 1801 11928 1835
rect 11962 1801 11987 1835
rect 11918 1793 11987 1801
rect 12017 1793 12083 1877
rect 12113 1793 12155 1877
rect 12185 1847 12251 1877
rect 12185 1813 12195 1847
rect 12229 1813 12251 1847
rect 12185 1793 12251 1813
rect 12281 1852 12340 1877
rect 12281 1818 12296 1852
rect 12330 1818 12340 1852
rect 12281 1793 12340 1818
rect 12370 1835 12424 1877
rect 12370 1801 12380 1835
rect 12414 1801 12424 1835
rect 12370 1793 12424 1801
rect 12454 1852 12508 1877
rect 12454 1818 12464 1852
rect 12498 1818 12508 1852
rect 12454 1793 12508 1818
rect 12538 1839 12590 1877
rect 12538 1805 12548 1839
rect 12582 1805 12590 1839
rect 12538 1793 12590 1805
rect 12644 1852 12696 1877
rect 12644 1818 12652 1852
rect 12686 1818 12696 1852
rect 12644 1793 12696 1818
rect 12726 1835 12780 1877
rect 12726 1801 12736 1835
rect 12770 1801 12780 1835
rect 12726 1793 12780 1801
rect 12810 1852 12864 1877
rect 12810 1818 12820 1852
rect 12854 1818 12864 1852
rect 12810 1793 12864 1818
rect 12894 1852 12948 1877
rect 12894 1818 12904 1852
rect 12938 1818 12948 1852
rect 12894 1793 12948 1818
rect 12978 1793 13038 1877
rect 13068 1843 13137 1877
rect 13068 1809 13093 1843
rect 13127 1809 13137 1843
rect 13068 1793 13137 1809
rect 13167 1952 13219 1993
rect 13167 1918 13177 1952
rect 13211 1918 13219 1952
rect 13167 1858 13219 1918
rect 13167 1824 13177 1858
rect 13211 1824 13219 1858
rect 13167 1793 13219 1824
rect 13788 1955 13840 1993
rect 13788 1921 13796 1955
rect 13830 1921 13840 1955
rect 13788 1865 13840 1921
rect 13788 1831 13796 1865
rect 13830 1831 13840 1865
rect 13788 1793 13840 1831
rect 13870 1877 13922 1993
rect 15037 1877 15089 1993
rect 13870 1835 13939 1877
rect 13870 1801 13880 1835
rect 13914 1801 13939 1835
rect 13870 1793 13939 1801
rect 13969 1793 14035 1877
rect 14065 1793 14107 1877
rect 14137 1847 14203 1877
rect 14137 1813 14147 1847
rect 14181 1813 14203 1847
rect 14137 1793 14203 1813
rect 14233 1852 14292 1877
rect 14233 1818 14248 1852
rect 14282 1818 14292 1852
rect 14233 1793 14292 1818
rect 14322 1835 14376 1877
rect 14322 1801 14332 1835
rect 14366 1801 14376 1835
rect 14322 1793 14376 1801
rect 14406 1852 14460 1877
rect 14406 1818 14416 1852
rect 14450 1818 14460 1852
rect 14406 1793 14460 1818
rect 14490 1839 14542 1877
rect 14490 1805 14500 1839
rect 14534 1805 14542 1839
rect 14490 1793 14542 1805
rect 14596 1852 14648 1877
rect 14596 1818 14604 1852
rect 14638 1818 14648 1852
rect 14596 1793 14648 1818
rect 14678 1835 14732 1877
rect 14678 1801 14688 1835
rect 14722 1801 14732 1835
rect 14678 1793 14732 1801
rect 14762 1852 14816 1877
rect 14762 1818 14772 1852
rect 14806 1818 14816 1852
rect 14762 1793 14816 1818
rect 14846 1852 14900 1877
rect 14846 1818 14856 1852
rect 14890 1818 14900 1852
rect 14846 1793 14900 1818
rect 14930 1793 14990 1877
rect 15020 1843 15089 1877
rect 15020 1809 15045 1843
rect 15079 1809 15089 1843
rect 15020 1793 15089 1809
rect 15119 1952 15171 1993
rect 15119 1918 15129 1952
rect 15163 1918 15171 1952
rect 15119 1858 15171 1918
rect 15119 1824 15129 1858
rect 15163 1824 15171 1858
rect 15119 1793 15171 1824
rect 15852 1955 15904 1993
rect 15852 1921 15860 1955
rect 15894 1921 15904 1955
rect 15852 1865 15904 1921
rect 15852 1831 15860 1865
rect 15894 1831 15904 1865
rect 15852 1793 15904 1831
rect 15934 1877 15986 1993
rect 17101 1877 17153 1993
rect 15934 1835 16003 1877
rect 15934 1801 15944 1835
rect 15978 1801 16003 1835
rect 15934 1793 16003 1801
rect 16033 1793 16099 1877
rect 16129 1793 16171 1877
rect 16201 1847 16267 1877
rect 16201 1813 16211 1847
rect 16245 1813 16267 1847
rect 16201 1793 16267 1813
rect 16297 1852 16356 1877
rect 16297 1818 16312 1852
rect 16346 1818 16356 1852
rect 16297 1793 16356 1818
rect 16386 1835 16440 1877
rect 16386 1801 16396 1835
rect 16430 1801 16440 1835
rect 16386 1793 16440 1801
rect 16470 1852 16524 1877
rect 16470 1818 16480 1852
rect 16514 1818 16524 1852
rect 16470 1793 16524 1818
rect 16554 1839 16606 1877
rect 16554 1805 16564 1839
rect 16598 1805 16606 1839
rect 16554 1793 16606 1805
rect 16660 1852 16712 1877
rect 16660 1818 16668 1852
rect 16702 1818 16712 1852
rect 16660 1793 16712 1818
rect 16742 1835 16796 1877
rect 16742 1801 16752 1835
rect 16786 1801 16796 1835
rect 16742 1793 16796 1801
rect 16826 1852 16880 1877
rect 16826 1818 16836 1852
rect 16870 1818 16880 1852
rect 16826 1793 16880 1818
rect 16910 1852 16964 1877
rect 16910 1818 16920 1852
rect 16954 1818 16964 1852
rect 16910 1793 16964 1818
rect 16994 1793 17054 1877
rect 17084 1843 17153 1877
rect 17084 1809 17109 1843
rect 17143 1809 17153 1843
rect 17084 1793 17153 1809
rect 17183 1952 17235 1993
rect 17183 1918 17193 1952
rect 17227 1918 17235 1952
rect 17183 1858 17235 1918
rect 17183 1824 17193 1858
rect 17227 1824 17235 1858
rect 17183 1793 17235 1824
<< ndiffc >>
rect 9377 16107 9411 16141
rect 9461 16129 9495 16163
rect 9545 16107 9579 16141
rect 9713 16109 9747 16143
rect 9813 16109 9847 16143
rect 9903 16180 9937 16214
rect 9903 16112 9937 16146
rect 9503 15389 9537 15423
rect 9695 15361 9729 15395
rect 9779 15361 9813 15395
rect 11509 15259 11543 15293
rect 11950 15319 11984 15353
rect 11950 15251 11984 15285
rect 12049 15319 12083 15353
rect 12049 15251 12083 15285
rect 10687 14779 10721 14813
rect 10879 14751 10913 14785
rect 10963 14751 10997 14785
rect 9387 14543 9421 14577
rect 9471 14565 9505 14599
rect 9555 14543 9589 14577
rect 9723 14545 9757 14579
rect 9823 14545 9857 14579
rect 9913 14616 9947 14650
rect 9913 14548 9947 14582
rect 9513 13825 9547 13859
rect 9705 13797 9739 13831
rect 9789 13797 9823 13831
rect 10725 13793 10759 13827
rect 11166 13853 11200 13887
rect 11166 13785 11200 13819
rect 11265 13853 11299 13887
rect 11265 13785 11299 13819
rect 12623 13793 12657 13827
rect 12713 13787 12747 13821
rect 12803 13773 12837 13807
rect 12887 13787 12921 13821
rect 12981 13773 13015 13807
rect 13069 13811 13103 13845
rect 11724 13421 11758 13455
rect 11808 13421 11842 13455
rect 11904 13421 11938 13455
rect 11989 13481 12023 13515
rect 11989 13413 12023 13447
rect 9379 12875 9413 12909
rect 9463 12897 9497 12931
rect 9547 12875 9581 12909
rect 9715 12877 9749 12911
rect 9815 12877 9849 12911
rect 9905 12948 9939 12982
rect 10849 12943 10883 12977
rect 11121 12959 11155 12993
rect 11205 12969 11239 13003
rect 9905 12880 9939 12914
rect 9505 12157 9539 12191
rect 9697 12129 9731 12163
rect 9781 12129 9815 12163
rect 10881 11951 10915 11985
rect 11073 11923 11107 11957
rect 11157 11923 11191 11957
rect 9389 11311 9423 11345
rect 9473 11333 9507 11367
rect 9557 11311 9591 11345
rect 9725 11313 9759 11347
rect 9825 11313 9859 11347
rect 9915 11384 9949 11418
rect 9915 11316 9949 11350
rect 9515 10593 9549 10627
rect 9707 10565 9741 10599
rect 9791 10565 9825 10599
rect 6194 6503 6228 6537
rect 6194 6435 6228 6469
rect 6278 6503 6312 6537
rect 6278 6435 6312 6469
rect 10088 5839 10122 5873
rect 10187 5879 10221 5913
rect 10439 5867 10473 5901
rect 10540 5862 10574 5896
rect 10624 5879 10658 5913
rect 10708 5862 10742 5896
rect 10792 5870 10826 5904
rect 10896 5862 10930 5896
rect 10980 5879 11014 5913
rect 11064 5862 11098 5896
rect 11148 5862 11182 5896
rect 11337 5875 11371 5909
rect 1906 5419 1940 5453
rect 2005 5459 2039 5493
rect 2257 5447 2291 5481
rect 2358 5442 2392 5476
rect 2442 5459 2476 5493
rect 2526 5442 2560 5476
rect 2610 5450 2644 5484
rect 2714 5442 2748 5476
rect 2798 5459 2832 5493
rect 2882 5442 2916 5476
rect 2966 5442 3000 5476
rect 3155 5455 3189 5489
rect 3239 5419 3273 5453
rect 4040 5411 4074 5445
rect 4139 5451 4173 5485
rect 4391 5439 4425 5473
rect 4492 5434 4526 5468
rect 4576 5451 4610 5485
rect 4660 5434 4694 5468
rect 4744 5442 4778 5476
rect 4848 5434 4882 5468
rect 4932 5451 4966 5485
rect 5016 5434 5050 5468
rect 5100 5434 5134 5468
rect 5289 5447 5323 5481
rect 5373 5411 5407 5445
rect 5992 5411 6026 5445
rect 6091 5451 6125 5485
rect 6343 5439 6377 5473
rect 6444 5434 6478 5468
rect 6528 5451 6562 5485
rect 6612 5434 6646 5468
rect 6696 5442 6730 5476
rect 6800 5434 6834 5468
rect 6884 5451 6918 5485
rect 6968 5434 7002 5468
rect 7052 5434 7086 5468
rect 7241 5447 7275 5481
rect 7325 5411 7359 5445
rect 7994 5417 8028 5451
rect 8093 5457 8127 5491
rect 8345 5445 8379 5479
rect 8446 5440 8480 5474
rect 8530 5457 8564 5491
rect 8614 5440 8648 5474
rect 8698 5448 8732 5482
rect 8802 5440 8836 5474
rect 8886 5457 8920 5491
rect 8970 5440 9004 5474
rect 9054 5440 9088 5474
rect 9243 5453 9277 5487
rect 11421 5839 11455 5873
rect 12150 5827 12184 5861
rect 12249 5867 12283 5901
rect 12501 5855 12535 5889
rect 12602 5850 12636 5884
rect 12686 5867 12720 5901
rect 12770 5850 12804 5884
rect 12854 5858 12888 5892
rect 12958 5850 12992 5884
rect 13042 5867 13076 5901
rect 13126 5850 13160 5884
rect 13210 5850 13244 5884
rect 13399 5863 13433 5897
rect 9327 5417 9361 5451
rect 13483 5827 13517 5861
rect 14108 5835 14142 5869
rect 14207 5875 14241 5909
rect 14459 5863 14493 5897
rect 14560 5858 14594 5892
rect 14644 5875 14678 5909
rect 14728 5858 14762 5892
rect 14812 5866 14846 5900
rect 14916 5858 14950 5892
rect 15000 5875 15034 5909
rect 15084 5858 15118 5892
rect 15168 5858 15202 5892
rect 15357 5871 15391 5905
rect 15441 5835 15475 5869
rect 16102 5841 16136 5875
rect 16201 5881 16235 5915
rect 16453 5869 16487 5903
rect 16554 5864 16588 5898
rect 16638 5881 16672 5915
rect 16722 5864 16756 5898
rect 16806 5872 16840 5906
rect 16910 5864 16944 5898
rect 16994 5881 17028 5915
rect 17078 5864 17112 5898
rect 17162 5864 17196 5898
rect 17351 5877 17385 5911
rect 17435 5841 17469 5875
rect 10116 4965 10150 4999
rect 10215 5005 10249 5039
rect 10467 4993 10501 5027
rect 10568 4988 10602 5022
rect 10652 5005 10686 5039
rect 10736 4988 10770 5022
rect 10820 4996 10854 5030
rect 10924 4988 10958 5022
rect 11008 5005 11042 5039
rect 11092 4988 11126 5022
rect 11176 4988 11210 5022
rect 11365 5001 11399 5035
rect 11449 4965 11483 4999
rect 12386 4921 12420 4955
rect 12485 4961 12519 4995
rect 12737 4949 12771 4983
rect 12838 4944 12872 4978
rect 12922 4961 12956 4995
rect 13006 4944 13040 4978
rect 13090 4952 13124 4986
rect 13194 4944 13228 4978
rect 13278 4961 13312 4995
rect 13362 4944 13396 4978
rect 13446 4944 13480 4978
rect 13635 4957 13669 4991
rect 13719 4921 13753 4955
rect 14388 4915 14422 4949
rect 14487 4955 14521 4989
rect 14739 4943 14773 4977
rect 14840 4938 14874 4972
rect 14924 4955 14958 4989
rect 15008 4938 15042 4972
rect 15092 4946 15126 4980
rect 15196 4938 15230 4972
rect 15280 4955 15314 4989
rect 15364 4938 15398 4972
rect 15448 4938 15482 4972
rect 15637 4951 15671 4985
rect 15721 4915 15755 4949
rect 16410 4897 16444 4931
rect 16509 4937 16543 4971
rect 16761 4925 16795 4959
rect 16862 4920 16896 4954
rect 16946 4937 16980 4971
rect 17030 4920 17064 4954
rect 17114 4928 17148 4962
rect 17218 4920 17252 4954
rect 17302 4937 17336 4971
rect 17386 4920 17420 4954
rect 17470 4920 17504 4954
rect 17659 4933 17693 4967
rect 17743 4897 17777 4931
rect 1876 2159 1910 2193
rect 1975 2199 2009 2233
rect 2227 2187 2261 2221
rect 2328 2182 2362 2216
rect 2412 2199 2446 2233
rect 2496 2182 2530 2216
rect 2580 2190 2614 2224
rect 2684 2182 2718 2216
rect 2768 2199 2802 2233
rect 2852 2182 2886 2216
rect 2936 2182 2970 2216
rect 3125 2195 3159 2229
rect 3209 2159 3243 2193
rect 3946 2155 3980 2189
rect 4045 2195 4079 2229
rect 4297 2183 4331 2217
rect 4398 2178 4432 2212
rect 4482 2195 4516 2229
rect 4566 2178 4600 2212
rect 4650 2186 4684 2220
rect 4754 2178 4788 2212
rect 4838 2195 4872 2229
rect 4922 2178 4956 2212
rect 5006 2178 5040 2212
rect 5195 2191 5229 2225
rect 5279 2155 5313 2189
rect 5898 2155 5932 2189
rect 5997 2195 6031 2229
rect 6249 2183 6283 2217
rect 6350 2178 6384 2212
rect 6434 2195 6468 2229
rect 6518 2178 6552 2212
rect 6602 2186 6636 2220
rect 6706 2178 6740 2212
rect 6790 2195 6824 2229
rect 6874 2178 6908 2212
rect 6958 2178 6992 2212
rect 7147 2191 7181 2225
rect 7231 2155 7265 2189
rect 7900 2161 7934 2195
rect 7999 2201 8033 2235
rect 8251 2189 8285 2223
rect 8352 2184 8386 2218
rect 8436 2201 8470 2235
rect 8520 2184 8554 2218
rect 8604 2192 8638 2226
rect 8708 2184 8742 2218
rect 8792 2201 8826 2235
rect 8876 2184 8910 2218
rect 8960 2184 8994 2218
rect 9149 2197 9183 2231
rect 9233 2161 9267 2195
rect 9852 2161 9886 2195
rect 9951 2201 9985 2235
rect 10203 2189 10237 2223
rect 10304 2184 10338 2218
rect 10388 2201 10422 2235
rect 10472 2184 10506 2218
rect 10556 2192 10590 2226
rect 10660 2184 10694 2218
rect 10744 2201 10778 2235
rect 10828 2184 10862 2218
rect 10912 2184 10946 2218
rect 11101 2197 11135 2231
rect 11185 2161 11219 2195
rect 11844 2161 11878 2195
rect 11943 2201 11977 2235
rect 12195 2189 12229 2223
rect 12296 2184 12330 2218
rect 12380 2201 12414 2235
rect 12464 2184 12498 2218
rect 12548 2192 12582 2226
rect 12652 2184 12686 2218
rect 12736 2201 12770 2235
rect 12820 2184 12854 2218
rect 12904 2184 12938 2218
rect 13093 2197 13127 2231
rect 13177 2161 13211 2195
rect 13796 2161 13830 2195
rect 13895 2201 13929 2235
rect 14147 2189 14181 2223
rect 14248 2184 14282 2218
rect 14332 2201 14366 2235
rect 14416 2184 14450 2218
rect 14500 2192 14534 2226
rect 14604 2184 14638 2218
rect 14688 2201 14722 2235
rect 14772 2184 14806 2218
rect 14856 2184 14890 2218
rect 15045 2197 15079 2231
rect 15129 2161 15163 2195
rect 15860 2161 15894 2195
rect 15959 2201 15993 2235
rect 16211 2189 16245 2223
rect 16312 2184 16346 2218
rect 16396 2201 16430 2235
rect 16480 2184 16514 2218
rect 16564 2192 16598 2226
rect 16668 2184 16702 2218
rect 16752 2201 16786 2235
rect 16836 2184 16870 2218
rect 16920 2184 16954 2218
rect 17109 2197 17143 2231
rect 17193 2161 17227 2195
<< pdiffc >>
rect 9377 16497 9411 16531
rect 9377 16429 9411 16463
rect 9545 16487 9579 16521
rect 9545 16419 9579 16453
rect 9629 16487 9663 16521
rect 9629 16419 9663 16453
rect 9713 16487 9747 16521
rect 9817 16487 9851 16521
rect 9817 16419 9851 16453
rect 9901 16489 9935 16523
rect 9901 16421 9935 16455
rect 9901 16353 9935 16387
rect 9503 15711 9537 15745
rect 9587 15711 9621 15745
rect 9695 15753 9729 15787
rect 9695 15685 9729 15719
rect 9799 15753 9833 15787
rect 9799 15685 9833 15719
rect 11509 15643 11543 15677
rect 11601 15635 11635 15669
rect 11703 15643 11737 15677
rect 11798 15635 11832 15669
rect 11949 15643 11983 15677
rect 11949 15575 11983 15609
rect 12049 15643 12083 15677
rect 12049 15575 12083 15609
rect 12049 15507 12083 15541
rect 10687 15101 10721 15135
rect 10771 15101 10805 15135
rect 10879 15143 10913 15177
rect 10879 15075 10913 15109
rect 9387 14933 9421 14967
rect 9387 14865 9421 14899
rect 9555 14923 9589 14957
rect 9555 14855 9589 14889
rect 9639 14923 9673 14957
rect 9639 14855 9673 14889
rect 9723 14923 9757 14957
rect 9827 14923 9861 14957
rect 9827 14855 9861 14889
rect 9911 14925 9945 14959
rect 9911 14857 9945 14891
rect 10983 15143 11017 15177
rect 10983 15075 11017 15109
rect 9911 14789 9945 14823
rect 9513 14147 9547 14181
rect 9597 14147 9631 14181
rect 9705 14189 9739 14223
rect 9705 14121 9739 14155
rect 9809 14189 9843 14223
rect 9809 14121 9843 14155
rect 10725 14177 10759 14211
rect 10817 14169 10851 14203
rect 10919 14177 10953 14211
rect 11014 14169 11048 14203
rect 11165 14177 11199 14211
rect 11165 14109 11199 14143
rect 11265 14177 11299 14211
rect 11265 14109 11299 14143
rect 12984 14161 13018 14195
rect 12984 14093 13018 14127
rect 11265 14041 11299 14075
rect 12623 14030 12657 14064
rect 13069 14130 13103 14164
rect 13069 14062 13103 14096
rect 11905 13787 11939 13821
rect 11736 13667 11770 13701
rect 11905 13719 11939 13753
rect 12005 13803 12039 13837
rect 12005 13735 12039 13769
rect 9379 13265 9413 13299
rect 9379 13197 9413 13231
rect 9547 13255 9581 13289
rect 9547 13187 9581 13221
rect 9631 13255 9665 13289
rect 9631 13187 9665 13221
rect 9715 13255 9749 13289
rect 9819 13255 9853 13289
rect 9819 13187 9853 13221
rect 11121 13335 11155 13369
rect 9903 13257 9937 13291
rect 9903 13189 9937 13223
rect 10849 13196 10883 13230
rect 10933 13226 10967 13260
rect 11026 13207 11060 13241
rect 9903 13121 9937 13155
rect 11205 13321 11239 13355
rect 11205 13253 11239 13287
rect 9505 12479 9539 12513
rect 9589 12479 9623 12513
rect 9697 12521 9731 12555
rect 9697 12453 9731 12487
rect 9801 12521 9835 12555
rect 9801 12453 9835 12487
rect 10881 12273 10915 12307
rect 10965 12273 10999 12307
rect 11073 12315 11107 12349
rect 11073 12247 11107 12281
rect 11177 12315 11211 12349
rect 11177 12247 11211 12281
rect 9389 11701 9423 11735
rect 9389 11633 9423 11667
rect 9557 11691 9591 11725
rect 9557 11623 9591 11657
rect 9641 11691 9675 11725
rect 9641 11623 9675 11657
rect 9725 11691 9759 11725
rect 9829 11691 9863 11725
rect 9829 11623 9863 11657
rect 9913 11693 9947 11727
rect 9913 11625 9947 11659
rect 9913 11557 9947 11591
rect 9515 10915 9549 10949
rect 9599 10915 9633 10949
rect 9707 10957 9741 10991
rect 9707 10889 9741 10923
rect 9811 10957 9845 10991
rect 9811 10889 9845 10923
rect 6194 6251 6228 6285
rect 6194 6183 6228 6217
rect 6194 6115 6228 6149
rect 6278 6251 6312 6285
rect 6278 6183 6312 6217
rect 6278 6115 6312 6149
rect 10088 5599 10122 5633
rect 1906 5179 1940 5213
rect 1906 5089 1940 5123
rect 10088 5509 10122 5543
rect 1990 5059 2024 5093
rect 2257 5071 2291 5105
rect 2358 5076 2392 5110
rect 2442 5059 2476 5093
rect 2526 5076 2560 5110
rect 2610 5063 2644 5097
rect 2714 5076 2748 5110
rect 2798 5059 2832 5093
rect 2882 5076 2916 5110
rect 2966 5076 3000 5110
rect 3155 5067 3189 5101
rect 3239 5176 3273 5210
rect 3239 5082 3273 5116
rect 4040 5171 4074 5205
rect 4040 5081 4074 5115
rect 4124 5051 4158 5085
rect 4391 5063 4425 5097
rect 4492 5068 4526 5102
rect 4576 5051 4610 5085
rect 4660 5068 4694 5102
rect 4744 5055 4778 5089
rect 4848 5068 4882 5102
rect 4932 5051 4966 5085
rect 5016 5068 5050 5102
rect 5100 5068 5134 5102
rect 5289 5059 5323 5093
rect 5373 5168 5407 5202
rect 5373 5074 5407 5108
rect 5992 5171 6026 5205
rect 5992 5081 6026 5115
rect 6076 5051 6110 5085
rect 6343 5063 6377 5097
rect 6444 5068 6478 5102
rect 6528 5051 6562 5085
rect 6612 5068 6646 5102
rect 6696 5055 6730 5089
rect 6800 5068 6834 5102
rect 6884 5051 6918 5085
rect 6968 5068 7002 5102
rect 7052 5068 7086 5102
rect 7241 5059 7275 5093
rect 7325 5168 7359 5202
rect 7325 5074 7359 5108
rect 7994 5177 8028 5211
rect 7994 5087 8028 5121
rect 10172 5479 10206 5513
rect 10439 5491 10473 5525
rect 10540 5496 10574 5530
rect 10624 5479 10658 5513
rect 10708 5496 10742 5530
rect 10792 5483 10826 5517
rect 10896 5496 10930 5530
rect 10980 5479 11014 5513
rect 11064 5496 11098 5530
rect 11148 5496 11182 5530
rect 11337 5487 11371 5521
rect 11421 5596 11455 5630
rect 11421 5502 11455 5536
rect 12150 5587 12184 5621
rect 12150 5497 12184 5531
rect 12234 5467 12268 5501
rect 12501 5479 12535 5513
rect 12602 5484 12636 5518
rect 12686 5467 12720 5501
rect 12770 5484 12804 5518
rect 12854 5471 12888 5505
rect 12958 5484 12992 5518
rect 13042 5467 13076 5501
rect 13126 5484 13160 5518
rect 13210 5484 13244 5518
rect 13399 5475 13433 5509
rect 13483 5584 13517 5618
rect 13483 5490 13517 5524
rect 14108 5595 14142 5629
rect 14108 5505 14142 5539
rect 14192 5475 14226 5509
rect 14459 5487 14493 5521
rect 14560 5492 14594 5526
rect 14644 5475 14678 5509
rect 14728 5492 14762 5526
rect 14812 5479 14846 5513
rect 14916 5492 14950 5526
rect 15000 5475 15034 5509
rect 15084 5492 15118 5526
rect 15168 5492 15202 5526
rect 15357 5483 15391 5517
rect 15441 5592 15475 5626
rect 15441 5498 15475 5532
rect 16102 5601 16136 5635
rect 16102 5511 16136 5545
rect 16186 5481 16220 5515
rect 16453 5493 16487 5527
rect 16554 5498 16588 5532
rect 16638 5481 16672 5515
rect 16722 5498 16756 5532
rect 16806 5485 16840 5519
rect 16910 5498 16944 5532
rect 16994 5481 17028 5515
rect 17078 5498 17112 5532
rect 17162 5498 17196 5532
rect 17351 5489 17385 5523
rect 17435 5598 17469 5632
rect 17435 5504 17469 5538
rect 8078 5057 8112 5091
rect 8345 5069 8379 5103
rect 8446 5074 8480 5108
rect 8530 5057 8564 5091
rect 8614 5074 8648 5108
rect 8698 5061 8732 5095
rect 8802 5074 8836 5108
rect 8886 5057 8920 5091
rect 8970 5074 9004 5108
rect 9054 5074 9088 5108
rect 9243 5065 9277 5099
rect 9327 5174 9361 5208
rect 9327 5080 9361 5114
rect 10116 4725 10150 4759
rect 10116 4635 10150 4669
rect 10200 4605 10234 4639
rect 10467 4617 10501 4651
rect 10568 4622 10602 4656
rect 10652 4605 10686 4639
rect 10736 4622 10770 4656
rect 10820 4609 10854 4643
rect 10924 4622 10958 4656
rect 11008 4605 11042 4639
rect 11092 4622 11126 4656
rect 11176 4622 11210 4656
rect 11365 4613 11399 4647
rect 11449 4722 11483 4756
rect 11449 4628 11483 4662
rect 12386 4681 12420 4715
rect 12386 4591 12420 4625
rect 12470 4561 12504 4595
rect 12737 4573 12771 4607
rect 12838 4578 12872 4612
rect 12922 4561 12956 4595
rect 13006 4578 13040 4612
rect 13090 4565 13124 4599
rect 13194 4578 13228 4612
rect 13278 4561 13312 4595
rect 13362 4578 13396 4612
rect 13446 4578 13480 4612
rect 13635 4569 13669 4603
rect 13719 4678 13753 4712
rect 13719 4584 13753 4618
rect 14388 4675 14422 4709
rect 14388 4585 14422 4619
rect 14472 4555 14506 4589
rect 14739 4567 14773 4601
rect 14840 4572 14874 4606
rect 14924 4555 14958 4589
rect 15008 4572 15042 4606
rect 15092 4559 15126 4593
rect 15196 4572 15230 4606
rect 15280 4555 15314 4589
rect 15364 4572 15398 4606
rect 15448 4572 15482 4606
rect 15637 4563 15671 4597
rect 15721 4672 15755 4706
rect 15721 4578 15755 4612
rect 16410 4657 16444 4691
rect 16410 4567 16444 4601
rect 16494 4537 16528 4571
rect 16761 4549 16795 4583
rect 16862 4554 16896 4588
rect 16946 4537 16980 4571
rect 17030 4554 17064 4588
rect 17114 4541 17148 4575
rect 17218 4554 17252 4588
rect 17302 4537 17336 4571
rect 17386 4554 17420 4588
rect 17470 4554 17504 4588
rect 17659 4545 17693 4579
rect 17743 4654 17777 4688
rect 17743 4560 17777 4594
rect 1876 1919 1910 1953
rect 1876 1829 1910 1863
rect 1960 1799 1994 1833
rect 2227 1811 2261 1845
rect 2328 1816 2362 1850
rect 2412 1799 2446 1833
rect 2496 1816 2530 1850
rect 2580 1803 2614 1837
rect 2684 1816 2718 1850
rect 2768 1799 2802 1833
rect 2852 1816 2886 1850
rect 2936 1816 2970 1850
rect 3125 1807 3159 1841
rect 3209 1916 3243 1950
rect 3209 1822 3243 1856
rect 3946 1915 3980 1949
rect 3946 1825 3980 1859
rect 4030 1795 4064 1829
rect 4297 1807 4331 1841
rect 4398 1812 4432 1846
rect 4482 1795 4516 1829
rect 4566 1812 4600 1846
rect 4650 1799 4684 1833
rect 4754 1812 4788 1846
rect 4838 1795 4872 1829
rect 4922 1812 4956 1846
rect 5006 1812 5040 1846
rect 5195 1803 5229 1837
rect 5279 1912 5313 1946
rect 5279 1818 5313 1852
rect 5898 1915 5932 1949
rect 5898 1825 5932 1859
rect 5982 1795 6016 1829
rect 6249 1807 6283 1841
rect 6350 1812 6384 1846
rect 6434 1795 6468 1829
rect 6518 1812 6552 1846
rect 6602 1799 6636 1833
rect 6706 1812 6740 1846
rect 6790 1795 6824 1829
rect 6874 1812 6908 1846
rect 6958 1812 6992 1846
rect 7147 1803 7181 1837
rect 7231 1912 7265 1946
rect 7231 1818 7265 1852
rect 7900 1921 7934 1955
rect 7900 1831 7934 1865
rect 7984 1801 8018 1835
rect 8251 1813 8285 1847
rect 8352 1818 8386 1852
rect 8436 1801 8470 1835
rect 8520 1818 8554 1852
rect 8604 1805 8638 1839
rect 8708 1818 8742 1852
rect 8792 1801 8826 1835
rect 8876 1818 8910 1852
rect 8960 1818 8994 1852
rect 9149 1809 9183 1843
rect 9233 1918 9267 1952
rect 9233 1824 9267 1858
rect 9852 1921 9886 1955
rect 9852 1831 9886 1865
rect 9936 1801 9970 1835
rect 10203 1813 10237 1847
rect 10304 1818 10338 1852
rect 10388 1801 10422 1835
rect 10472 1818 10506 1852
rect 10556 1805 10590 1839
rect 10660 1818 10694 1852
rect 10744 1801 10778 1835
rect 10828 1818 10862 1852
rect 10912 1818 10946 1852
rect 11101 1809 11135 1843
rect 11185 1918 11219 1952
rect 11185 1824 11219 1858
rect 11844 1921 11878 1955
rect 11844 1831 11878 1865
rect 11928 1801 11962 1835
rect 12195 1813 12229 1847
rect 12296 1818 12330 1852
rect 12380 1801 12414 1835
rect 12464 1818 12498 1852
rect 12548 1805 12582 1839
rect 12652 1818 12686 1852
rect 12736 1801 12770 1835
rect 12820 1818 12854 1852
rect 12904 1818 12938 1852
rect 13093 1809 13127 1843
rect 13177 1918 13211 1952
rect 13177 1824 13211 1858
rect 13796 1921 13830 1955
rect 13796 1831 13830 1865
rect 13880 1801 13914 1835
rect 14147 1813 14181 1847
rect 14248 1818 14282 1852
rect 14332 1801 14366 1835
rect 14416 1818 14450 1852
rect 14500 1805 14534 1839
rect 14604 1818 14638 1852
rect 14688 1801 14722 1835
rect 14772 1818 14806 1852
rect 14856 1818 14890 1852
rect 15045 1809 15079 1843
rect 15129 1918 15163 1952
rect 15129 1824 15163 1858
rect 15860 1921 15894 1955
rect 15860 1831 15894 1865
rect 15944 1801 15978 1835
rect 16211 1813 16245 1847
rect 16312 1818 16346 1852
rect 16396 1801 16430 1835
rect 16480 1818 16514 1852
rect 16564 1805 16598 1839
rect 16668 1818 16702 1852
rect 16752 1801 16786 1835
rect 16836 1818 16870 1852
rect 16920 1818 16954 1852
rect 17109 1809 17143 1843
rect 17193 1918 17227 1952
rect 17193 1824 17227 1858
<< poly >>
rect 9421 16543 9451 16569
rect 9505 16543 9535 16569
rect 9589 16543 9619 16569
rect 9673 16543 9703 16569
rect 9861 16543 9891 16569
rect 9421 16311 9451 16343
rect 9505 16311 9535 16343
rect 9589 16311 9619 16343
rect 9673 16311 9703 16343
rect 9861 16311 9891 16343
rect 9409 16295 9463 16311
rect 9409 16261 9419 16295
rect 9453 16261 9463 16295
rect 9409 16245 9463 16261
rect 9505 16295 9619 16311
rect 9505 16261 9536 16295
rect 9570 16261 9619 16295
rect 9505 16245 9619 16261
rect 9661 16295 9715 16311
rect 9661 16261 9671 16295
rect 9705 16261 9715 16295
rect 9661 16245 9715 16261
rect 9757 16295 9891 16311
rect 9757 16261 9767 16295
rect 9801 16278 9891 16295
rect 9801 16261 9887 16278
rect 9757 16245 9887 16261
rect 9421 16223 9451 16245
rect 9505 16223 9535 16245
rect 9589 16223 9619 16245
rect 9673 16223 9703 16245
rect 9857 16223 9887 16245
rect 9421 16067 9451 16093
rect 9505 16067 9535 16093
rect 9589 16067 9619 16093
rect 9673 16067 9703 16093
rect 9857 16067 9887 16093
rect 9739 15799 9769 15825
rect 9547 15757 9577 15783
rect 9631 15757 9661 15783
rect 9547 15567 9577 15673
rect 9490 15551 9577 15567
rect 9490 15517 9506 15551
rect 9540 15517 9577 15551
rect 9490 15501 9577 15517
rect 9547 15461 9577 15501
rect 9631 15567 9661 15673
rect 11553 15689 11583 15715
rect 11653 15689 11683 15715
rect 11757 15689 11787 15715
rect 11843 15689 11873 15715
rect 12009 15689 12039 15715
rect 9739 15567 9769 15599
rect 9631 15551 9697 15567
rect 9631 15517 9647 15551
rect 9681 15517 9697 15551
rect 9631 15501 9697 15517
rect 9739 15551 9805 15567
rect 9739 15517 9755 15551
rect 9789 15517 9805 15551
rect 9739 15501 9805 15517
rect 9631 15461 9661 15501
rect 9739 15479 9769 15501
rect 9547 15351 9577 15377
rect 9631 15351 9661 15377
rect 11553 15457 11583 15605
rect 11653 15457 11683 15605
rect 11757 15457 11787 15605
rect 11843 15457 11873 15605
rect 12009 15457 12039 15489
rect 11495 15441 11583 15457
rect 11495 15407 11505 15441
rect 11539 15407 11583 15441
rect 11495 15391 11583 15407
rect 9739 15323 9769 15349
rect 11553 15323 11583 15391
rect 11641 15441 11695 15457
rect 11641 15407 11651 15441
rect 11685 15407 11695 15441
rect 11641 15391 11695 15407
rect 11747 15441 11801 15457
rect 11747 15407 11757 15441
rect 11791 15407 11801 15441
rect 11747 15391 11801 15407
rect 11843 15441 11907 15457
rect 11843 15407 11853 15441
rect 11887 15407 11907 15441
rect 11843 15391 11907 15407
rect 11954 15441 12039 15457
rect 11954 15407 11964 15441
rect 11998 15407 12039 15441
rect 11954 15391 12039 15407
rect 11641 15323 11671 15391
rect 11747 15323 11777 15391
rect 11843 15323 11873 15391
rect 12009 15369 12039 15391
rect 10923 15189 10953 15215
rect 11553 15213 11583 15239
rect 11641 15213 11671 15239
rect 11747 15213 11777 15239
rect 11843 15213 11873 15239
rect 12009 15213 12039 15239
rect 10731 15147 10761 15173
rect 10815 15147 10845 15173
rect 9431 14979 9461 15005
rect 9515 14979 9545 15005
rect 9599 14979 9629 15005
rect 9683 14979 9713 15005
rect 9871 14979 9901 15005
rect 10731 14957 10761 15063
rect 10674 14941 10761 14957
rect 10674 14907 10690 14941
rect 10724 14907 10761 14941
rect 10674 14891 10761 14907
rect 10731 14851 10761 14891
rect 10815 14957 10845 15063
rect 10923 14957 10953 14989
rect 10815 14941 10881 14957
rect 10815 14907 10831 14941
rect 10865 14907 10881 14941
rect 10815 14891 10881 14907
rect 10923 14941 10989 14957
rect 10923 14907 10939 14941
rect 10973 14907 10989 14941
rect 10923 14891 10989 14907
rect 10815 14851 10845 14891
rect 10923 14869 10953 14891
rect 9431 14747 9461 14779
rect 9515 14747 9545 14779
rect 9599 14747 9629 14779
rect 9683 14747 9713 14779
rect 9871 14747 9901 14779
rect 9419 14731 9473 14747
rect 9419 14697 9429 14731
rect 9463 14697 9473 14731
rect 9419 14681 9473 14697
rect 9515 14731 9629 14747
rect 9515 14697 9546 14731
rect 9580 14697 9629 14731
rect 9515 14681 9629 14697
rect 9671 14731 9725 14747
rect 9671 14697 9681 14731
rect 9715 14697 9725 14731
rect 9671 14681 9725 14697
rect 9767 14731 9901 14747
rect 10731 14741 10761 14767
rect 10815 14741 10845 14767
rect 9767 14697 9777 14731
rect 9811 14714 9901 14731
rect 9811 14697 9897 14714
rect 10923 14713 10953 14739
rect 9767 14681 9897 14697
rect 9431 14659 9461 14681
rect 9515 14659 9545 14681
rect 9599 14659 9629 14681
rect 9683 14659 9713 14681
rect 9867 14659 9897 14681
rect 9431 14503 9461 14529
rect 9515 14503 9545 14529
rect 9599 14503 9629 14529
rect 9683 14503 9713 14529
rect 9867 14503 9897 14529
rect 9749 14235 9779 14261
rect 9557 14193 9587 14219
rect 9641 14193 9671 14219
rect 9557 14003 9587 14109
rect 9500 13987 9587 14003
rect 9500 13953 9516 13987
rect 9550 13953 9587 13987
rect 9500 13937 9587 13953
rect 9557 13897 9587 13937
rect 9641 14003 9671 14109
rect 10769 14223 10799 14249
rect 10869 14223 10899 14249
rect 10973 14223 11003 14249
rect 11059 14223 11089 14249
rect 11225 14223 11255 14249
rect 9749 14003 9779 14035
rect 9641 13987 9707 14003
rect 9641 13953 9657 13987
rect 9691 13953 9707 13987
rect 9641 13937 9707 13953
rect 9749 13987 9815 14003
rect 10769 13991 10799 14139
rect 10869 13991 10899 14139
rect 10973 13991 11003 14139
rect 11059 13991 11089 14139
rect 13029 14207 13059 14233
rect 12829 14183 12895 14193
rect 12829 14149 12845 14183
rect 12879 14149 12895 14183
rect 12829 14139 12895 14149
rect 12667 14091 12697 14117
rect 12763 14091 12793 14117
rect 12835 14091 12865 14139
rect 12931 14091 12961 14117
rect 11225 13991 11255 14023
rect 9749 13953 9765 13987
rect 9799 13953 9815 13987
rect 9749 13937 9815 13953
rect 10711 13975 10799 13991
rect 10711 13941 10721 13975
rect 10755 13941 10799 13975
rect 9641 13897 9671 13937
rect 9749 13915 9779 13937
rect 10711 13925 10799 13941
rect 9557 13787 9587 13813
rect 9641 13787 9671 13813
rect 10769 13857 10799 13925
rect 10857 13975 10911 13991
rect 10857 13941 10867 13975
rect 10901 13941 10911 13975
rect 10857 13925 10911 13941
rect 10963 13975 11017 13991
rect 10963 13941 10973 13975
rect 11007 13941 11017 13975
rect 10963 13925 11017 13941
rect 11059 13975 11123 13991
rect 11059 13941 11069 13975
rect 11103 13941 11123 13975
rect 11059 13925 11123 13941
rect 11170 13975 11255 13991
rect 12667 13975 12697 14007
rect 12763 13975 12793 14007
rect 11170 13941 11180 13975
rect 11214 13941 11255 13975
rect 11170 13925 11255 13941
rect 10857 13857 10887 13925
rect 10963 13857 10993 13925
rect 11059 13857 11089 13925
rect 11225 13903 11255 13925
rect 12613 13959 12697 13975
rect 12613 13925 12623 13959
rect 12657 13925 12697 13959
rect 12613 13909 12697 13925
rect 12739 13959 12793 13975
rect 12739 13925 12749 13959
rect 12783 13925 12793 13959
rect 12739 13909 12793 13925
rect 9749 13759 9779 13785
rect 11949 13849 11979 13875
rect 10769 13747 10799 13773
rect 10857 13747 10887 13773
rect 10963 13747 10993 13773
rect 11059 13747 11089 13773
rect 11225 13747 11255 13773
rect 11780 13733 11810 13759
rect 11852 13733 11882 13759
rect 12667 13847 12697 13909
rect 12763 13847 12793 13909
rect 12835 13892 12865 14007
rect 12931 13975 12961 14007
rect 13029 13975 13059 14007
rect 12915 13959 12969 13975
rect 12915 13925 12925 13959
rect 12959 13925 12969 13959
rect 12915 13909 12969 13925
rect 13011 13959 13066 13975
rect 13011 13925 13021 13959
rect 13055 13925 13066 13959
rect 13011 13909 13066 13925
rect 12835 13891 12876 13892
rect 12835 13862 12877 13891
rect 12847 13847 12877 13862
rect 12931 13847 12961 13909
rect 13029 13887 13059 13909
rect 12667 13737 12697 13763
rect 12763 13737 12793 13763
rect 12847 13737 12877 13763
rect 12931 13737 12961 13763
rect 13029 13731 13059 13757
rect 11780 13617 11810 13649
rect 11710 13601 11810 13617
rect 11710 13567 11726 13601
rect 11760 13567 11810 13601
rect 11710 13551 11810 13567
rect 11852 13617 11882 13649
rect 11949 13617 11979 13649
rect 11852 13601 11906 13617
rect 11852 13567 11862 13601
rect 11896 13567 11906 13601
rect 11852 13551 11906 13567
rect 11949 13601 12015 13617
rect 11949 13567 11965 13601
rect 11999 13567 12015 13601
rect 11949 13551 12015 13567
rect 11768 13483 11798 13551
rect 11852 13483 11882 13551
rect 11949 13529 11979 13551
rect 11165 13381 11195 13407
rect 10977 13360 11031 13376
rect 9423 13311 9453 13337
rect 9507 13311 9537 13337
rect 9591 13311 9621 13337
rect 9675 13311 9705 13337
rect 9863 13311 9893 13337
rect 10977 13326 10987 13360
rect 11021 13326 11031 13360
rect 10977 13310 11031 13326
rect 10893 13268 10923 13309
rect 10977 13268 11007 13310
rect 11070 13268 11100 13294
rect 10893 13135 10923 13184
rect 10977 13166 11007 13184
rect 9423 13079 9453 13111
rect 9507 13079 9537 13111
rect 9591 13079 9621 13111
rect 9675 13079 9705 13111
rect 9863 13079 9893 13111
rect 9411 13063 9465 13079
rect 9411 13029 9421 13063
rect 9455 13029 9465 13063
rect 9411 13013 9465 13029
rect 9507 13063 9621 13079
rect 9507 13029 9538 13063
rect 9572 13029 9621 13063
rect 9507 13013 9621 13029
rect 9663 13063 9717 13079
rect 9663 13029 9673 13063
rect 9707 13029 9717 13063
rect 9663 13013 9717 13029
rect 9759 13063 9893 13079
rect 9759 13029 9769 13063
rect 9803 13046 9893 13063
rect 10839 13087 10923 13135
rect 10839 13053 10849 13087
rect 10883 13053 10923 13087
rect 9803 13029 9889 13046
rect 10839 13030 10923 13053
rect 9759 13013 9889 13029
rect 10893 13015 10923 13030
rect 10965 13141 11007 13166
rect 11070 13143 11100 13184
rect 11768 13373 11798 13399
rect 11852 13373 11882 13399
rect 11949 13373 11979 13399
rect 11165 13149 11195 13181
rect 10965 13015 10995 13141
rect 11049 13127 11103 13143
rect 11049 13110 11059 13127
rect 11037 13093 11059 13110
rect 11093 13093 11103 13127
rect 11037 13077 11103 13093
rect 11145 13133 11199 13149
rect 11145 13099 11155 13133
rect 11189 13099 11199 13133
rect 11145 13083 11199 13099
rect 11037 13054 11079 13077
rect 11165 13061 11195 13083
rect 11037 13030 11074 13054
rect 11037 13015 11067 13030
rect 9423 12991 9453 13013
rect 9507 12991 9537 13013
rect 9591 12991 9621 13013
rect 9675 12991 9705 13013
rect 9859 12991 9889 13013
rect 10893 12905 10923 12931
rect 10965 12905 10995 12931
rect 11037 12905 11067 12931
rect 11165 12905 11195 12931
rect 9423 12835 9453 12861
rect 9507 12835 9537 12861
rect 9591 12835 9621 12861
rect 9675 12835 9705 12861
rect 9859 12835 9889 12861
rect 9741 12567 9771 12593
rect 9549 12525 9579 12551
rect 9633 12525 9663 12551
rect 9549 12335 9579 12441
rect 9492 12319 9579 12335
rect 9492 12285 9508 12319
rect 9542 12285 9579 12319
rect 9492 12269 9579 12285
rect 9549 12229 9579 12269
rect 9633 12335 9663 12441
rect 9741 12335 9771 12367
rect 11117 12361 11147 12387
rect 9633 12319 9699 12335
rect 9633 12285 9649 12319
rect 9683 12285 9699 12319
rect 9633 12269 9699 12285
rect 9741 12319 9807 12335
rect 10925 12319 10955 12345
rect 11009 12319 11039 12345
rect 9741 12285 9757 12319
rect 9791 12285 9807 12319
rect 9741 12269 9807 12285
rect 9633 12229 9663 12269
rect 9741 12247 9771 12269
rect 9549 12119 9579 12145
rect 9633 12119 9663 12145
rect 10925 12129 10955 12235
rect 9741 12091 9771 12117
rect 10868 12113 10955 12129
rect 10868 12079 10884 12113
rect 10918 12079 10955 12113
rect 10868 12063 10955 12079
rect 10925 12023 10955 12063
rect 11009 12129 11039 12235
rect 11117 12129 11147 12161
rect 11009 12113 11075 12129
rect 11009 12079 11025 12113
rect 11059 12079 11075 12113
rect 11009 12063 11075 12079
rect 11117 12113 11183 12129
rect 11117 12079 11133 12113
rect 11167 12079 11183 12113
rect 11117 12063 11183 12079
rect 11009 12023 11039 12063
rect 11117 12041 11147 12063
rect 10925 11913 10955 11939
rect 11009 11913 11039 11939
rect 11117 11885 11147 11911
rect 9433 11747 9463 11773
rect 9517 11747 9547 11773
rect 9601 11747 9631 11773
rect 9685 11747 9715 11773
rect 9873 11747 9903 11773
rect 9433 11515 9463 11547
rect 9517 11515 9547 11547
rect 9601 11515 9631 11547
rect 9685 11515 9715 11547
rect 9873 11515 9903 11547
rect 9421 11499 9475 11515
rect 9421 11465 9431 11499
rect 9465 11465 9475 11499
rect 9421 11449 9475 11465
rect 9517 11499 9631 11515
rect 9517 11465 9548 11499
rect 9582 11465 9631 11499
rect 9517 11449 9631 11465
rect 9673 11499 9727 11515
rect 9673 11465 9683 11499
rect 9717 11465 9727 11499
rect 9673 11449 9727 11465
rect 9769 11499 9903 11515
rect 9769 11465 9779 11499
rect 9813 11482 9903 11499
rect 9813 11465 9899 11482
rect 9769 11449 9899 11465
rect 9433 11427 9463 11449
rect 9517 11427 9547 11449
rect 9601 11427 9631 11449
rect 9685 11427 9715 11449
rect 9869 11427 9899 11449
rect 9433 11271 9463 11297
rect 9517 11271 9547 11297
rect 9601 11271 9631 11297
rect 9685 11271 9715 11297
rect 9869 11271 9899 11297
rect 9751 11003 9781 11029
rect 9559 10961 9589 10987
rect 9643 10961 9673 10987
rect 9559 10771 9589 10877
rect 9502 10755 9589 10771
rect 9502 10721 9518 10755
rect 9552 10721 9589 10755
rect 9502 10705 9589 10721
rect 9559 10665 9589 10705
rect 9643 10771 9673 10877
rect 9751 10771 9781 10803
rect 9643 10755 9709 10771
rect 9643 10721 9659 10755
rect 9693 10721 9709 10755
rect 9643 10705 9709 10721
rect 9751 10755 9817 10771
rect 9751 10721 9767 10755
rect 9801 10721 9817 10755
rect 9751 10705 9817 10721
rect 9643 10665 9673 10705
rect 9751 10683 9781 10705
rect 9559 10555 9589 10581
rect 9643 10555 9673 10581
rect 9751 10527 9781 10553
rect 6238 6553 6268 6579
rect 6238 6401 6268 6423
rect 6238 6385 6324 6401
rect 6238 6351 6274 6385
rect 6308 6351 6324 6385
rect 6238 6335 6324 6351
rect 6238 6303 6268 6335
rect 6238 6077 6268 6103
rect 10132 5921 10162 5947
rect 10231 5921 10261 5947
rect 10327 5921 10357 5947
rect 10399 5921 10429 5947
rect 10495 5921 10525 5947
rect 10584 5921 10614 5947
rect 10668 5921 10698 5947
rect 10752 5921 10782 5947
rect 10940 5921 10970 5947
rect 11024 5921 11054 5947
rect 11108 5921 11138 5947
rect 11192 5921 11222 5947
rect 11282 5921 11312 5947
rect 11381 5921 11411 5947
rect 10132 5769 10162 5791
rect 10231 5777 10261 5837
rect 10132 5753 10186 5769
rect 10132 5719 10142 5753
rect 10176 5719 10186 5753
rect 10132 5703 10186 5719
rect 10231 5761 10285 5777
rect 10231 5727 10241 5761
rect 10275 5727 10285 5761
rect 10231 5711 10285 5727
rect 10132 5671 10162 5703
rect 1950 5501 1980 5527
rect 2049 5501 2079 5527
rect 2145 5501 2175 5527
rect 2217 5501 2247 5527
rect 2313 5501 2343 5527
rect 2402 5501 2432 5527
rect 2486 5501 2516 5527
rect 2570 5501 2600 5527
rect 2758 5501 2788 5527
rect 2842 5501 2872 5527
rect 2926 5501 2956 5527
rect 3010 5501 3040 5527
rect 3100 5501 3130 5527
rect 3199 5501 3229 5527
rect 1950 5349 1980 5371
rect 2049 5357 2079 5417
rect 1950 5333 2004 5349
rect 1950 5299 1960 5333
rect 1994 5299 2004 5333
rect 1950 5283 2004 5299
rect 2049 5341 2103 5357
rect 2049 5307 2059 5341
rect 2093 5307 2103 5341
rect 2049 5291 2103 5307
rect 1950 5251 1980 5283
rect 2049 5135 2079 5291
rect 2145 5245 2175 5417
rect 2121 5229 2175 5245
rect 2121 5195 2131 5229
rect 2165 5195 2175 5229
rect 2121 5179 2175 5195
rect 2145 5135 2175 5179
rect 2217 5245 2247 5417
rect 2313 5373 2343 5417
rect 2402 5373 2432 5417
rect 2486 5402 2516 5417
rect 2289 5357 2343 5373
rect 2289 5323 2299 5357
rect 2333 5323 2343 5357
rect 2289 5307 2343 5323
rect 2389 5357 2443 5373
rect 2389 5323 2399 5357
rect 2433 5323 2443 5357
rect 2389 5307 2443 5323
rect 2485 5372 2516 5402
rect 2570 5402 2600 5417
rect 2758 5402 2788 5417
rect 2570 5372 2788 5402
rect 2217 5229 2271 5245
rect 2217 5195 2227 5229
rect 2261 5195 2271 5229
rect 2217 5179 2271 5195
rect 2217 5135 2247 5179
rect 2313 5135 2343 5307
rect 2402 5135 2432 5307
rect 2485 5261 2515 5372
rect 2570 5357 2611 5372
rect 2581 5261 2611 5357
rect 2842 5342 2872 5417
rect 2926 5343 2956 5417
rect 2818 5326 2872 5342
rect 2818 5292 2828 5326
rect 2862 5292 2872 5326
rect 2818 5276 2872 5292
rect 2914 5327 2968 5343
rect 2914 5293 2924 5327
rect 2958 5293 2968 5327
rect 2914 5277 2968 5293
rect 2474 5245 2528 5261
rect 2474 5211 2484 5245
rect 2518 5211 2528 5245
rect 2474 5195 2528 5211
rect 2581 5245 2645 5261
rect 2581 5211 2601 5245
rect 2635 5211 2645 5245
rect 2486 5135 2516 5195
rect 2581 5180 2645 5211
rect 2570 5150 2788 5180
rect 2570 5135 2600 5150
rect 2758 5135 2788 5150
rect 2842 5135 2872 5276
rect 2926 5135 2956 5277
rect 3010 5238 3040 5417
rect 3100 5349 3130 5417
rect 4084 5493 4114 5519
rect 4183 5493 4213 5519
rect 4279 5493 4309 5519
rect 4351 5493 4381 5519
rect 4447 5493 4477 5519
rect 4536 5493 4566 5519
rect 4620 5493 4650 5519
rect 4704 5493 4734 5519
rect 4892 5493 4922 5519
rect 4976 5493 5006 5519
rect 5060 5493 5090 5519
rect 5144 5493 5174 5519
rect 5234 5493 5264 5519
rect 5333 5493 5363 5519
rect 6036 5493 6066 5519
rect 6135 5493 6165 5519
rect 6231 5493 6261 5519
rect 6303 5493 6333 5519
rect 6399 5493 6429 5519
rect 6488 5493 6518 5519
rect 6572 5493 6602 5519
rect 6656 5493 6686 5519
rect 6844 5493 6874 5519
rect 6928 5493 6958 5519
rect 7012 5493 7042 5519
rect 7096 5493 7126 5519
rect 7186 5493 7216 5519
rect 7285 5493 7315 5519
rect 8038 5499 8068 5525
rect 8137 5499 8167 5525
rect 8233 5499 8263 5525
rect 8305 5499 8335 5525
rect 8401 5499 8431 5525
rect 8490 5499 8520 5525
rect 8574 5499 8604 5525
rect 8658 5499 8688 5525
rect 8846 5499 8876 5525
rect 8930 5499 8960 5525
rect 9014 5499 9044 5525
rect 9098 5499 9128 5525
rect 9188 5499 9218 5525
rect 9287 5499 9317 5525
rect 3199 5349 3229 5371
rect 3082 5333 3136 5349
rect 3082 5299 3092 5333
rect 3126 5299 3136 5333
rect 3082 5283 3136 5299
rect 3178 5333 3232 5349
rect 3178 5299 3188 5333
rect 3222 5299 3232 5333
rect 3178 5283 3232 5299
rect 4084 5341 4114 5363
rect 4183 5349 4213 5409
rect 4084 5325 4138 5341
rect 4084 5291 4094 5325
rect 4128 5291 4138 5325
rect 3004 5222 3058 5238
rect 3004 5188 3014 5222
rect 3048 5188 3058 5222
rect 3004 5172 3058 5188
rect 3010 5135 3040 5172
rect 3100 5135 3130 5283
rect 3199 5251 3229 5283
rect 4084 5275 4138 5291
rect 4183 5333 4237 5349
rect 4183 5299 4193 5333
rect 4227 5299 4237 5333
rect 4183 5283 4237 5299
rect 4084 5243 4114 5275
rect 1950 5025 1980 5051
rect 2049 5025 2079 5051
rect 2145 5025 2175 5051
rect 2217 5025 2247 5051
rect 2313 5025 2343 5051
rect 2402 5025 2432 5051
rect 2486 5025 2516 5051
rect 2570 5025 2600 5051
rect 2758 5025 2788 5051
rect 2842 5025 2872 5051
rect 2926 5025 2956 5051
rect 3010 5025 3040 5051
rect 3100 5025 3130 5051
rect 3199 5025 3229 5051
rect 4183 5127 4213 5283
rect 4279 5237 4309 5409
rect 4255 5221 4309 5237
rect 4255 5187 4265 5221
rect 4299 5187 4309 5221
rect 4255 5171 4309 5187
rect 4279 5127 4309 5171
rect 4351 5237 4381 5409
rect 4447 5365 4477 5409
rect 4536 5365 4566 5409
rect 4620 5394 4650 5409
rect 4423 5349 4477 5365
rect 4423 5315 4433 5349
rect 4467 5315 4477 5349
rect 4423 5299 4477 5315
rect 4523 5349 4577 5365
rect 4523 5315 4533 5349
rect 4567 5315 4577 5349
rect 4523 5299 4577 5315
rect 4619 5364 4650 5394
rect 4704 5394 4734 5409
rect 4892 5394 4922 5409
rect 4704 5364 4922 5394
rect 4351 5221 4405 5237
rect 4351 5187 4361 5221
rect 4395 5187 4405 5221
rect 4351 5171 4405 5187
rect 4351 5127 4381 5171
rect 4447 5127 4477 5299
rect 4536 5127 4566 5299
rect 4619 5253 4649 5364
rect 4704 5349 4745 5364
rect 4715 5253 4745 5349
rect 4976 5334 5006 5409
rect 5060 5335 5090 5409
rect 4952 5318 5006 5334
rect 4952 5284 4962 5318
rect 4996 5284 5006 5318
rect 4952 5268 5006 5284
rect 5048 5319 5102 5335
rect 5048 5285 5058 5319
rect 5092 5285 5102 5319
rect 5048 5269 5102 5285
rect 4608 5237 4662 5253
rect 4608 5203 4618 5237
rect 4652 5203 4662 5237
rect 4608 5187 4662 5203
rect 4715 5237 4779 5253
rect 4715 5203 4735 5237
rect 4769 5203 4779 5237
rect 4620 5127 4650 5187
rect 4715 5172 4779 5203
rect 4704 5142 4922 5172
rect 4704 5127 4734 5142
rect 4892 5127 4922 5142
rect 4976 5127 5006 5268
rect 5060 5127 5090 5269
rect 5144 5230 5174 5409
rect 5234 5341 5264 5409
rect 5333 5341 5363 5363
rect 6036 5341 6066 5363
rect 6135 5349 6165 5409
rect 5216 5325 5270 5341
rect 5216 5291 5226 5325
rect 5260 5291 5270 5325
rect 5216 5275 5270 5291
rect 5312 5325 5366 5341
rect 5312 5291 5322 5325
rect 5356 5291 5366 5325
rect 5312 5275 5366 5291
rect 6036 5325 6090 5341
rect 6036 5291 6046 5325
rect 6080 5291 6090 5325
rect 6036 5275 6090 5291
rect 6135 5333 6189 5349
rect 6135 5299 6145 5333
rect 6179 5299 6189 5333
rect 6135 5283 6189 5299
rect 5138 5214 5192 5230
rect 5138 5180 5148 5214
rect 5182 5180 5192 5214
rect 5138 5164 5192 5180
rect 5144 5127 5174 5164
rect 5234 5127 5264 5275
rect 5333 5243 5363 5275
rect 6036 5243 6066 5275
rect 6135 5127 6165 5283
rect 6231 5237 6261 5409
rect 6207 5221 6261 5237
rect 6207 5187 6217 5221
rect 6251 5187 6261 5221
rect 6207 5171 6261 5187
rect 6231 5127 6261 5171
rect 6303 5237 6333 5409
rect 6399 5365 6429 5409
rect 6488 5365 6518 5409
rect 6572 5394 6602 5409
rect 6375 5349 6429 5365
rect 6375 5315 6385 5349
rect 6419 5315 6429 5349
rect 6375 5299 6429 5315
rect 6475 5349 6529 5365
rect 6475 5315 6485 5349
rect 6519 5315 6529 5349
rect 6475 5299 6529 5315
rect 6571 5364 6602 5394
rect 6656 5394 6686 5409
rect 6844 5394 6874 5409
rect 6656 5364 6874 5394
rect 6303 5221 6357 5237
rect 6303 5187 6313 5221
rect 6347 5187 6357 5221
rect 6303 5171 6357 5187
rect 6303 5127 6333 5171
rect 6399 5127 6429 5299
rect 6488 5127 6518 5299
rect 6571 5253 6601 5364
rect 6656 5349 6697 5364
rect 6667 5253 6697 5349
rect 6928 5334 6958 5409
rect 7012 5335 7042 5409
rect 6904 5318 6958 5334
rect 6904 5284 6914 5318
rect 6948 5284 6958 5318
rect 6904 5268 6958 5284
rect 7000 5319 7054 5335
rect 7000 5285 7010 5319
rect 7044 5285 7054 5319
rect 7000 5269 7054 5285
rect 6560 5237 6614 5253
rect 6560 5203 6570 5237
rect 6604 5203 6614 5237
rect 6560 5187 6614 5203
rect 6667 5237 6731 5253
rect 6667 5203 6687 5237
rect 6721 5203 6731 5237
rect 6572 5127 6602 5187
rect 6667 5172 6731 5203
rect 6656 5142 6874 5172
rect 6656 5127 6686 5142
rect 6844 5127 6874 5142
rect 6928 5127 6958 5268
rect 7012 5127 7042 5269
rect 7096 5230 7126 5409
rect 7186 5341 7216 5409
rect 7285 5341 7315 5363
rect 8038 5347 8068 5369
rect 8137 5355 8167 5415
rect 7168 5325 7222 5341
rect 7168 5291 7178 5325
rect 7212 5291 7222 5325
rect 7168 5275 7222 5291
rect 7264 5325 7318 5341
rect 7264 5291 7274 5325
rect 7308 5291 7318 5325
rect 7264 5275 7318 5291
rect 8038 5331 8092 5347
rect 8038 5297 8048 5331
rect 8082 5297 8092 5331
rect 8038 5281 8092 5297
rect 8137 5339 8191 5355
rect 8137 5305 8147 5339
rect 8181 5305 8191 5339
rect 8137 5289 8191 5305
rect 7090 5214 7144 5230
rect 7090 5180 7100 5214
rect 7134 5180 7144 5214
rect 7090 5164 7144 5180
rect 7096 5127 7126 5164
rect 7186 5127 7216 5275
rect 7285 5243 7315 5275
rect 8038 5249 8068 5281
rect 8137 5133 8167 5289
rect 8233 5243 8263 5415
rect 8209 5227 8263 5243
rect 8209 5193 8219 5227
rect 8253 5193 8263 5227
rect 8209 5177 8263 5193
rect 8233 5133 8263 5177
rect 8305 5243 8335 5415
rect 8401 5371 8431 5415
rect 8490 5371 8520 5415
rect 8574 5400 8604 5415
rect 8377 5355 8431 5371
rect 8377 5321 8387 5355
rect 8421 5321 8431 5355
rect 8377 5305 8431 5321
rect 8477 5355 8531 5371
rect 8477 5321 8487 5355
rect 8521 5321 8531 5355
rect 8477 5305 8531 5321
rect 8573 5370 8604 5400
rect 8658 5400 8688 5415
rect 8846 5400 8876 5415
rect 8658 5370 8876 5400
rect 8305 5227 8359 5243
rect 8305 5193 8315 5227
rect 8349 5193 8359 5227
rect 8305 5177 8359 5193
rect 8305 5133 8335 5177
rect 8401 5133 8431 5305
rect 8490 5133 8520 5305
rect 8573 5259 8603 5370
rect 8658 5355 8699 5370
rect 8669 5259 8699 5355
rect 8930 5340 8960 5415
rect 9014 5341 9044 5415
rect 8906 5324 8960 5340
rect 8906 5290 8916 5324
rect 8950 5290 8960 5324
rect 8906 5274 8960 5290
rect 9002 5325 9056 5341
rect 9002 5291 9012 5325
rect 9046 5291 9056 5325
rect 9002 5275 9056 5291
rect 8562 5243 8616 5259
rect 8562 5209 8572 5243
rect 8606 5209 8616 5243
rect 8562 5193 8616 5209
rect 8669 5243 8733 5259
rect 8669 5209 8689 5243
rect 8723 5209 8733 5243
rect 8574 5133 8604 5193
rect 8669 5178 8733 5209
rect 8658 5148 8876 5178
rect 8658 5133 8688 5148
rect 8846 5133 8876 5148
rect 8930 5133 8960 5274
rect 9014 5133 9044 5275
rect 9098 5236 9128 5415
rect 9188 5347 9218 5415
rect 10231 5555 10261 5711
rect 10327 5665 10357 5837
rect 10303 5649 10357 5665
rect 10303 5615 10313 5649
rect 10347 5615 10357 5649
rect 10303 5599 10357 5615
rect 10327 5555 10357 5599
rect 10399 5665 10429 5837
rect 10495 5793 10525 5837
rect 10584 5793 10614 5837
rect 10668 5822 10698 5837
rect 10471 5777 10525 5793
rect 10471 5743 10481 5777
rect 10515 5743 10525 5777
rect 10471 5727 10525 5743
rect 10571 5777 10625 5793
rect 10571 5743 10581 5777
rect 10615 5743 10625 5777
rect 10571 5727 10625 5743
rect 10667 5792 10698 5822
rect 10752 5822 10782 5837
rect 10940 5822 10970 5837
rect 10752 5792 10970 5822
rect 10399 5649 10453 5665
rect 10399 5615 10409 5649
rect 10443 5615 10453 5649
rect 10399 5599 10453 5615
rect 10399 5555 10429 5599
rect 10495 5555 10525 5727
rect 10584 5555 10614 5727
rect 10667 5681 10697 5792
rect 10752 5777 10793 5792
rect 10763 5681 10793 5777
rect 11024 5762 11054 5837
rect 11108 5763 11138 5837
rect 11000 5746 11054 5762
rect 11000 5712 11010 5746
rect 11044 5712 11054 5746
rect 11000 5696 11054 5712
rect 11096 5747 11150 5763
rect 11096 5713 11106 5747
rect 11140 5713 11150 5747
rect 11096 5697 11150 5713
rect 10656 5665 10710 5681
rect 10656 5631 10666 5665
rect 10700 5631 10710 5665
rect 10656 5615 10710 5631
rect 10763 5665 10827 5681
rect 10763 5631 10783 5665
rect 10817 5631 10827 5665
rect 10668 5555 10698 5615
rect 10763 5600 10827 5631
rect 10752 5570 10970 5600
rect 10752 5555 10782 5570
rect 10940 5555 10970 5570
rect 11024 5555 11054 5696
rect 11108 5555 11138 5697
rect 11192 5658 11222 5837
rect 11282 5769 11312 5837
rect 12194 5909 12224 5935
rect 12293 5909 12323 5935
rect 12389 5909 12419 5935
rect 12461 5909 12491 5935
rect 12557 5909 12587 5935
rect 12646 5909 12676 5935
rect 12730 5909 12760 5935
rect 12814 5909 12844 5935
rect 13002 5909 13032 5935
rect 13086 5909 13116 5935
rect 13170 5909 13200 5935
rect 13254 5909 13284 5935
rect 13344 5909 13374 5935
rect 13443 5909 13473 5935
rect 14152 5917 14182 5943
rect 14251 5917 14281 5943
rect 14347 5917 14377 5943
rect 14419 5917 14449 5943
rect 14515 5917 14545 5943
rect 14604 5917 14634 5943
rect 14688 5917 14718 5943
rect 14772 5917 14802 5943
rect 14960 5917 14990 5943
rect 15044 5917 15074 5943
rect 15128 5917 15158 5943
rect 15212 5917 15242 5943
rect 15302 5917 15332 5943
rect 15401 5917 15431 5943
rect 16146 5923 16176 5949
rect 16245 5923 16275 5949
rect 16341 5923 16371 5949
rect 16413 5923 16443 5949
rect 16509 5923 16539 5949
rect 16598 5923 16628 5949
rect 16682 5923 16712 5949
rect 16766 5923 16796 5949
rect 16954 5923 16984 5949
rect 17038 5923 17068 5949
rect 17122 5923 17152 5949
rect 17206 5923 17236 5949
rect 17296 5923 17326 5949
rect 17395 5923 17425 5949
rect 11381 5769 11411 5791
rect 11264 5753 11318 5769
rect 11264 5719 11274 5753
rect 11308 5719 11318 5753
rect 11264 5703 11318 5719
rect 11360 5753 11414 5769
rect 11360 5719 11370 5753
rect 11404 5719 11414 5753
rect 11360 5703 11414 5719
rect 12194 5757 12224 5779
rect 12293 5765 12323 5825
rect 12194 5741 12248 5757
rect 12194 5707 12204 5741
rect 12238 5707 12248 5741
rect 11186 5642 11240 5658
rect 11186 5608 11196 5642
rect 11230 5608 11240 5642
rect 11186 5592 11240 5608
rect 11192 5555 11222 5592
rect 11282 5555 11312 5703
rect 11381 5671 11411 5703
rect 12194 5691 12248 5707
rect 12293 5749 12347 5765
rect 12293 5715 12303 5749
rect 12337 5715 12347 5749
rect 12293 5699 12347 5715
rect 12194 5659 12224 5691
rect 10132 5445 10162 5471
rect 10231 5445 10261 5471
rect 10327 5445 10357 5471
rect 10399 5445 10429 5471
rect 10495 5445 10525 5471
rect 10584 5445 10614 5471
rect 10668 5445 10698 5471
rect 10752 5445 10782 5471
rect 10940 5445 10970 5471
rect 11024 5445 11054 5471
rect 11108 5445 11138 5471
rect 11192 5445 11222 5471
rect 11282 5445 11312 5471
rect 11381 5445 11411 5471
rect 12293 5543 12323 5699
rect 12389 5653 12419 5825
rect 12365 5637 12419 5653
rect 12365 5603 12375 5637
rect 12409 5603 12419 5637
rect 12365 5587 12419 5603
rect 12389 5543 12419 5587
rect 12461 5653 12491 5825
rect 12557 5781 12587 5825
rect 12646 5781 12676 5825
rect 12730 5810 12760 5825
rect 12533 5765 12587 5781
rect 12533 5731 12543 5765
rect 12577 5731 12587 5765
rect 12533 5715 12587 5731
rect 12633 5765 12687 5781
rect 12633 5731 12643 5765
rect 12677 5731 12687 5765
rect 12633 5715 12687 5731
rect 12729 5780 12760 5810
rect 12814 5810 12844 5825
rect 13002 5810 13032 5825
rect 12814 5780 13032 5810
rect 12461 5637 12515 5653
rect 12461 5603 12471 5637
rect 12505 5603 12515 5637
rect 12461 5587 12515 5603
rect 12461 5543 12491 5587
rect 12557 5543 12587 5715
rect 12646 5543 12676 5715
rect 12729 5669 12759 5780
rect 12814 5765 12855 5780
rect 12825 5669 12855 5765
rect 13086 5750 13116 5825
rect 13170 5751 13200 5825
rect 13062 5734 13116 5750
rect 13062 5700 13072 5734
rect 13106 5700 13116 5734
rect 13062 5684 13116 5700
rect 13158 5735 13212 5751
rect 13158 5701 13168 5735
rect 13202 5701 13212 5735
rect 13158 5685 13212 5701
rect 12718 5653 12772 5669
rect 12718 5619 12728 5653
rect 12762 5619 12772 5653
rect 12718 5603 12772 5619
rect 12825 5653 12889 5669
rect 12825 5619 12845 5653
rect 12879 5619 12889 5653
rect 12730 5543 12760 5603
rect 12825 5588 12889 5619
rect 12814 5558 13032 5588
rect 12814 5543 12844 5558
rect 13002 5543 13032 5558
rect 13086 5543 13116 5684
rect 13170 5543 13200 5685
rect 13254 5646 13284 5825
rect 13344 5757 13374 5825
rect 13443 5757 13473 5779
rect 14152 5765 14182 5787
rect 14251 5773 14281 5833
rect 13326 5741 13380 5757
rect 13326 5707 13336 5741
rect 13370 5707 13380 5741
rect 13326 5691 13380 5707
rect 13422 5741 13476 5757
rect 13422 5707 13432 5741
rect 13466 5707 13476 5741
rect 13422 5691 13476 5707
rect 14152 5749 14206 5765
rect 14152 5715 14162 5749
rect 14196 5715 14206 5749
rect 14152 5699 14206 5715
rect 14251 5757 14305 5773
rect 14251 5723 14261 5757
rect 14295 5723 14305 5757
rect 14251 5707 14305 5723
rect 13248 5630 13302 5646
rect 13248 5596 13258 5630
rect 13292 5596 13302 5630
rect 13248 5580 13302 5596
rect 13254 5543 13284 5580
rect 13344 5543 13374 5691
rect 13443 5659 13473 5691
rect 14152 5667 14182 5699
rect 14251 5551 14281 5707
rect 14347 5661 14377 5833
rect 14323 5645 14377 5661
rect 14323 5611 14333 5645
rect 14367 5611 14377 5645
rect 14323 5595 14377 5611
rect 14347 5551 14377 5595
rect 14419 5661 14449 5833
rect 14515 5789 14545 5833
rect 14604 5789 14634 5833
rect 14688 5818 14718 5833
rect 14491 5773 14545 5789
rect 14491 5739 14501 5773
rect 14535 5739 14545 5773
rect 14491 5723 14545 5739
rect 14591 5773 14645 5789
rect 14591 5739 14601 5773
rect 14635 5739 14645 5773
rect 14591 5723 14645 5739
rect 14687 5788 14718 5818
rect 14772 5818 14802 5833
rect 14960 5818 14990 5833
rect 14772 5788 14990 5818
rect 14419 5645 14473 5661
rect 14419 5611 14429 5645
rect 14463 5611 14473 5645
rect 14419 5595 14473 5611
rect 14419 5551 14449 5595
rect 14515 5551 14545 5723
rect 14604 5551 14634 5723
rect 14687 5677 14717 5788
rect 14772 5773 14813 5788
rect 14783 5677 14813 5773
rect 15044 5758 15074 5833
rect 15128 5759 15158 5833
rect 15020 5742 15074 5758
rect 15020 5708 15030 5742
rect 15064 5708 15074 5742
rect 15020 5692 15074 5708
rect 15116 5743 15170 5759
rect 15116 5709 15126 5743
rect 15160 5709 15170 5743
rect 15116 5693 15170 5709
rect 14676 5661 14730 5677
rect 14676 5627 14686 5661
rect 14720 5627 14730 5661
rect 14676 5611 14730 5627
rect 14783 5661 14847 5677
rect 14783 5627 14803 5661
rect 14837 5627 14847 5661
rect 14688 5551 14718 5611
rect 14783 5596 14847 5627
rect 14772 5566 14990 5596
rect 14772 5551 14802 5566
rect 14960 5551 14990 5566
rect 15044 5551 15074 5692
rect 15128 5551 15158 5693
rect 15212 5654 15242 5833
rect 15302 5765 15332 5833
rect 15401 5765 15431 5787
rect 16146 5771 16176 5793
rect 16245 5779 16275 5839
rect 15284 5749 15338 5765
rect 15284 5715 15294 5749
rect 15328 5715 15338 5749
rect 15284 5699 15338 5715
rect 15380 5749 15434 5765
rect 15380 5715 15390 5749
rect 15424 5715 15434 5749
rect 15380 5699 15434 5715
rect 16146 5755 16200 5771
rect 16146 5721 16156 5755
rect 16190 5721 16200 5755
rect 16146 5705 16200 5721
rect 16245 5763 16299 5779
rect 16245 5729 16255 5763
rect 16289 5729 16299 5763
rect 16245 5713 16299 5729
rect 15206 5638 15260 5654
rect 15206 5604 15216 5638
rect 15250 5604 15260 5638
rect 15206 5588 15260 5604
rect 15212 5551 15242 5588
rect 15302 5551 15332 5699
rect 15401 5667 15431 5699
rect 16146 5673 16176 5705
rect 16245 5557 16275 5713
rect 16341 5667 16371 5839
rect 16317 5651 16371 5667
rect 16317 5617 16327 5651
rect 16361 5617 16371 5651
rect 16317 5601 16371 5617
rect 16341 5557 16371 5601
rect 16413 5667 16443 5839
rect 16509 5795 16539 5839
rect 16598 5795 16628 5839
rect 16682 5824 16712 5839
rect 16485 5779 16539 5795
rect 16485 5745 16495 5779
rect 16529 5745 16539 5779
rect 16485 5729 16539 5745
rect 16585 5779 16639 5795
rect 16585 5745 16595 5779
rect 16629 5745 16639 5779
rect 16585 5729 16639 5745
rect 16681 5794 16712 5824
rect 16766 5824 16796 5839
rect 16954 5824 16984 5839
rect 16766 5794 16984 5824
rect 16413 5651 16467 5667
rect 16413 5617 16423 5651
rect 16457 5617 16467 5651
rect 16413 5601 16467 5617
rect 16413 5557 16443 5601
rect 16509 5557 16539 5729
rect 16598 5557 16628 5729
rect 16681 5683 16711 5794
rect 16766 5779 16807 5794
rect 16777 5683 16807 5779
rect 17038 5764 17068 5839
rect 17122 5765 17152 5839
rect 17014 5748 17068 5764
rect 17014 5714 17024 5748
rect 17058 5714 17068 5748
rect 17014 5698 17068 5714
rect 17110 5749 17164 5765
rect 17110 5715 17120 5749
rect 17154 5715 17164 5749
rect 17110 5699 17164 5715
rect 16670 5667 16724 5683
rect 16670 5633 16680 5667
rect 16714 5633 16724 5667
rect 16670 5617 16724 5633
rect 16777 5667 16841 5683
rect 16777 5633 16797 5667
rect 16831 5633 16841 5667
rect 16682 5557 16712 5617
rect 16777 5602 16841 5633
rect 16766 5572 16984 5602
rect 16766 5557 16796 5572
rect 16954 5557 16984 5572
rect 17038 5557 17068 5698
rect 17122 5557 17152 5699
rect 17206 5660 17236 5839
rect 17296 5771 17326 5839
rect 17395 5771 17425 5793
rect 17278 5755 17332 5771
rect 17278 5721 17288 5755
rect 17322 5721 17332 5755
rect 17278 5705 17332 5721
rect 17374 5755 17428 5771
rect 17374 5721 17384 5755
rect 17418 5721 17428 5755
rect 17374 5705 17428 5721
rect 17200 5644 17254 5660
rect 17200 5610 17210 5644
rect 17244 5610 17254 5644
rect 17200 5594 17254 5610
rect 17206 5557 17236 5594
rect 17296 5557 17326 5705
rect 17395 5673 17425 5705
rect 12194 5433 12224 5459
rect 12293 5433 12323 5459
rect 12389 5433 12419 5459
rect 12461 5433 12491 5459
rect 12557 5433 12587 5459
rect 12646 5433 12676 5459
rect 12730 5433 12760 5459
rect 12814 5433 12844 5459
rect 13002 5433 13032 5459
rect 13086 5433 13116 5459
rect 13170 5433 13200 5459
rect 13254 5433 13284 5459
rect 13344 5433 13374 5459
rect 13443 5433 13473 5459
rect 14152 5441 14182 5467
rect 14251 5441 14281 5467
rect 14347 5441 14377 5467
rect 14419 5441 14449 5467
rect 14515 5441 14545 5467
rect 14604 5441 14634 5467
rect 14688 5441 14718 5467
rect 14772 5441 14802 5467
rect 14960 5441 14990 5467
rect 15044 5441 15074 5467
rect 15128 5441 15158 5467
rect 15212 5441 15242 5467
rect 15302 5441 15332 5467
rect 15401 5441 15431 5467
rect 16146 5447 16176 5473
rect 16245 5447 16275 5473
rect 16341 5447 16371 5473
rect 16413 5447 16443 5473
rect 16509 5447 16539 5473
rect 16598 5447 16628 5473
rect 16682 5447 16712 5473
rect 16766 5447 16796 5473
rect 16954 5447 16984 5473
rect 17038 5447 17068 5473
rect 17122 5447 17152 5473
rect 17206 5447 17236 5473
rect 17296 5447 17326 5473
rect 17395 5447 17425 5473
rect 9287 5347 9317 5369
rect 9170 5331 9224 5347
rect 9170 5297 9180 5331
rect 9214 5297 9224 5331
rect 9170 5281 9224 5297
rect 9266 5331 9320 5347
rect 9266 5297 9276 5331
rect 9310 5297 9320 5331
rect 9266 5281 9320 5297
rect 9092 5220 9146 5236
rect 9092 5186 9102 5220
rect 9136 5186 9146 5220
rect 9092 5170 9146 5186
rect 9098 5133 9128 5170
rect 9188 5133 9218 5281
rect 9287 5249 9317 5281
rect 4084 5017 4114 5043
rect 4183 5017 4213 5043
rect 4279 5017 4309 5043
rect 4351 5017 4381 5043
rect 4447 5017 4477 5043
rect 4536 5017 4566 5043
rect 4620 5017 4650 5043
rect 4704 5017 4734 5043
rect 4892 5017 4922 5043
rect 4976 5017 5006 5043
rect 5060 5017 5090 5043
rect 5144 5017 5174 5043
rect 5234 5017 5264 5043
rect 5333 5017 5363 5043
rect 6036 5017 6066 5043
rect 6135 5017 6165 5043
rect 6231 5017 6261 5043
rect 6303 5017 6333 5043
rect 6399 5017 6429 5043
rect 6488 5017 6518 5043
rect 6572 5017 6602 5043
rect 6656 5017 6686 5043
rect 6844 5017 6874 5043
rect 6928 5017 6958 5043
rect 7012 5017 7042 5043
rect 7096 5017 7126 5043
rect 7186 5017 7216 5043
rect 7285 5017 7315 5043
rect 8038 5023 8068 5049
rect 8137 5023 8167 5049
rect 8233 5023 8263 5049
rect 8305 5023 8335 5049
rect 8401 5023 8431 5049
rect 8490 5023 8520 5049
rect 8574 5023 8604 5049
rect 8658 5023 8688 5049
rect 8846 5023 8876 5049
rect 8930 5023 8960 5049
rect 9014 5023 9044 5049
rect 9098 5023 9128 5049
rect 9188 5023 9218 5049
rect 9287 5023 9317 5049
rect 10160 5047 10190 5073
rect 10259 5047 10289 5073
rect 10355 5047 10385 5073
rect 10427 5047 10457 5073
rect 10523 5047 10553 5073
rect 10612 5047 10642 5073
rect 10696 5047 10726 5073
rect 10780 5047 10810 5073
rect 10968 5047 10998 5073
rect 11052 5047 11082 5073
rect 11136 5047 11166 5073
rect 11220 5047 11250 5073
rect 11310 5047 11340 5073
rect 11409 5047 11439 5073
rect 10160 4895 10190 4917
rect 10259 4903 10289 4963
rect 10160 4879 10214 4895
rect 10160 4845 10170 4879
rect 10204 4845 10214 4879
rect 10160 4829 10214 4845
rect 10259 4887 10313 4903
rect 10259 4853 10269 4887
rect 10303 4853 10313 4887
rect 10259 4837 10313 4853
rect 10160 4797 10190 4829
rect 10259 4681 10289 4837
rect 10355 4791 10385 4963
rect 10331 4775 10385 4791
rect 10331 4741 10341 4775
rect 10375 4741 10385 4775
rect 10331 4725 10385 4741
rect 10355 4681 10385 4725
rect 10427 4791 10457 4963
rect 10523 4919 10553 4963
rect 10612 4919 10642 4963
rect 10696 4948 10726 4963
rect 10499 4903 10553 4919
rect 10499 4869 10509 4903
rect 10543 4869 10553 4903
rect 10499 4853 10553 4869
rect 10599 4903 10653 4919
rect 10599 4869 10609 4903
rect 10643 4869 10653 4903
rect 10599 4853 10653 4869
rect 10695 4918 10726 4948
rect 10780 4948 10810 4963
rect 10968 4948 10998 4963
rect 10780 4918 10998 4948
rect 10427 4775 10481 4791
rect 10427 4741 10437 4775
rect 10471 4741 10481 4775
rect 10427 4725 10481 4741
rect 10427 4681 10457 4725
rect 10523 4681 10553 4853
rect 10612 4681 10642 4853
rect 10695 4807 10725 4918
rect 10780 4903 10821 4918
rect 10791 4807 10821 4903
rect 11052 4888 11082 4963
rect 11136 4889 11166 4963
rect 11028 4872 11082 4888
rect 11028 4838 11038 4872
rect 11072 4838 11082 4872
rect 11028 4822 11082 4838
rect 11124 4873 11178 4889
rect 11124 4839 11134 4873
rect 11168 4839 11178 4873
rect 11124 4823 11178 4839
rect 10684 4791 10738 4807
rect 10684 4757 10694 4791
rect 10728 4757 10738 4791
rect 10684 4741 10738 4757
rect 10791 4791 10855 4807
rect 10791 4757 10811 4791
rect 10845 4757 10855 4791
rect 10696 4681 10726 4741
rect 10791 4726 10855 4757
rect 10780 4696 10998 4726
rect 10780 4681 10810 4696
rect 10968 4681 10998 4696
rect 11052 4681 11082 4822
rect 11136 4681 11166 4823
rect 11220 4784 11250 4963
rect 11310 4895 11340 4963
rect 12430 5003 12460 5029
rect 12529 5003 12559 5029
rect 12625 5003 12655 5029
rect 12697 5003 12727 5029
rect 12793 5003 12823 5029
rect 12882 5003 12912 5029
rect 12966 5003 12996 5029
rect 13050 5003 13080 5029
rect 13238 5003 13268 5029
rect 13322 5003 13352 5029
rect 13406 5003 13436 5029
rect 13490 5003 13520 5029
rect 13580 5003 13610 5029
rect 13679 5003 13709 5029
rect 11409 4895 11439 4917
rect 11292 4879 11346 4895
rect 11292 4845 11302 4879
rect 11336 4845 11346 4879
rect 11292 4829 11346 4845
rect 11388 4879 11442 4895
rect 11388 4845 11398 4879
rect 11432 4845 11442 4879
rect 11388 4829 11442 4845
rect 12430 4851 12460 4873
rect 12529 4859 12559 4919
rect 12430 4835 12484 4851
rect 11214 4768 11268 4784
rect 11214 4734 11224 4768
rect 11258 4734 11268 4768
rect 11214 4718 11268 4734
rect 11220 4681 11250 4718
rect 11310 4681 11340 4829
rect 11409 4797 11439 4829
rect 12430 4801 12440 4835
rect 12474 4801 12484 4835
rect 12430 4785 12484 4801
rect 12529 4843 12583 4859
rect 12529 4809 12539 4843
rect 12573 4809 12583 4843
rect 12529 4793 12583 4809
rect 12430 4753 12460 4785
rect 10160 4571 10190 4597
rect 10259 4571 10289 4597
rect 10355 4571 10385 4597
rect 10427 4571 10457 4597
rect 10523 4571 10553 4597
rect 10612 4571 10642 4597
rect 10696 4571 10726 4597
rect 10780 4571 10810 4597
rect 10968 4571 10998 4597
rect 11052 4571 11082 4597
rect 11136 4571 11166 4597
rect 11220 4571 11250 4597
rect 11310 4571 11340 4597
rect 11409 4571 11439 4597
rect 12529 4637 12559 4793
rect 12625 4747 12655 4919
rect 12601 4731 12655 4747
rect 12601 4697 12611 4731
rect 12645 4697 12655 4731
rect 12601 4681 12655 4697
rect 12625 4637 12655 4681
rect 12697 4747 12727 4919
rect 12793 4875 12823 4919
rect 12882 4875 12912 4919
rect 12966 4904 12996 4919
rect 12769 4859 12823 4875
rect 12769 4825 12779 4859
rect 12813 4825 12823 4859
rect 12769 4809 12823 4825
rect 12869 4859 12923 4875
rect 12869 4825 12879 4859
rect 12913 4825 12923 4859
rect 12869 4809 12923 4825
rect 12965 4874 12996 4904
rect 13050 4904 13080 4919
rect 13238 4904 13268 4919
rect 13050 4874 13268 4904
rect 12697 4731 12751 4747
rect 12697 4697 12707 4731
rect 12741 4697 12751 4731
rect 12697 4681 12751 4697
rect 12697 4637 12727 4681
rect 12793 4637 12823 4809
rect 12882 4637 12912 4809
rect 12965 4763 12995 4874
rect 13050 4859 13091 4874
rect 13061 4763 13091 4859
rect 13322 4844 13352 4919
rect 13406 4845 13436 4919
rect 13298 4828 13352 4844
rect 13298 4794 13308 4828
rect 13342 4794 13352 4828
rect 13298 4778 13352 4794
rect 13394 4829 13448 4845
rect 13394 4795 13404 4829
rect 13438 4795 13448 4829
rect 13394 4779 13448 4795
rect 12954 4747 13008 4763
rect 12954 4713 12964 4747
rect 12998 4713 13008 4747
rect 12954 4697 13008 4713
rect 13061 4747 13125 4763
rect 13061 4713 13081 4747
rect 13115 4713 13125 4747
rect 12966 4637 12996 4697
rect 13061 4682 13125 4713
rect 13050 4652 13268 4682
rect 13050 4637 13080 4652
rect 13238 4637 13268 4652
rect 13322 4637 13352 4778
rect 13406 4637 13436 4779
rect 13490 4740 13520 4919
rect 13580 4851 13610 4919
rect 14432 4997 14462 5023
rect 14531 4997 14561 5023
rect 14627 4997 14657 5023
rect 14699 4997 14729 5023
rect 14795 4997 14825 5023
rect 14884 4997 14914 5023
rect 14968 4997 14998 5023
rect 15052 4997 15082 5023
rect 15240 4997 15270 5023
rect 15324 4997 15354 5023
rect 15408 4997 15438 5023
rect 15492 4997 15522 5023
rect 15582 4997 15612 5023
rect 15681 4997 15711 5023
rect 13679 4851 13709 4873
rect 13562 4835 13616 4851
rect 13562 4801 13572 4835
rect 13606 4801 13616 4835
rect 13562 4785 13616 4801
rect 13658 4835 13712 4851
rect 13658 4801 13668 4835
rect 13702 4801 13712 4835
rect 13658 4785 13712 4801
rect 14432 4845 14462 4867
rect 14531 4853 14561 4913
rect 14432 4829 14486 4845
rect 14432 4795 14442 4829
rect 14476 4795 14486 4829
rect 13484 4724 13538 4740
rect 13484 4690 13494 4724
rect 13528 4690 13538 4724
rect 13484 4674 13538 4690
rect 13490 4637 13520 4674
rect 13580 4637 13610 4785
rect 13679 4753 13709 4785
rect 14432 4779 14486 4795
rect 14531 4837 14585 4853
rect 14531 4803 14541 4837
rect 14575 4803 14585 4837
rect 14531 4787 14585 4803
rect 14432 4747 14462 4779
rect 12430 4527 12460 4553
rect 12529 4527 12559 4553
rect 12625 4527 12655 4553
rect 12697 4527 12727 4553
rect 12793 4527 12823 4553
rect 12882 4527 12912 4553
rect 12966 4527 12996 4553
rect 13050 4527 13080 4553
rect 13238 4527 13268 4553
rect 13322 4527 13352 4553
rect 13406 4527 13436 4553
rect 13490 4527 13520 4553
rect 13580 4527 13610 4553
rect 13679 4527 13709 4553
rect 14531 4631 14561 4787
rect 14627 4741 14657 4913
rect 14603 4725 14657 4741
rect 14603 4691 14613 4725
rect 14647 4691 14657 4725
rect 14603 4675 14657 4691
rect 14627 4631 14657 4675
rect 14699 4741 14729 4913
rect 14795 4869 14825 4913
rect 14884 4869 14914 4913
rect 14968 4898 14998 4913
rect 14771 4853 14825 4869
rect 14771 4819 14781 4853
rect 14815 4819 14825 4853
rect 14771 4803 14825 4819
rect 14871 4853 14925 4869
rect 14871 4819 14881 4853
rect 14915 4819 14925 4853
rect 14871 4803 14925 4819
rect 14967 4868 14998 4898
rect 15052 4898 15082 4913
rect 15240 4898 15270 4913
rect 15052 4868 15270 4898
rect 14699 4725 14753 4741
rect 14699 4691 14709 4725
rect 14743 4691 14753 4725
rect 14699 4675 14753 4691
rect 14699 4631 14729 4675
rect 14795 4631 14825 4803
rect 14884 4631 14914 4803
rect 14967 4757 14997 4868
rect 15052 4853 15093 4868
rect 15063 4757 15093 4853
rect 15324 4838 15354 4913
rect 15408 4839 15438 4913
rect 15300 4822 15354 4838
rect 15300 4788 15310 4822
rect 15344 4788 15354 4822
rect 15300 4772 15354 4788
rect 15396 4823 15450 4839
rect 15396 4789 15406 4823
rect 15440 4789 15450 4823
rect 15396 4773 15450 4789
rect 14956 4741 15010 4757
rect 14956 4707 14966 4741
rect 15000 4707 15010 4741
rect 14956 4691 15010 4707
rect 15063 4741 15127 4757
rect 15063 4707 15083 4741
rect 15117 4707 15127 4741
rect 14968 4631 14998 4691
rect 15063 4676 15127 4707
rect 15052 4646 15270 4676
rect 15052 4631 15082 4646
rect 15240 4631 15270 4646
rect 15324 4631 15354 4772
rect 15408 4631 15438 4773
rect 15492 4734 15522 4913
rect 15582 4845 15612 4913
rect 16454 4979 16484 5005
rect 16553 4979 16583 5005
rect 16649 4979 16679 5005
rect 16721 4979 16751 5005
rect 16817 4979 16847 5005
rect 16906 4979 16936 5005
rect 16990 4979 17020 5005
rect 17074 4979 17104 5005
rect 17262 4979 17292 5005
rect 17346 4979 17376 5005
rect 17430 4979 17460 5005
rect 17514 4979 17544 5005
rect 17604 4979 17634 5005
rect 17703 4979 17733 5005
rect 15681 4845 15711 4867
rect 15564 4829 15618 4845
rect 15564 4795 15574 4829
rect 15608 4795 15618 4829
rect 15564 4779 15618 4795
rect 15660 4829 15714 4845
rect 15660 4795 15670 4829
rect 15704 4795 15714 4829
rect 15660 4779 15714 4795
rect 16454 4827 16484 4849
rect 16553 4835 16583 4895
rect 16454 4811 16508 4827
rect 15486 4718 15540 4734
rect 15486 4684 15496 4718
rect 15530 4684 15540 4718
rect 15486 4668 15540 4684
rect 15492 4631 15522 4668
rect 15582 4631 15612 4779
rect 15681 4747 15711 4779
rect 16454 4777 16464 4811
rect 16498 4777 16508 4811
rect 16454 4761 16508 4777
rect 16553 4819 16607 4835
rect 16553 4785 16563 4819
rect 16597 4785 16607 4819
rect 16553 4769 16607 4785
rect 16454 4729 16484 4761
rect 14432 4521 14462 4547
rect 14531 4521 14561 4547
rect 14627 4521 14657 4547
rect 14699 4521 14729 4547
rect 14795 4521 14825 4547
rect 14884 4521 14914 4547
rect 14968 4521 14998 4547
rect 15052 4521 15082 4547
rect 15240 4521 15270 4547
rect 15324 4521 15354 4547
rect 15408 4521 15438 4547
rect 15492 4521 15522 4547
rect 15582 4521 15612 4547
rect 15681 4521 15711 4547
rect 16553 4613 16583 4769
rect 16649 4723 16679 4895
rect 16625 4707 16679 4723
rect 16625 4673 16635 4707
rect 16669 4673 16679 4707
rect 16625 4657 16679 4673
rect 16649 4613 16679 4657
rect 16721 4723 16751 4895
rect 16817 4851 16847 4895
rect 16906 4851 16936 4895
rect 16990 4880 17020 4895
rect 16793 4835 16847 4851
rect 16793 4801 16803 4835
rect 16837 4801 16847 4835
rect 16793 4785 16847 4801
rect 16893 4835 16947 4851
rect 16893 4801 16903 4835
rect 16937 4801 16947 4835
rect 16893 4785 16947 4801
rect 16989 4850 17020 4880
rect 17074 4880 17104 4895
rect 17262 4880 17292 4895
rect 17074 4850 17292 4880
rect 16721 4707 16775 4723
rect 16721 4673 16731 4707
rect 16765 4673 16775 4707
rect 16721 4657 16775 4673
rect 16721 4613 16751 4657
rect 16817 4613 16847 4785
rect 16906 4613 16936 4785
rect 16989 4739 17019 4850
rect 17074 4835 17115 4850
rect 17085 4739 17115 4835
rect 17346 4820 17376 4895
rect 17430 4821 17460 4895
rect 17322 4804 17376 4820
rect 17322 4770 17332 4804
rect 17366 4770 17376 4804
rect 17322 4754 17376 4770
rect 17418 4805 17472 4821
rect 17418 4771 17428 4805
rect 17462 4771 17472 4805
rect 17418 4755 17472 4771
rect 16978 4723 17032 4739
rect 16978 4689 16988 4723
rect 17022 4689 17032 4723
rect 16978 4673 17032 4689
rect 17085 4723 17149 4739
rect 17085 4689 17105 4723
rect 17139 4689 17149 4723
rect 16990 4613 17020 4673
rect 17085 4658 17149 4689
rect 17074 4628 17292 4658
rect 17074 4613 17104 4628
rect 17262 4613 17292 4628
rect 17346 4613 17376 4754
rect 17430 4613 17460 4755
rect 17514 4716 17544 4895
rect 17604 4827 17634 4895
rect 17703 4827 17733 4849
rect 17586 4811 17640 4827
rect 17586 4777 17596 4811
rect 17630 4777 17640 4811
rect 17586 4761 17640 4777
rect 17682 4811 17736 4827
rect 17682 4777 17692 4811
rect 17726 4777 17736 4811
rect 17682 4761 17736 4777
rect 17508 4700 17562 4716
rect 17508 4666 17518 4700
rect 17552 4666 17562 4700
rect 17508 4650 17562 4666
rect 17514 4613 17544 4650
rect 17604 4613 17634 4761
rect 17703 4729 17733 4761
rect 16454 4503 16484 4529
rect 16553 4503 16583 4529
rect 16649 4503 16679 4529
rect 16721 4503 16751 4529
rect 16817 4503 16847 4529
rect 16906 4503 16936 4529
rect 16990 4503 17020 4529
rect 17074 4503 17104 4529
rect 17262 4503 17292 4529
rect 17346 4503 17376 4529
rect 17430 4503 17460 4529
rect 17514 4503 17544 4529
rect 17604 4503 17634 4529
rect 17703 4503 17733 4529
rect 1920 2241 1950 2267
rect 2019 2241 2049 2267
rect 2115 2241 2145 2267
rect 2187 2241 2217 2267
rect 2283 2241 2313 2267
rect 2372 2241 2402 2267
rect 2456 2241 2486 2267
rect 2540 2241 2570 2267
rect 2728 2241 2758 2267
rect 2812 2241 2842 2267
rect 2896 2241 2926 2267
rect 2980 2241 3010 2267
rect 3070 2241 3100 2267
rect 3169 2241 3199 2267
rect 1920 2089 1950 2111
rect 2019 2097 2049 2157
rect 1920 2073 1974 2089
rect 1920 2039 1930 2073
rect 1964 2039 1974 2073
rect 1920 2023 1974 2039
rect 2019 2081 2073 2097
rect 2019 2047 2029 2081
rect 2063 2047 2073 2081
rect 2019 2031 2073 2047
rect 1920 1991 1950 2023
rect 2019 1875 2049 2031
rect 2115 1985 2145 2157
rect 2091 1969 2145 1985
rect 2091 1935 2101 1969
rect 2135 1935 2145 1969
rect 2091 1919 2145 1935
rect 2115 1875 2145 1919
rect 2187 1985 2217 2157
rect 2283 2113 2313 2157
rect 2372 2113 2402 2157
rect 2456 2142 2486 2157
rect 2259 2097 2313 2113
rect 2259 2063 2269 2097
rect 2303 2063 2313 2097
rect 2259 2047 2313 2063
rect 2359 2097 2413 2113
rect 2359 2063 2369 2097
rect 2403 2063 2413 2097
rect 2359 2047 2413 2063
rect 2455 2112 2486 2142
rect 2540 2142 2570 2157
rect 2728 2142 2758 2157
rect 2540 2112 2758 2142
rect 2187 1969 2241 1985
rect 2187 1935 2197 1969
rect 2231 1935 2241 1969
rect 2187 1919 2241 1935
rect 2187 1875 2217 1919
rect 2283 1875 2313 2047
rect 2372 1875 2402 2047
rect 2455 2001 2485 2112
rect 2540 2097 2581 2112
rect 2551 2001 2581 2097
rect 2812 2082 2842 2157
rect 2896 2083 2926 2157
rect 2788 2066 2842 2082
rect 2788 2032 2798 2066
rect 2832 2032 2842 2066
rect 2788 2016 2842 2032
rect 2884 2067 2938 2083
rect 2884 2033 2894 2067
rect 2928 2033 2938 2067
rect 2884 2017 2938 2033
rect 2444 1985 2498 2001
rect 2444 1951 2454 1985
rect 2488 1951 2498 1985
rect 2444 1935 2498 1951
rect 2551 1985 2615 2001
rect 2551 1951 2571 1985
rect 2605 1951 2615 1985
rect 2456 1875 2486 1935
rect 2551 1920 2615 1951
rect 2540 1890 2758 1920
rect 2540 1875 2570 1890
rect 2728 1875 2758 1890
rect 2812 1875 2842 2016
rect 2896 1875 2926 2017
rect 2980 1978 3010 2157
rect 3070 2089 3100 2157
rect 3990 2237 4020 2263
rect 4089 2237 4119 2263
rect 4185 2237 4215 2263
rect 4257 2237 4287 2263
rect 4353 2237 4383 2263
rect 4442 2237 4472 2263
rect 4526 2237 4556 2263
rect 4610 2237 4640 2263
rect 4798 2237 4828 2263
rect 4882 2237 4912 2263
rect 4966 2237 4996 2263
rect 5050 2237 5080 2263
rect 5140 2237 5170 2263
rect 5239 2237 5269 2263
rect 5942 2237 5972 2263
rect 6041 2237 6071 2263
rect 6137 2237 6167 2263
rect 6209 2237 6239 2263
rect 6305 2237 6335 2263
rect 6394 2237 6424 2263
rect 6478 2237 6508 2263
rect 6562 2237 6592 2263
rect 6750 2237 6780 2263
rect 6834 2237 6864 2263
rect 6918 2237 6948 2263
rect 7002 2237 7032 2263
rect 7092 2237 7122 2263
rect 7191 2237 7221 2263
rect 7944 2243 7974 2269
rect 8043 2243 8073 2269
rect 8139 2243 8169 2269
rect 8211 2243 8241 2269
rect 8307 2243 8337 2269
rect 8396 2243 8426 2269
rect 8480 2243 8510 2269
rect 8564 2243 8594 2269
rect 8752 2243 8782 2269
rect 8836 2243 8866 2269
rect 8920 2243 8950 2269
rect 9004 2243 9034 2269
rect 9094 2243 9124 2269
rect 9193 2243 9223 2269
rect 9896 2243 9926 2269
rect 9995 2243 10025 2269
rect 10091 2243 10121 2269
rect 10163 2243 10193 2269
rect 10259 2243 10289 2269
rect 10348 2243 10378 2269
rect 10432 2243 10462 2269
rect 10516 2243 10546 2269
rect 10704 2243 10734 2269
rect 10788 2243 10818 2269
rect 10872 2243 10902 2269
rect 10956 2243 10986 2269
rect 11046 2243 11076 2269
rect 11145 2243 11175 2269
rect 11888 2243 11918 2269
rect 11987 2243 12017 2269
rect 12083 2243 12113 2269
rect 12155 2243 12185 2269
rect 12251 2243 12281 2269
rect 12340 2243 12370 2269
rect 12424 2243 12454 2269
rect 12508 2243 12538 2269
rect 12696 2243 12726 2269
rect 12780 2243 12810 2269
rect 12864 2243 12894 2269
rect 12948 2243 12978 2269
rect 13038 2243 13068 2269
rect 13137 2243 13167 2269
rect 13840 2243 13870 2269
rect 13939 2243 13969 2269
rect 14035 2243 14065 2269
rect 14107 2243 14137 2269
rect 14203 2243 14233 2269
rect 14292 2243 14322 2269
rect 14376 2243 14406 2269
rect 14460 2243 14490 2269
rect 14648 2243 14678 2269
rect 14732 2243 14762 2269
rect 14816 2243 14846 2269
rect 14900 2243 14930 2269
rect 14990 2243 15020 2269
rect 15089 2243 15119 2269
rect 15904 2243 15934 2269
rect 16003 2243 16033 2269
rect 16099 2243 16129 2269
rect 16171 2243 16201 2269
rect 16267 2243 16297 2269
rect 16356 2243 16386 2269
rect 16440 2243 16470 2269
rect 16524 2243 16554 2269
rect 16712 2243 16742 2269
rect 16796 2243 16826 2269
rect 16880 2243 16910 2269
rect 16964 2243 16994 2269
rect 17054 2243 17084 2269
rect 17153 2243 17183 2269
rect 3169 2089 3199 2111
rect 3052 2073 3106 2089
rect 3052 2039 3062 2073
rect 3096 2039 3106 2073
rect 3052 2023 3106 2039
rect 3148 2073 3202 2089
rect 3148 2039 3158 2073
rect 3192 2039 3202 2073
rect 3148 2023 3202 2039
rect 3990 2085 4020 2107
rect 4089 2093 4119 2153
rect 3990 2069 4044 2085
rect 3990 2035 4000 2069
rect 4034 2035 4044 2069
rect 2974 1962 3028 1978
rect 2974 1928 2984 1962
rect 3018 1928 3028 1962
rect 2974 1912 3028 1928
rect 2980 1875 3010 1912
rect 3070 1875 3100 2023
rect 3169 1991 3199 2023
rect 3990 2019 4044 2035
rect 4089 2077 4143 2093
rect 4089 2043 4099 2077
rect 4133 2043 4143 2077
rect 4089 2027 4143 2043
rect 3990 1987 4020 2019
rect 1920 1765 1950 1791
rect 2019 1765 2049 1791
rect 2115 1765 2145 1791
rect 2187 1765 2217 1791
rect 2283 1765 2313 1791
rect 2372 1765 2402 1791
rect 2456 1765 2486 1791
rect 2540 1765 2570 1791
rect 2728 1765 2758 1791
rect 2812 1765 2842 1791
rect 2896 1765 2926 1791
rect 2980 1765 3010 1791
rect 3070 1765 3100 1791
rect 3169 1765 3199 1791
rect 4089 1871 4119 2027
rect 4185 1981 4215 2153
rect 4161 1965 4215 1981
rect 4161 1931 4171 1965
rect 4205 1931 4215 1965
rect 4161 1915 4215 1931
rect 4185 1871 4215 1915
rect 4257 1981 4287 2153
rect 4353 2109 4383 2153
rect 4442 2109 4472 2153
rect 4526 2138 4556 2153
rect 4329 2093 4383 2109
rect 4329 2059 4339 2093
rect 4373 2059 4383 2093
rect 4329 2043 4383 2059
rect 4429 2093 4483 2109
rect 4429 2059 4439 2093
rect 4473 2059 4483 2093
rect 4429 2043 4483 2059
rect 4525 2108 4556 2138
rect 4610 2138 4640 2153
rect 4798 2138 4828 2153
rect 4610 2108 4828 2138
rect 4257 1965 4311 1981
rect 4257 1931 4267 1965
rect 4301 1931 4311 1965
rect 4257 1915 4311 1931
rect 4257 1871 4287 1915
rect 4353 1871 4383 2043
rect 4442 1871 4472 2043
rect 4525 1997 4555 2108
rect 4610 2093 4651 2108
rect 4621 1997 4651 2093
rect 4882 2078 4912 2153
rect 4966 2079 4996 2153
rect 4858 2062 4912 2078
rect 4858 2028 4868 2062
rect 4902 2028 4912 2062
rect 4858 2012 4912 2028
rect 4954 2063 5008 2079
rect 4954 2029 4964 2063
rect 4998 2029 5008 2063
rect 4954 2013 5008 2029
rect 4514 1981 4568 1997
rect 4514 1947 4524 1981
rect 4558 1947 4568 1981
rect 4514 1931 4568 1947
rect 4621 1981 4685 1997
rect 4621 1947 4641 1981
rect 4675 1947 4685 1981
rect 4526 1871 4556 1931
rect 4621 1916 4685 1947
rect 4610 1886 4828 1916
rect 4610 1871 4640 1886
rect 4798 1871 4828 1886
rect 4882 1871 4912 2012
rect 4966 1871 4996 2013
rect 5050 1974 5080 2153
rect 5140 2085 5170 2153
rect 5239 2085 5269 2107
rect 5942 2085 5972 2107
rect 6041 2093 6071 2153
rect 5122 2069 5176 2085
rect 5122 2035 5132 2069
rect 5166 2035 5176 2069
rect 5122 2019 5176 2035
rect 5218 2069 5272 2085
rect 5218 2035 5228 2069
rect 5262 2035 5272 2069
rect 5218 2019 5272 2035
rect 5942 2069 5996 2085
rect 5942 2035 5952 2069
rect 5986 2035 5996 2069
rect 5942 2019 5996 2035
rect 6041 2077 6095 2093
rect 6041 2043 6051 2077
rect 6085 2043 6095 2077
rect 6041 2027 6095 2043
rect 5044 1958 5098 1974
rect 5044 1924 5054 1958
rect 5088 1924 5098 1958
rect 5044 1908 5098 1924
rect 5050 1871 5080 1908
rect 5140 1871 5170 2019
rect 5239 1987 5269 2019
rect 5942 1987 5972 2019
rect 6041 1871 6071 2027
rect 6137 1981 6167 2153
rect 6113 1965 6167 1981
rect 6113 1931 6123 1965
rect 6157 1931 6167 1965
rect 6113 1915 6167 1931
rect 6137 1871 6167 1915
rect 6209 1981 6239 2153
rect 6305 2109 6335 2153
rect 6394 2109 6424 2153
rect 6478 2138 6508 2153
rect 6281 2093 6335 2109
rect 6281 2059 6291 2093
rect 6325 2059 6335 2093
rect 6281 2043 6335 2059
rect 6381 2093 6435 2109
rect 6381 2059 6391 2093
rect 6425 2059 6435 2093
rect 6381 2043 6435 2059
rect 6477 2108 6508 2138
rect 6562 2138 6592 2153
rect 6750 2138 6780 2153
rect 6562 2108 6780 2138
rect 6209 1965 6263 1981
rect 6209 1931 6219 1965
rect 6253 1931 6263 1965
rect 6209 1915 6263 1931
rect 6209 1871 6239 1915
rect 6305 1871 6335 2043
rect 6394 1871 6424 2043
rect 6477 1997 6507 2108
rect 6562 2093 6603 2108
rect 6573 1997 6603 2093
rect 6834 2078 6864 2153
rect 6918 2079 6948 2153
rect 6810 2062 6864 2078
rect 6810 2028 6820 2062
rect 6854 2028 6864 2062
rect 6810 2012 6864 2028
rect 6906 2063 6960 2079
rect 6906 2029 6916 2063
rect 6950 2029 6960 2063
rect 6906 2013 6960 2029
rect 6466 1981 6520 1997
rect 6466 1947 6476 1981
rect 6510 1947 6520 1981
rect 6466 1931 6520 1947
rect 6573 1981 6637 1997
rect 6573 1947 6593 1981
rect 6627 1947 6637 1981
rect 6478 1871 6508 1931
rect 6573 1916 6637 1947
rect 6562 1886 6780 1916
rect 6562 1871 6592 1886
rect 6750 1871 6780 1886
rect 6834 1871 6864 2012
rect 6918 1871 6948 2013
rect 7002 1974 7032 2153
rect 7092 2085 7122 2153
rect 7191 2085 7221 2107
rect 7944 2091 7974 2113
rect 8043 2099 8073 2159
rect 7074 2069 7128 2085
rect 7074 2035 7084 2069
rect 7118 2035 7128 2069
rect 7074 2019 7128 2035
rect 7170 2069 7224 2085
rect 7170 2035 7180 2069
rect 7214 2035 7224 2069
rect 7170 2019 7224 2035
rect 7944 2075 7998 2091
rect 7944 2041 7954 2075
rect 7988 2041 7998 2075
rect 7944 2025 7998 2041
rect 8043 2083 8097 2099
rect 8043 2049 8053 2083
rect 8087 2049 8097 2083
rect 8043 2033 8097 2049
rect 6996 1958 7050 1974
rect 6996 1924 7006 1958
rect 7040 1924 7050 1958
rect 6996 1908 7050 1924
rect 7002 1871 7032 1908
rect 7092 1871 7122 2019
rect 7191 1987 7221 2019
rect 7944 1993 7974 2025
rect 8043 1877 8073 2033
rect 8139 1987 8169 2159
rect 8115 1971 8169 1987
rect 8115 1937 8125 1971
rect 8159 1937 8169 1971
rect 8115 1921 8169 1937
rect 8139 1877 8169 1921
rect 8211 1987 8241 2159
rect 8307 2115 8337 2159
rect 8396 2115 8426 2159
rect 8480 2144 8510 2159
rect 8283 2099 8337 2115
rect 8283 2065 8293 2099
rect 8327 2065 8337 2099
rect 8283 2049 8337 2065
rect 8383 2099 8437 2115
rect 8383 2065 8393 2099
rect 8427 2065 8437 2099
rect 8383 2049 8437 2065
rect 8479 2114 8510 2144
rect 8564 2144 8594 2159
rect 8752 2144 8782 2159
rect 8564 2114 8782 2144
rect 8211 1971 8265 1987
rect 8211 1937 8221 1971
rect 8255 1937 8265 1971
rect 8211 1921 8265 1937
rect 8211 1877 8241 1921
rect 8307 1877 8337 2049
rect 8396 1877 8426 2049
rect 8479 2003 8509 2114
rect 8564 2099 8605 2114
rect 8575 2003 8605 2099
rect 8836 2084 8866 2159
rect 8920 2085 8950 2159
rect 8812 2068 8866 2084
rect 8812 2034 8822 2068
rect 8856 2034 8866 2068
rect 8812 2018 8866 2034
rect 8908 2069 8962 2085
rect 8908 2035 8918 2069
rect 8952 2035 8962 2069
rect 8908 2019 8962 2035
rect 8468 1987 8522 2003
rect 8468 1953 8478 1987
rect 8512 1953 8522 1987
rect 8468 1937 8522 1953
rect 8575 1987 8639 2003
rect 8575 1953 8595 1987
rect 8629 1953 8639 1987
rect 8480 1877 8510 1937
rect 8575 1922 8639 1953
rect 8564 1892 8782 1922
rect 8564 1877 8594 1892
rect 8752 1877 8782 1892
rect 8836 1877 8866 2018
rect 8920 1877 8950 2019
rect 9004 1980 9034 2159
rect 9094 2091 9124 2159
rect 9193 2091 9223 2113
rect 9896 2091 9926 2113
rect 9995 2099 10025 2159
rect 9076 2075 9130 2091
rect 9076 2041 9086 2075
rect 9120 2041 9130 2075
rect 9076 2025 9130 2041
rect 9172 2075 9226 2091
rect 9172 2041 9182 2075
rect 9216 2041 9226 2075
rect 9172 2025 9226 2041
rect 9896 2075 9950 2091
rect 9896 2041 9906 2075
rect 9940 2041 9950 2075
rect 9896 2025 9950 2041
rect 9995 2083 10049 2099
rect 9995 2049 10005 2083
rect 10039 2049 10049 2083
rect 9995 2033 10049 2049
rect 8998 1964 9052 1980
rect 8998 1930 9008 1964
rect 9042 1930 9052 1964
rect 8998 1914 9052 1930
rect 9004 1877 9034 1914
rect 9094 1877 9124 2025
rect 9193 1993 9223 2025
rect 9896 1993 9926 2025
rect 9995 1877 10025 2033
rect 10091 1987 10121 2159
rect 10067 1971 10121 1987
rect 10067 1937 10077 1971
rect 10111 1937 10121 1971
rect 10067 1921 10121 1937
rect 10091 1877 10121 1921
rect 10163 1987 10193 2159
rect 10259 2115 10289 2159
rect 10348 2115 10378 2159
rect 10432 2144 10462 2159
rect 10235 2099 10289 2115
rect 10235 2065 10245 2099
rect 10279 2065 10289 2099
rect 10235 2049 10289 2065
rect 10335 2099 10389 2115
rect 10335 2065 10345 2099
rect 10379 2065 10389 2099
rect 10335 2049 10389 2065
rect 10431 2114 10462 2144
rect 10516 2144 10546 2159
rect 10704 2144 10734 2159
rect 10516 2114 10734 2144
rect 10163 1971 10217 1987
rect 10163 1937 10173 1971
rect 10207 1937 10217 1971
rect 10163 1921 10217 1937
rect 10163 1877 10193 1921
rect 10259 1877 10289 2049
rect 10348 1877 10378 2049
rect 10431 2003 10461 2114
rect 10516 2099 10557 2114
rect 10527 2003 10557 2099
rect 10788 2084 10818 2159
rect 10872 2085 10902 2159
rect 10764 2068 10818 2084
rect 10764 2034 10774 2068
rect 10808 2034 10818 2068
rect 10764 2018 10818 2034
rect 10860 2069 10914 2085
rect 10860 2035 10870 2069
rect 10904 2035 10914 2069
rect 10860 2019 10914 2035
rect 10420 1987 10474 2003
rect 10420 1953 10430 1987
rect 10464 1953 10474 1987
rect 10420 1937 10474 1953
rect 10527 1987 10591 2003
rect 10527 1953 10547 1987
rect 10581 1953 10591 1987
rect 10432 1877 10462 1937
rect 10527 1922 10591 1953
rect 10516 1892 10734 1922
rect 10516 1877 10546 1892
rect 10704 1877 10734 1892
rect 10788 1877 10818 2018
rect 10872 1877 10902 2019
rect 10956 1980 10986 2159
rect 11046 2091 11076 2159
rect 11145 2091 11175 2113
rect 11888 2091 11918 2113
rect 11987 2099 12017 2159
rect 11028 2075 11082 2091
rect 11028 2041 11038 2075
rect 11072 2041 11082 2075
rect 11028 2025 11082 2041
rect 11124 2075 11178 2091
rect 11124 2041 11134 2075
rect 11168 2041 11178 2075
rect 11124 2025 11178 2041
rect 11888 2075 11942 2091
rect 11888 2041 11898 2075
rect 11932 2041 11942 2075
rect 11888 2025 11942 2041
rect 11987 2083 12041 2099
rect 11987 2049 11997 2083
rect 12031 2049 12041 2083
rect 11987 2033 12041 2049
rect 10950 1964 11004 1980
rect 10950 1930 10960 1964
rect 10994 1930 11004 1964
rect 10950 1914 11004 1930
rect 10956 1877 10986 1914
rect 11046 1877 11076 2025
rect 11145 1993 11175 2025
rect 11888 1993 11918 2025
rect 11987 1877 12017 2033
rect 12083 1987 12113 2159
rect 12059 1971 12113 1987
rect 12059 1937 12069 1971
rect 12103 1937 12113 1971
rect 12059 1921 12113 1937
rect 12083 1877 12113 1921
rect 12155 1987 12185 2159
rect 12251 2115 12281 2159
rect 12340 2115 12370 2159
rect 12424 2144 12454 2159
rect 12227 2099 12281 2115
rect 12227 2065 12237 2099
rect 12271 2065 12281 2099
rect 12227 2049 12281 2065
rect 12327 2099 12381 2115
rect 12327 2065 12337 2099
rect 12371 2065 12381 2099
rect 12327 2049 12381 2065
rect 12423 2114 12454 2144
rect 12508 2144 12538 2159
rect 12696 2144 12726 2159
rect 12508 2114 12726 2144
rect 12155 1971 12209 1987
rect 12155 1937 12165 1971
rect 12199 1937 12209 1971
rect 12155 1921 12209 1937
rect 12155 1877 12185 1921
rect 12251 1877 12281 2049
rect 12340 1877 12370 2049
rect 12423 2003 12453 2114
rect 12508 2099 12549 2114
rect 12519 2003 12549 2099
rect 12780 2084 12810 2159
rect 12864 2085 12894 2159
rect 12756 2068 12810 2084
rect 12756 2034 12766 2068
rect 12800 2034 12810 2068
rect 12756 2018 12810 2034
rect 12852 2069 12906 2085
rect 12852 2035 12862 2069
rect 12896 2035 12906 2069
rect 12852 2019 12906 2035
rect 12412 1987 12466 2003
rect 12412 1953 12422 1987
rect 12456 1953 12466 1987
rect 12412 1937 12466 1953
rect 12519 1987 12583 2003
rect 12519 1953 12539 1987
rect 12573 1953 12583 1987
rect 12424 1877 12454 1937
rect 12519 1922 12583 1953
rect 12508 1892 12726 1922
rect 12508 1877 12538 1892
rect 12696 1877 12726 1892
rect 12780 1877 12810 2018
rect 12864 1877 12894 2019
rect 12948 1980 12978 2159
rect 13038 2091 13068 2159
rect 13137 2091 13167 2113
rect 13840 2091 13870 2113
rect 13939 2099 13969 2159
rect 13020 2075 13074 2091
rect 13020 2041 13030 2075
rect 13064 2041 13074 2075
rect 13020 2025 13074 2041
rect 13116 2075 13170 2091
rect 13116 2041 13126 2075
rect 13160 2041 13170 2075
rect 13116 2025 13170 2041
rect 13840 2075 13894 2091
rect 13840 2041 13850 2075
rect 13884 2041 13894 2075
rect 13840 2025 13894 2041
rect 13939 2083 13993 2099
rect 13939 2049 13949 2083
rect 13983 2049 13993 2083
rect 13939 2033 13993 2049
rect 12942 1964 12996 1980
rect 12942 1930 12952 1964
rect 12986 1930 12996 1964
rect 12942 1914 12996 1930
rect 12948 1877 12978 1914
rect 13038 1877 13068 2025
rect 13137 1993 13167 2025
rect 13840 1993 13870 2025
rect 13939 1877 13969 2033
rect 14035 1987 14065 2159
rect 14011 1971 14065 1987
rect 14011 1937 14021 1971
rect 14055 1937 14065 1971
rect 14011 1921 14065 1937
rect 14035 1877 14065 1921
rect 14107 1987 14137 2159
rect 14203 2115 14233 2159
rect 14292 2115 14322 2159
rect 14376 2144 14406 2159
rect 14179 2099 14233 2115
rect 14179 2065 14189 2099
rect 14223 2065 14233 2099
rect 14179 2049 14233 2065
rect 14279 2099 14333 2115
rect 14279 2065 14289 2099
rect 14323 2065 14333 2099
rect 14279 2049 14333 2065
rect 14375 2114 14406 2144
rect 14460 2144 14490 2159
rect 14648 2144 14678 2159
rect 14460 2114 14678 2144
rect 14107 1971 14161 1987
rect 14107 1937 14117 1971
rect 14151 1937 14161 1971
rect 14107 1921 14161 1937
rect 14107 1877 14137 1921
rect 14203 1877 14233 2049
rect 14292 1877 14322 2049
rect 14375 2003 14405 2114
rect 14460 2099 14501 2114
rect 14471 2003 14501 2099
rect 14732 2084 14762 2159
rect 14816 2085 14846 2159
rect 14708 2068 14762 2084
rect 14708 2034 14718 2068
rect 14752 2034 14762 2068
rect 14708 2018 14762 2034
rect 14804 2069 14858 2085
rect 14804 2035 14814 2069
rect 14848 2035 14858 2069
rect 14804 2019 14858 2035
rect 14364 1987 14418 2003
rect 14364 1953 14374 1987
rect 14408 1953 14418 1987
rect 14364 1937 14418 1953
rect 14471 1987 14535 2003
rect 14471 1953 14491 1987
rect 14525 1953 14535 1987
rect 14376 1877 14406 1937
rect 14471 1922 14535 1953
rect 14460 1892 14678 1922
rect 14460 1877 14490 1892
rect 14648 1877 14678 1892
rect 14732 1877 14762 2018
rect 14816 1877 14846 2019
rect 14900 1980 14930 2159
rect 14990 2091 15020 2159
rect 15089 2091 15119 2113
rect 15904 2091 15934 2113
rect 16003 2099 16033 2159
rect 14972 2075 15026 2091
rect 14972 2041 14982 2075
rect 15016 2041 15026 2075
rect 14972 2025 15026 2041
rect 15068 2075 15122 2091
rect 15068 2041 15078 2075
rect 15112 2041 15122 2075
rect 15068 2025 15122 2041
rect 15904 2075 15958 2091
rect 15904 2041 15914 2075
rect 15948 2041 15958 2075
rect 15904 2025 15958 2041
rect 16003 2083 16057 2099
rect 16003 2049 16013 2083
rect 16047 2049 16057 2083
rect 16003 2033 16057 2049
rect 14894 1964 14948 1980
rect 14894 1930 14904 1964
rect 14938 1930 14948 1964
rect 14894 1914 14948 1930
rect 14900 1877 14930 1914
rect 14990 1877 15020 2025
rect 15089 1993 15119 2025
rect 15904 1993 15934 2025
rect 16003 1877 16033 2033
rect 16099 1987 16129 2159
rect 16075 1971 16129 1987
rect 16075 1937 16085 1971
rect 16119 1937 16129 1971
rect 16075 1921 16129 1937
rect 16099 1877 16129 1921
rect 16171 1987 16201 2159
rect 16267 2115 16297 2159
rect 16356 2115 16386 2159
rect 16440 2144 16470 2159
rect 16243 2099 16297 2115
rect 16243 2065 16253 2099
rect 16287 2065 16297 2099
rect 16243 2049 16297 2065
rect 16343 2099 16397 2115
rect 16343 2065 16353 2099
rect 16387 2065 16397 2099
rect 16343 2049 16397 2065
rect 16439 2114 16470 2144
rect 16524 2144 16554 2159
rect 16712 2144 16742 2159
rect 16524 2114 16742 2144
rect 16171 1971 16225 1987
rect 16171 1937 16181 1971
rect 16215 1937 16225 1971
rect 16171 1921 16225 1937
rect 16171 1877 16201 1921
rect 16267 1877 16297 2049
rect 16356 1877 16386 2049
rect 16439 2003 16469 2114
rect 16524 2099 16565 2114
rect 16535 2003 16565 2099
rect 16796 2084 16826 2159
rect 16880 2085 16910 2159
rect 16772 2068 16826 2084
rect 16772 2034 16782 2068
rect 16816 2034 16826 2068
rect 16772 2018 16826 2034
rect 16868 2069 16922 2085
rect 16868 2035 16878 2069
rect 16912 2035 16922 2069
rect 16868 2019 16922 2035
rect 16428 1987 16482 2003
rect 16428 1953 16438 1987
rect 16472 1953 16482 1987
rect 16428 1937 16482 1953
rect 16535 1987 16599 2003
rect 16535 1953 16555 1987
rect 16589 1953 16599 1987
rect 16440 1877 16470 1937
rect 16535 1922 16599 1953
rect 16524 1892 16742 1922
rect 16524 1877 16554 1892
rect 16712 1877 16742 1892
rect 16796 1877 16826 2018
rect 16880 1877 16910 2019
rect 16964 1980 16994 2159
rect 17054 2091 17084 2159
rect 17153 2091 17183 2113
rect 17036 2075 17090 2091
rect 17036 2041 17046 2075
rect 17080 2041 17090 2075
rect 17036 2025 17090 2041
rect 17132 2075 17186 2091
rect 17132 2041 17142 2075
rect 17176 2041 17186 2075
rect 17132 2025 17186 2041
rect 16958 1964 17012 1980
rect 16958 1930 16968 1964
rect 17002 1930 17012 1964
rect 16958 1914 17012 1930
rect 16964 1877 16994 1914
rect 17054 1877 17084 2025
rect 17153 1993 17183 2025
rect 3990 1761 4020 1787
rect 4089 1761 4119 1787
rect 4185 1761 4215 1787
rect 4257 1761 4287 1787
rect 4353 1761 4383 1787
rect 4442 1761 4472 1787
rect 4526 1761 4556 1787
rect 4610 1761 4640 1787
rect 4798 1761 4828 1787
rect 4882 1761 4912 1787
rect 4966 1761 4996 1787
rect 5050 1761 5080 1787
rect 5140 1761 5170 1787
rect 5239 1761 5269 1787
rect 5942 1761 5972 1787
rect 6041 1761 6071 1787
rect 6137 1761 6167 1787
rect 6209 1761 6239 1787
rect 6305 1761 6335 1787
rect 6394 1761 6424 1787
rect 6478 1761 6508 1787
rect 6562 1761 6592 1787
rect 6750 1761 6780 1787
rect 6834 1761 6864 1787
rect 6918 1761 6948 1787
rect 7002 1761 7032 1787
rect 7092 1761 7122 1787
rect 7191 1761 7221 1787
rect 7944 1767 7974 1793
rect 8043 1767 8073 1793
rect 8139 1767 8169 1793
rect 8211 1767 8241 1793
rect 8307 1767 8337 1793
rect 8396 1767 8426 1793
rect 8480 1767 8510 1793
rect 8564 1767 8594 1793
rect 8752 1767 8782 1793
rect 8836 1767 8866 1793
rect 8920 1767 8950 1793
rect 9004 1767 9034 1793
rect 9094 1767 9124 1793
rect 9193 1767 9223 1793
rect 9896 1767 9926 1793
rect 9995 1767 10025 1793
rect 10091 1767 10121 1793
rect 10163 1767 10193 1793
rect 10259 1767 10289 1793
rect 10348 1767 10378 1793
rect 10432 1767 10462 1793
rect 10516 1767 10546 1793
rect 10704 1767 10734 1793
rect 10788 1767 10818 1793
rect 10872 1767 10902 1793
rect 10956 1767 10986 1793
rect 11046 1767 11076 1793
rect 11145 1767 11175 1793
rect 11888 1767 11918 1793
rect 11987 1767 12017 1793
rect 12083 1767 12113 1793
rect 12155 1767 12185 1793
rect 12251 1767 12281 1793
rect 12340 1767 12370 1793
rect 12424 1767 12454 1793
rect 12508 1767 12538 1793
rect 12696 1767 12726 1793
rect 12780 1767 12810 1793
rect 12864 1767 12894 1793
rect 12948 1767 12978 1793
rect 13038 1767 13068 1793
rect 13137 1767 13167 1793
rect 13840 1767 13870 1793
rect 13939 1767 13969 1793
rect 14035 1767 14065 1793
rect 14107 1767 14137 1793
rect 14203 1767 14233 1793
rect 14292 1767 14322 1793
rect 14376 1767 14406 1793
rect 14460 1767 14490 1793
rect 14648 1767 14678 1793
rect 14732 1767 14762 1793
rect 14816 1767 14846 1793
rect 14900 1767 14930 1793
rect 14990 1767 15020 1793
rect 15089 1767 15119 1793
rect 15904 1767 15934 1793
rect 16003 1767 16033 1793
rect 16099 1767 16129 1793
rect 16171 1767 16201 1793
rect 16267 1767 16297 1793
rect 16356 1767 16386 1793
rect 16440 1767 16470 1793
rect 16524 1767 16554 1793
rect 16712 1767 16742 1793
rect 16796 1767 16826 1793
rect 16880 1767 16910 1793
rect 16964 1767 16994 1793
rect 17054 1767 17084 1793
rect 17153 1767 17183 1793
<< polycont >>
rect 9419 16261 9453 16295
rect 9536 16261 9570 16295
rect 9671 16261 9705 16295
rect 9767 16261 9801 16295
rect 9506 15517 9540 15551
rect 9647 15517 9681 15551
rect 9755 15517 9789 15551
rect 11505 15407 11539 15441
rect 11651 15407 11685 15441
rect 11757 15407 11791 15441
rect 11853 15407 11887 15441
rect 11964 15407 11998 15441
rect 10690 14907 10724 14941
rect 10831 14907 10865 14941
rect 10939 14907 10973 14941
rect 9429 14697 9463 14731
rect 9546 14697 9580 14731
rect 9681 14697 9715 14731
rect 9777 14697 9811 14731
rect 9516 13953 9550 13987
rect 9657 13953 9691 13987
rect 12845 14149 12879 14183
rect 9765 13953 9799 13987
rect 10721 13941 10755 13975
rect 10867 13941 10901 13975
rect 10973 13941 11007 13975
rect 11069 13941 11103 13975
rect 11180 13941 11214 13975
rect 12623 13925 12657 13959
rect 12749 13925 12783 13959
rect 12925 13925 12959 13959
rect 13021 13925 13055 13959
rect 11726 13567 11760 13601
rect 11862 13567 11896 13601
rect 11965 13567 11999 13601
rect 10987 13326 11021 13360
rect 9421 13029 9455 13063
rect 9538 13029 9572 13063
rect 9673 13029 9707 13063
rect 9769 13029 9803 13063
rect 10849 13053 10883 13087
rect 11059 13093 11093 13127
rect 11155 13099 11189 13133
rect 9508 12285 9542 12319
rect 9649 12285 9683 12319
rect 9757 12285 9791 12319
rect 10884 12079 10918 12113
rect 11025 12079 11059 12113
rect 11133 12079 11167 12113
rect 9431 11465 9465 11499
rect 9548 11465 9582 11499
rect 9683 11465 9717 11499
rect 9779 11465 9813 11499
rect 9518 10721 9552 10755
rect 9659 10721 9693 10755
rect 9767 10721 9801 10755
rect 6274 6351 6308 6385
rect 10142 5719 10176 5753
rect 10241 5727 10275 5761
rect 1960 5299 1994 5333
rect 2059 5307 2093 5341
rect 2131 5195 2165 5229
rect 2299 5323 2333 5357
rect 2399 5323 2433 5357
rect 2227 5195 2261 5229
rect 2828 5292 2862 5326
rect 2924 5293 2958 5327
rect 2484 5211 2518 5245
rect 2601 5211 2635 5245
rect 3092 5299 3126 5333
rect 3188 5299 3222 5333
rect 4094 5291 4128 5325
rect 3014 5188 3048 5222
rect 4193 5299 4227 5333
rect 4265 5187 4299 5221
rect 4433 5315 4467 5349
rect 4533 5315 4567 5349
rect 4361 5187 4395 5221
rect 4962 5284 4996 5318
rect 5058 5285 5092 5319
rect 4618 5203 4652 5237
rect 4735 5203 4769 5237
rect 5226 5291 5260 5325
rect 5322 5291 5356 5325
rect 6046 5291 6080 5325
rect 6145 5299 6179 5333
rect 5148 5180 5182 5214
rect 6217 5187 6251 5221
rect 6385 5315 6419 5349
rect 6485 5315 6519 5349
rect 6313 5187 6347 5221
rect 6914 5284 6948 5318
rect 7010 5285 7044 5319
rect 6570 5203 6604 5237
rect 6687 5203 6721 5237
rect 7178 5291 7212 5325
rect 7274 5291 7308 5325
rect 8048 5297 8082 5331
rect 8147 5305 8181 5339
rect 7100 5180 7134 5214
rect 8219 5193 8253 5227
rect 8387 5321 8421 5355
rect 8487 5321 8521 5355
rect 8315 5193 8349 5227
rect 8916 5290 8950 5324
rect 9012 5291 9046 5325
rect 8572 5209 8606 5243
rect 8689 5209 8723 5243
rect 10313 5615 10347 5649
rect 10481 5743 10515 5777
rect 10581 5743 10615 5777
rect 10409 5615 10443 5649
rect 11010 5712 11044 5746
rect 11106 5713 11140 5747
rect 10666 5631 10700 5665
rect 10783 5631 10817 5665
rect 11274 5719 11308 5753
rect 11370 5719 11404 5753
rect 12204 5707 12238 5741
rect 11196 5608 11230 5642
rect 12303 5715 12337 5749
rect 12375 5603 12409 5637
rect 12543 5731 12577 5765
rect 12643 5731 12677 5765
rect 12471 5603 12505 5637
rect 13072 5700 13106 5734
rect 13168 5701 13202 5735
rect 12728 5619 12762 5653
rect 12845 5619 12879 5653
rect 13336 5707 13370 5741
rect 13432 5707 13466 5741
rect 14162 5715 14196 5749
rect 14261 5723 14295 5757
rect 13258 5596 13292 5630
rect 14333 5611 14367 5645
rect 14501 5739 14535 5773
rect 14601 5739 14635 5773
rect 14429 5611 14463 5645
rect 15030 5708 15064 5742
rect 15126 5709 15160 5743
rect 14686 5627 14720 5661
rect 14803 5627 14837 5661
rect 15294 5715 15328 5749
rect 15390 5715 15424 5749
rect 16156 5721 16190 5755
rect 16255 5729 16289 5763
rect 15216 5604 15250 5638
rect 16327 5617 16361 5651
rect 16495 5745 16529 5779
rect 16595 5745 16629 5779
rect 16423 5617 16457 5651
rect 17024 5714 17058 5748
rect 17120 5715 17154 5749
rect 16680 5633 16714 5667
rect 16797 5633 16831 5667
rect 17288 5721 17322 5755
rect 17384 5721 17418 5755
rect 17210 5610 17244 5644
rect 9180 5297 9214 5331
rect 9276 5297 9310 5331
rect 9102 5186 9136 5220
rect 10170 4845 10204 4879
rect 10269 4853 10303 4887
rect 10341 4741 10375 4775
rect 10509 4869 10543 4903
rect 10609 4869 10643 4903
rect 10437 4741 10471 4775
rect 11038 4838 11072 4872
rect 11134 4839 11168 4873
rect 10694 4757 10728 4791
rect 10811 4757 10845 4791
rect 11302 4845 11336 4879
rect 11398 4845 11432 4879
rect 11224 4734 11258 4768
rect 12440 4801 12474 4835
rect 12539 4809 12573 4843
rect 12611 4697 12645 4731
rect 12779 4825 12813 4859
rect 12879 4825 12913 4859
rect 12707 4697 12741 4731
rect 13308 4794 13342 4828
rect 13404 4795 13438 4829
rect 12964 4713 12998 4747
rect 13081 4713 13115 4747
rect 13572 4801 13606 4835
rect 13668 4801 13702 4835
rect 14442 4795 14476 4829
rect 13494 4690 13528 4724
rect 14541 4803 14575 4837
rect 14613 4691 14647 4725
rect 14781 4819 14815 4853
rect 14881 4819 14915 4853
rect 14709 4691 14743 4725
rect 15310 4788 15344 4822
rect 15406 4789 15440 4823
rect 14966 4707 15000 4741
rect 15083 4707 15117 4741
rect 15574 4795 15608 4829
rect 15670 4795 15704 4829
rect 15496 4684 15530 4718
rect 16464 4777 16498 4811
rect 16563 4785 16597 4819
rect 16635 4673 16669 4707
rect 16803 4801 16837 4835
rect 16903 4801 16937 4835
rect 16731 4673 16765 4707
rect 17332 4770 17366 4804
rect 17428 4771 17462 4805
rect 16988 4689 17022 4723
rect 17105 4689 17139 4723
rect 17596 4777 17630 4811
rect 17692 4777 17726 4811
rect 17518 4666 17552 4700
rect 1930 2039 1964 2073
rect 2029 2047 2063 2081
rect 2101 1935 2135 1969
rect 2269 2063 2303 2097
rect 2369 2063 2403 2097
rect 2197 1935 2231 1969
rect 2798 2032 2832 2066
rect 2894 2033 2928 2067
rect 2454 1951 2488 1985
rect 2571 1951 2605 1985
rect 3062 2039 3096 2073
rect 3158 2039 3192 2073
rect 4000 2035 4034 2069
rect 2984 1928 3018 1962
rect 4099 2043 4133 2077
rect 4171 1931 4205 1965
rect 4339 2059 4373 2093
rect 4439 2059 4473 2093
rect 4267 1931 4301 1965
rect 4868 2028 4902 2062
rect 4964 2029 4998 2063
rect 4524 1947 4558 1981
rect 4641 1947 4675 1981
rect 5132 2035 5166 2069
rect 5228 2035 5262 2069
rect 5952 2035 5986 2069
rect 6051 2043 6085 2077
rect 5054 1924 5088 1958
rect 6123 1931 6157 1965
rect 6291 2059 6325 2093
rect 6391 2059 6425 2093
rect 6219 1931 6253 1965
rect 6820 2028 6854 2062
rect 6916 2029 6950 2063
rect 6476 1947 6510 1981
rect 6593 1947 6627 1981
rect 7084 2035 7118 2069
rect 7180 2035 7214 2069
rect 7954 2041 7988 2075
rect 8053 2049 8087 2083
rect 7006 1924 7040 1958
rect 8125 1937 8159 1971
rect 8293 2065 8327 2099
rect 8393 2065 8427 2099
rect 8221 1937 8255 1971
rect 8822 2034 8856 2068
rect 8918 2035 8952 2069
rect 8478 1953 8512 1987
rect 8595 1953 8629 1987
rect 9086 2041 9120 2075
rect 9182 2041 9216 2075
rect 9906 2041 9940 2075
rect 10005 2049 10039 2083
rect 9008 1930 9042 1964
rect 10077 1937 10111 1971
rect 10245 2065 10279 2099
rect 10345 2065 10379 2099
rect 10173 1937 10207 1971
rect 10774 2034 10808 2068
rect 10870 2035 10904 2069
rect 10430 1953 10464 1987
rect 10547 1953 10581 1987
rect 11038 2041 11072 2075
rect 11134 2041 11168 2075
rect 11898 2041 11932 2075
rect 11997 2049 12031 2083
rect 10960 1930 10994 1964
rect 12069 1937 12103 1971
rect 12237 2065 12271 2099
rect 12337 2065 12371 2099
rect 12165 1937 12199 1971
rect 12766 2034 12800 2068
rect 12862 2035 12896 2069
rect 12422 1953 12456 1987
rect 12539 1953 12573 1987
rect 13030 2041 13064 2075
rect 13126 2041 13160 2075
rect 13850 2041 13884 2075
rect 13949 2049 13983 2083
rect 12952 1930 12986 1964
rect 14021 1937 14055 1971
rect 14189 2065 14223 2099
rect 14289 2065 14323 2099
rect 14117 1937 14151 1971
rect 14718 2034 14752 2068
rect 14814 2035 14848 2069
rect 14374 1953 14408 1987
rect 14491 1953 14525 1987
rect 14982 2041 15016 2075
rect 15078 2041 15112 2075
rect 15914 2041 15948 2075
rect 16013 2049 16047 2083
rect 14904 1930 14938 1964
rect 16085 1937 16119 1971
rect 16253 2065 16287 2099
rect 16353 2065 16387 2099
rect 16181 1937 16215 1971
rect 16782 2034 16816 2068
rect 16878 2035 16912 2069
rect 16438 1953 16472 1987
rect 16555 1953 16589 1987
rect 17046 2041 17080 2075
rect 17142 2041 17176 2075
rect 16968 1930 17002 1964
<< locali >>
rect 9334 16573 9363 16607
rect 9397 16573 9455 16607
rect 9489 16573 9547 16607
rect 9581 16573 9639 16607
rect 9673 16573 9731 16607
rect 9765 16573 9823 16607
rect 9857 16573 9915 16607
rect 9949 16573 9978 16607
rect 9351 16531 9427 16539
rect 9351 16497 9377 16531
rect 9411 16497 9427 16531
rect 9351 16463 9427 16497
rect 9351 16429 9377 16463
rect 9411 16429 9427 16463
rect 9351 16403 9427 16429
rect 9545 16521 9579 16573
rect 9545 16453 9579 16487
rect 9545 16403 9579 16419
rect 9613 16521 9679 16539
rect 9613 16487 9629 16521
rect 9663 16487 9679 16521
rect 9613 16453 9679 16487
rect 9713 16521 9747 16573
rect 9713 16471 9747 16487
rect 9781 16521 9861 16539
rect 9781 16487 9817 16521
rect 9851 16487 9861 16521
rect 9613 16419 9629 16453
rect 9663 16437 9679 16453
rect 9781 16453 9861 16487
rect 9781 16437 9817 16453
rect 9663 16419 9817 16437
rect 9851 16419 9861 16453
rect 9613 16403 9861 16419
rect 9897 16523 9961 16539
rect 9897 16489 9901 16523
rect 9935 16489 9961 16523
rect 9897 16455 9961 16489
rect 9897 16421 9901 16455
rect 9935 16421 9961 16455
rect 9351 16211 9385 16403
rect 9897 16394 9961 16421
rect 9897 16387 9910 16394
rect 9419 16335 9680 16369
rect 9897 16353 9901 16387
rect 9944 16356 9961 16394
rect 9935 16353 9961 16356
rect 9419 16296 9468 16335
rect 9419 16295 9420 16296
rect 9454 16262 9468 16296
rect 9453 16261 9468 16262
rect 9502 16298 9612 16301
rect 9502 16295 9540 16298
rect 9502 16261 9536 16295
rect 9574 16264 9612 16298
rect 9570 16261 9612 16264
rect 9646 16295 9680 16335
rect 9835 16319 9961 16353
rect 9755 16295 9801 16311
rect 9646 16261 9671 16295
rect 9705 16261 9721 16295
rect 9755 16261 9767 16295
rect 9419 16245 9468 16261
rect 9755 16211 9801 16261
rect 9351 16177 9801 16211
rect 9461 16163 9495 16177
rect 9361 16107 9377 16141
rect 9411 16107 9427 16141
rect 9835 16143 9869 16319
rect 9461 16113 9495 16129
rect 9361 16063 9427 16107
rect 9529 16107 9545 16141
rect 9579 16107 9595 16141
rect 9678 16109 9713 16143
rect 9747 16109 9813 16143
rect 9847 16109 9869 16143
rect 9903 16214 9961 16230
rect 9937 16180 9961 16214
rect 9903 16146 9961 16180
rect 9937 16112 9961 16146
rect 9529 16063 9595 16107
rect 9903 16063 9961 16112
rect 9334 16029 9363 16063
rect 9397 16029 9455 16063
rect 9489 16029 9547 16063
rect 9581 16029 9639 16063
rect 9673 16029 9731 16063
rect 9765 16029 9823 16063
rect 9857 16029 9915 16063
rect 9949 16029 9978 16063
rect 9432 15829 9461 15863
rect 9495 15829 9553 15863
rect 9587 15829 9645 15863
rect 9679 15829 9737 15863
rect 9771 15829 9829 15863
rect 9863 15829 9892 15863
rect 9489 15745 9545 15829
rect 9679 15787 9745 15829
rect 9489 15711 9503 15745
rect 9537 15711 9545 15745
rect 9489 15695 9545 15711
rect 9579 15745 9639 15761
rect 9579 15711 9587 15745
rect 9621 15711 9639 15745
rect 9579 15651 9639 15711
rect 9679 15753 9695 15787
rect 9729 15753 9745 15787
rect 9679 15719 9745 15753
rect 9679 15685 9695 15719
rect 9729 15685 9745 15719
rect 9783 15787 9875 15795
rect 9783 15753 9799 15787
rect 9833 15753 9875 15787
rect 9783 15719 9875 15753
rect 11474 15719 11503 15753
rect 11537 15719 11595 15753
rect 11629 15719 11687 15753
rect 11721 15719 11779 15753
rect 11813 15719 11871 15753
rect 11905 15719 11963 15753
rect 11997 15719 12055 15753
rect 12089 15719 12118 15753
rect 9783 15685 9799 15719
rect 9833 15685 9875 15719
rect 9452 15574 9505 15639
rect 9579 15617 9767 15651
rect 9452 15534 9454 15574
rect 9496 15567 9505 15574
rect 9733 15567 9767 15617
rect 9496 15551 9587 15567
rect 9496 15534 9506 15551
rect 9452 15517 9506 15534
rect 9540 15517 9587 15551
rect 9631 15564 9699 15567
rect 9631 15524 9644 15564
rect 9686 15524 9699 15564
rect 9631 15517 9647 15524
rect 9681 15517 9699 15524
rect 9733 15551 9791 15567
rect 9733 15517 9755 15551
rect 9789 15517 9791 15551
rect 9733 15501 9791 15517
rect 9733 15483 9767 15501
rect 9489 15445 9767 15483
rect 9825 15494 9875 15685
rect 11492 15677 11559 15719
rect 11492 15643 11509 15677
rect 11543 15643 11559 15677
rect 11593 15669 11643 15685
rect 11593 15635 11601 15669
rect 11635 15635 11643 15669
rect 9825 15460 9836 15494
rect 9872 15460 9875 15494
rect 9489 15423 9555 15445
rect 9489 15389 9503 15423
rect 9537 15389 9555 15423
rect 9825 15411 9875 15460
rect 9489 15373 9555 15389
rect 9679 15395 9729 15411
rect 9679 15361 9695 15395
rect 9679 15319 9729 15361
rect 9763 15395 9875 15411
rect 9763 15361 9779 15395
rect 9813 15361 9875 15395
rect 9763 15353 9875 15361
rect 11491 15441 11539 15607
rect 11593 15525 11643 15635
rect 11687 15677 11753 15719
rect 11687 15643 11703 15677
rect 11737 15643 11753 15677
rect 11687 15575 11753 15643
rect 11790 15669 11840 15685
rect 11790 15635 11798 15669
rect 11832 15635 11840 15669
rect 11790 15525 11840 15635
rect 11933 15677 11999 15719
rect 11933 15643 11949 15677
rect 11983 15643 11999 15677
rect 11933 15609 11999 15643
rect 12033 15677 12101 15685
rect 12033 15643 12049 15677
rect 12083 15643 12101 15677
rect 12033 15633 12101 15643
rect 11933 15575 11949 15609
rect 11983 15575 11999 15609
rect 11933 15559 11999 15575
rect 12049 15609 12101 15633
rect 12083 15575 12101 15609
rect 12049 15541 12101 15575
rect 11491 15407 11505 15441
rect 11491 15404 11539 15407
rect 11491 15368 11498 15404
rect 11534 15368 11539 15404
rect 11491 15345 11539 15368
rect 11573 15491 12011 15525
rect 9432 15285 9461 15319
rect 9495 15285 9553 15319
rect 9587 15285 9645 15319
rect 9679 15285 9737 15319
rect 9771 15285 9829 15319
rect 9863 15285 9892 15319
rect 11573 15309 11607 15491
rect 11948 15457 12011 15491
rect 12083 15507 12101 15541
rect 11508 15293 11607 15309
rect 11508 15259 11509 15293
rect 11543 15259 11607 15293
rect 11651 15441 11721 15457
rect 11685 15438 11721 15441
rect 11651 15402 11670 15407
rect 11704 15402 11721 15438
rect 11651 15264 11721 15402
rect 11757 15441 11817 15457
rect 11791 15407 11817 15441
rect 11757 15314 11817 15407
rect 11757 15280 11768 15314
rect 11802 15280 11817 15314
rect 11757 15263 11817 15280
rect 11853 15441 11909 15457
rect 11887 15407 11909 15441
rect 11948 15441 12014 15457
rect 11948 15407 11964 15441
rect 11998 15407 12014 15441
rect 12049 15436 12101 15507
rect 11853 15384 11909 15407
rect 11853 15348 11864 15384
rect 11898 15348 11909 15384
rect 12049 15402 12056 15436
rect 12090 15402 12101 15436
rect 11853 15263 11909 15348
rect 11945 15353 11999 15369
rect 12049 15353 12101 15402
rect 11945 15319 11950 15353
rect 11984 15319 11999 15353
rect 11945 15285 11999 15319
rect 10616 15219 10645 15253
rect 10679 15219 10737 15253
rect 10771 15219 10829 15253
rect 10863 15219 10921 15253
rect 10955 15219 11013 15253
rect 11047 15219 11076 15253
rect 11508 15243 11607 15259
rect 11945 15251 11950 15285
rect 11984 15251 11999 15285
rect 12033 15319 12049 15353
rect 12083 15319 12101 15353
rect 12033 15285 12101 15319
rect 12033 15251 12049 15285
rect 12083 15251 12101 15285
rect 10673 15135 10729 15219
rect 10863 15177 10929 15219
rect 11945 15209 11999 15251
rect 10673 15101 10687 15135
rect 10721 15101 10729 15135
rect 10673 15085 10729 15101
rect 10763 15135 10823 15151
rect 10763 15101 10771 15135
rect 10805 15101 10823 15135
rect 9344 15009 9373 15043
rect 9407 15009 9465 15043
rect 9499 15009 9557 15043
rect 9591 15009 9649 15043
rect 9683 15009 9741 15043
rect 9775 15009 9833 15043
rect 9867 15009 9925 15043
rect 9959 15009 9988 15043
rect 10763 15041 10823 15101
rect 10863 15143 10879 15177
rect 10913 15143 10929 15177
rect 10863 15109 10929 15143
rect 10863 15075 10879 15109
rect 10913 15075 10929 15109
rect 10967 15177 11059 15185
rect 10967 15143 10983 15177
rect 11017 15152 11059 15177
rect 11474 15175 11503 15209
rect 11537 15175 11595 15209
rect 11629 15175 11687 15209
rect 11721 15175 11779 15209
rect 11813 15175 11871 15209
rect 11905 15175 11963 15209
rect 11997 15175 12055 15209
rect 12089 15175 12118 15209
rect 10967 15116 11010 15143
rect 11050 15116 11059 15152
rect 10967 15109 11059 15116
rect 10967 15075 10983 15109
rect 11017 15075 11059 15109
rect 9361 14967 9437 14975
rect 9361 14933 9387 14967
rect 9421 14933 9437 14967
rect 9361 14899 9437 14933
rect 9361 14865 9387 14899
rect 9421 14865 9437 14899
rect 9361 14839 9437 14865
rect 9555 14957 9589 15009
rect 9555 14889 9589 14923
rect 9555 14839 9589 14855
rect 9623 14957 9689 14975
rect 9623 14923 9639 14957
rect 9673 14923 9689 14957
rect 9623 14889 9689 14923
rect 9723 14957 9757 15009
rect 9723 14907 9757 14923
rect 9791 14957 9871 14975
rect 9791 14923 9827 14957
rect 9861 14923 9871 14957
rect 9623 14855 9639 14889
rect 9673 14873 9689 14889
rect 9791 14889 9871 14923
rect 9791 14873 9827 14889
rect 9673 14855 9827 14873
rect 9861 14855 9871 14889
rect 9623 14839 9871 14855
rect 9907 14959 9971 14975
rect 9907 14925 9911 14959
rect 9945 14934 9971 14959
rect 9907 14900 9922 14925
rect 9956 14900 9971 14934
rect 10636 14957 10689 15029
rect 10763 15007 10951 15041
rect 10917 14957 10951 15007
rect 10636 14942 10771 14957
rect 10636 14907 10690 14942
rect 10724 14907 10771 14942
rect 10815 14942 10883 14957
rect 10815 14908 10830 14942
rect 10866 14908 10883 14942
rect 10815 14907 10831 14908
rect 10865 14907 10883 14908
rect 10917 14941 10975 14957
rect 10917 14907 10939 14941
rect 10973 14907 10975 14941
rect 9907 14891 9971 14900
rect 9907 14857 9911 14891
rect 9945 14857 9971 14891
rect 10917 14891 10975 14907
rect 10917 14873 10951 14891
rect 9361 14647 9395 14839
rect 9907 14823 9971 14857
rect 9429 14771 9690 14805
rect 9907 14789 9911 14823
rect 9945 14789 9971 14823
rect 9429 14732 9478 14771
rect 9429 14731 9430 14732
rect 9464 14698 9478 14732
rect 9463 14697 9478 14698
rect 9512 14734 9622 14737
rect 9512 14731 9550 14734
rect 9512 14697 9546 14731
rect 9584 14700 9622 14734
rect 9580 14697 9622 14700
rect 9656 14731 9690 14771
rect 9845 14755 9971 14789
rect 10673 14835 10951 14873
rect 10673 14813 10739 14835
rect 10673 14779 10687 14813
rect 10721 14779 10739 14813
rect 11009 14801 11059 15075
rect 10673 14763 10739 14779
rect 10863 14785 10913 14801
rect 9765 14731 9811 14747
rect 9656 14697 9681 14731
rect 9715 14697 9731 14731
rect 9765 14697 9777 14731
rect 9429 14681 9478 14697
rect 9765 14647 9811 14697
rect 9361 14613 9811 14647
rect 9471 14599 9505 14613
rect 9371 14543 9387 14577
rect 9421 14543 9437 14577
rect 9845 14579 9879 14755
rect 10863 14751 10879 14785
rect 10863 14709 10913 14751
rect 10947 14785 11059 14801
rect 10947 14751 10963 14785
rect 10997 14751 11059 14785
rect 10947 14743 11059 14751
rect 10616 14675 10645 14709
rect 10679 14675 10737 14709
rect 10771 14675 10829 14709
rect 10863 14675 10921 14709
rect 10955 14675 11013 14709
rect 11047 14675 11076 14709
rect 9471 14549 9505 14565
rect 9371 14499 9437 14543
rect 9539 14543 9555 14577
rect 9589 14543 9605 14577
rect 9688 14545 9723 14579
rect 9757 14545 9823 14579
rect 9857 14545 9879 14579
rect 9913 14650 9971 14666
rect 9947 14616 9971 14650
rect 9913 14582 9971 14616
rect 9947 14548 9971 14582
rect 9539 14499 9605 14543
rect 9913 14499 9971 14548
rect 9344 14465 9373 14499
rect 9407 14465 9465 14499
rect 9499 14465 9557 14499
rect 9591 14465 9649 14499
rect 9683 14465 9741 14499
rect 9775 14465 9833 14499
rect 9867 14465 9925 14499
rect 9959 14465 9988 14499
rect 9442 14265 9471 14299
rect 9505 14265 9563 14299
rect 9597 14265 9655 14299
rect 9689 14265 9747 14299
rect 9781 14265 9839 14299
rect 9873 14265 9902 14299
rect 9499 14181 9555 14265
rect 9689 14223 9755 14265
rect 10690 14253 10719 14287
rect 10753 14253 10811 14287
rect 10845 14253 10903 14287
rect 10937 14253 10995 14287
rect 11029 14253 11087 14287
rect 11121 14253 11179 14287
rect 11213 14253 11271 14287
rect 11305 14253 11334 14287
rect 9499 14147 9513 14181
rect 9547 14147 9555 14181
rect 9499 14131 9555 14147
rect 9589 14181 9649 14197
rect 9589 14147 9597 14181
rect 9631 14147 9649 14181
rect 9589 14087 9649 14147
rect 9689 14189 9705 14223
rect 9739 14189 9755 14223
rect 9689 14155 9755 14189
rect 9689 14121 9705 14155
rect 9739 14121 9755 14155
rect 9793 14223 9885 14231
rect 9793 14189 9809 14223
rect 9843 14189 9885 14223
rect 9793 14155 9885 14189
rect 10708 14211 10775 14253
rect 10708 14177 10725 14211
rect 10759 14177 10775 14211
rect 10809 14203 10859 14219
rect 9793 14121 9809 14155
rect 9843 14121 9885 14155
rect 10809 14169 10817 14203
rect 10851 14169 10859 14203
rect 9462 14010 9515 14075
rect 9589 14053 9777 14087
rect 9462 13970 9464 14010
rect 9506 14003 9515 14010
rect 9743 14003 9777 14053
rect 9506 13987 9597 14003
rect 9506 13970 9516 13987
rect 9462 13953 9516 13970
rect 9550 13953 9597 13987
rect 9641 14000 9709 14003
rect 9641 13960 9654 14000
rect 9696 13960 9709 14000
rect 9641 13953 9657 13960
rect 9691 13953 9709 13960
rect 9743 13987 9801 14003
rect 9743 13953 9765 13987
rect 9799 13953 9801 13987
rect 9743 13937 9801 13953
rect 9743 13919 9777 13937
rect 9499 13881 9777 13919
rect 9835 13888 9885 14121
rect 9499 13859 9565 13881
rect 9499 13825 9513 13859
rect 9547 13825 9565 13859
rect 9835 13854 9844 13888
rect 9880 13854 9885 13888
rect 10707 13980 10755 14141
rect 10809 14059 10859 14169
rect 10903 14211 10969 14253
rect 10903 14177 10919 14211
rect 10953 14177 10969 14211
rect 10903 14109 10969 14177
rect 11006 14203 11056 14219
rect 11006 14169 11014 14203
rect 11048 14169 11056 14203
rect 11006 14059 11056 14169
rect 11149 14211 11215 14253
rect 12588 14237 12617 14271
rect 12651 14237 12709 14271
rect 12743 14237 12801 14271
rect 12835 14237 12893 14271
rect 12927 14237 12985 14271
rect 13019 14237 13077 14271
rect 13111 14237 13140 14271
rect 11149 14177 11165 14211
rect 11199 14177 11215 14211
rect 11149 14143 11215 14177
rect 11249 14211 11317 14219
rect 11249 14177 11265 14211
rect 11299 14177 11317 14211
rect 12971 14195 13027 14237
rect 11249 14167 11317 14177
rect 11149 14109 11165 14143
rect 11199 14109 11215 14143
rect 11149 14093 11215 14109
rect 11265 14143 11317 14167
rect 11299 14109 11317 14143
rect 12606 14183 12937 14193
rect 12606 14170 12845 14183
rect 12606 14136 12762 14170
rect 12798 14149 12845 14170
rect 12879 14149 12937 14183
rect 12798 14136 12937 14149
rect 12606 14135 12937 14136
rect 12971 14161 12984 14195
rect 13018 14161 13027 14195
rect 11265 14075 11317 14109
rect 12971 14127 13027 14161
rect 10707 13946 10716 13980
rect 10750 13975 10755 13980
rect 10707 13941 10721 13946
rect 10707 13879 10755 13941
rect 10789 14025 11227 14059
rect 9835 13847 9885 13854
rect 9499 13809 9565 13825
rect 9689 13831 9739 13847
rect 9689 13797 9705 13831
rect 9689 13755 9739 13797
rect 9773 13831 9885 13847
rect 10789 13843 10823 14025
rect 11164 13991 11227 14025
rect 11299 14041 11317 14075
rect 9773 13797 9789 13831
rect 9823 13797 9885 13831
rect 9773 13789 9885 13797
rect 10724 13827 10823 13843
rect 10724 13793 10725 13827
rect 10759 13793 10823 13827
rect 10867 13975 10937 13991
rect 10901 13941 10937 13975
rect 10867 13884 10937 13941
rect 10867 13850 10886 13884
rect 10920 13850 10937 13884
rect 10867 13798 10937 13850
rect 10973 13975 11033 13991
rect 11007 13941 11033 13975
rect 10973 13924 11033 13941
rect 10973 13890 10984 13924
rect 11018 13890 11033 13924
rect 10973 13797 11033 13890
rect 11069 13975 11125 13991
rect 11103 13974 11125 13975
rect 11069 13936 11078 13941
rect 11114 13936 11125 13974
rect 11164 13975 11230 13991
rect 11164 13941 11180 13975
rect 11214 13941 11230 13975
rect 11069 13797 11125 13936
rect 11161 13887 11215 13903
rect 11265 13887 11317 14041
rect 12606 14067 12924 14101
rect 12971 14093 12984 14127
rect 13018 14093 13027 14127
rect 12971 14077 13027 14093
rect 13069 14164 13123 14203
rect 13103 14130 13123 14164
rect 13069 14096 13123 14130
rect 13103 14080 13123 14096
rect 12606 14064 12670 14067
rect 12606 14030 12623 14064
rect 12657 14030 12670 14064
rect 12890 14043 12924 14067
rect 12606 14009 12670 14030
rect 12606 13959 12676 13975
rect 12606 13942 12623 13959
rect 12657 13942 12676 13959
rect 11161 13853 11166 13887
rect 11200 13853 11215 13887
rect 11161 13819 11215 13853
rect 10724 13777 10823 13793
rect 11161 13785 11166 13819
rect 11200 13785 11215 13819
rect 11249 13856 11265 13887
rect 11249 13818 11260 13856
rect 11299 13853 11317 13887
rect 11660 13879 11689 13913
rect 11723 13879 11781 13913
rect 11815 13879 11873 13913
rect 11907 13879 11965 13913
rect 11999 13879 12057 13913
rect 12091 13879 12120 13913
rect 12606 13908 12618 13942
rect 12658 13908 12676 13942
rect 12710 13964 12852 14033
rect 12890 14009 13035 14043
rect 13069 14040 13078 14062
rect 13120 14040 13123 14080
rect 13069 14009 13123 14040
rect 13001 13975 13035 14009
rect 12710 13922 12746 13964
rect 12796 13922 12852 13964
rect 12710 13909 12852 13922
rect 12886 13960 12967 13975
rect 12886 13924 12918 13960
rect 12956 13959 12967 13960
rect 12959 13925 12967 13959
rect 12956 13924 12967 13925
rect 12886 13909 12967 13924
rect 13001 13959 13055 13975
rect 13001 13925 13021 13959
rect 13001 13909 13055 13925
rect 11298 13819 11317 13853
rect 11249 13785 11265 13818
rect 11299 13785 11317 13819
rect 11889 13821 11955 13879
rect 12606 13861 12676 13908
rect 13001 13875 13035 13909
rect 11889 13787 11905 13821
rect 11939 13787 11955 13821
rect 9442 13721 9471 13755
rect 9505 13721 9563 13755
rect 9597 13721 9655 13755
rect 9689 13721 9747 13755
rect 9781 13721 9839 13755
rect 9873 13721 9902 13755
rect 11161 13743 11215 13785
rect 11889 13753 11955 13787
rect 10690 13709 10719 13743
rect 10753 13709 10811 13743
rect 10845 13709 10903 13743
rect 10937 13709 10995 13743
rect 11029 13709 11087 13743
rect 11121 13709 11179 13743
rect 11213 13709 11271 13743
rect 11305 13709 11334 13743
rect 11714 13701 11792 13720
rect 11889 13719 11905 13753
rect 11939 13719 11955 13753
rect 11989 13837 12096 13845
rect 11989 13803 12005 13837
rect 12039 13803 12096 13837
rect 12713 13841 13035 13875
rect 13089 13862 13123 14009
rect 13069 13845 13123 13862
rect 11989 13769 12096 13803
rect 11989 13735 12005 13769
rect 12039 13768 12096 13769
rect 11989 13734 12028 13735
rect 12062 13734 12096 13768
rect 11989 13721 12096 13734
rect 12607 13793 12623 13827
rect 12657 13793 12673 13827
rect 12607 13727 12673 13793
rect 12713 13821 12747 13841
rect 12887 13821 12921 13841
rect 12713 13771 12747 13787
rect 12787 13773 12803 13807
rect 12837 13773 12853 13807
rect 12787 13727 12853 13773
rect 13103 13811 13123 13845
rect 12887 13771 12921 13787
rect 12955 13773 12981 13807
rect 13015 13773 13031 13807
rect 13069 13793 13123 13811
rect 12955 13727 13031 13773
rect 11714 13667 11736 13701
rect 11770 13685 11792 13701
rect 11770 13667 11999 13685
rect 11714 13651 11999 13667
rect 11689 13601 11760 13617
rect 11689 13567 11726 13601
rect 11689 13558 11760 13567
rect 11689 13524 11700 13558
rect 11734 13524 11760 13558
rect 11689 13505 11760 13524
rect 11794 13471 11828 13651
rect 11862 13608 11915 13617
rect 11862 13601 11878 13608
rect 11912 13574 11915 13608
rect 11896 13567 11915 13574
rect 11862 13505 11915 13567
rect 11965 13601 11999 13651
rect 11965 13551 11999 13567
rect 12033 13517 12096 13721
rect 12588 13693 12617 13727
rect 12651 13693 12709 13727
rect 12743 13693 12801 13727
rect 12835 13693 12893 13727
rect 12927 13693 12985 13727
rect 13019 13693 13077 13727
rect 13111 13693 13140 13727
rect 11973 13515 12096 13517
rect 11973 13481 11989 13515
rect 12023 13481 12096 13515
rect 11710 13455 11758 13471
rect 10814 13411 10843 13445
rect 10877 13411 10935 13445
rect 10969 13411 11027 13445
rect 11061 13411 11119 13445
rect 11153 13411 11211 13445
rect 11245 13411 11274 13445
rect 11710 13421 11724 13455
rect 9336 13341 9365 13375
rect 9399 13341 9457 13375
rect 9491 13341 9549 13375
rect 9583 13341 9641 13375
rect 9675 13341 9733 13375
rect 9767 13341 9825 13375
rect 9859 13341 9917 13375
rect 9951 13341 9980 13375
rect 9353 13299 9429 13307
rect 9353 13265 9379 13299
rect 9413 13265 9429 13299
rect 9353 13231 9429 13265
rect 9353 13197 9379 13231
rect 9413 13197 9429 13231
rect 9353 13171 9429 13197
rect 9547 13289 9581 13341
rect 9547 13221 9581 13255
rect 9547 13171 9581 13187
rect 9615 13289 9681 13307
rect 9615 13255 9631 13289
rect 9665 13255 9681 13289
rect 9615 13221 9681 13255
rect 9715 13289 9749 13341
rect 9715 13239 9749 13255
rect 9783 13289 9863 13307
rect 9783 13255 9819 13289
rect 9853 13255 9863 13289
rect 9615 13187 9631 13221
rect 9665 13205 9681 13221
rect 9783 13221 9863 13255
rect 9783 13205 9819 13221
rect 9665 13187 9819 13205
rect 9853 13187 9863 13221
rect 9615 13171 9863 13187
rect 9899 13291 9963 13307
rect 9899 13257 9903 13291
rect 9937 13257 9963 13291
rect 10831 13300 10952 13411
rect 10987 13360 11083 13377
rect 11021 13338 11083 13360
rect 10987 13309 11012 13326
rect 11048 13309 11083 13338
rect 11117 13369 11168 13411
rect 11117 13335 11121 13369
rect 11155 13335 11168 13369
rect 11117 13302 11168 13335
rect 11202 13355 11257 13377
rect 11710 13369 11758 13421
rect 11794 13455 11850 13471
rect 11794 13421 11808 13455
rect 11842 13421 11850 13455
rect 11794 13405 11850 13421
rect 11896 13455 11939 13471
rect 11896 13421 11904 13455
rect 11938 13421 11939 13455
rect 11896 13369 11939 13421
rect 11973 13447 12096 13481
rect 11973 13413 11989 13447
rect 12023 13413 12096 13447
rect 11973 13403 12096 13413
rect 11202 13321 11205 13355
rect 11239 13321 11257 13355
rect 11660 13335 11689 13369
rect 11723 13335 11781 13369
rect 11815 13335 11873 13369
rect 11907 13335 11965 13369
rect 11999 13335 12057 13369
rect 12091 13335 12120 13369
rect 10831 13280 10954 13300
rect 9899 13224 9963 13257
rect 10917 13275 10954 13280
rect 11202 13287 11257 13321
rect 10917 13260 10983 13275
rect 9899 13223 9914 13224
rect 9899 13189 9903 13223
rect 9948 13190 9963 13224
rect 9937 13189 9963 13190
rect 9353 12979 9387 13171
rect 9899 13155 9963 13189
rect 9421 13103 9682 13137
rect 9899 13121 9903 13155
rect 9937 13121 9963 13155
rect 10831 13230 10883 13246
rect 10831 13196 10849 13230
rect 10917 13226 10933 13260
rect 10967 13226 10983 13260
rect 11017 13241 11168 13261
rect 11017 13211 11026 13241
rect 11014 13207 11026 13211
rect 11060 13207 11168 13241
rect 11202 13253 11205 13287
rect 11239 13282 11257 13287
rect 11202 13244 11208 13253
rect 11246 13244 11257 13282
rect 11202 13237 11257 13244
rect 11014 13204 11168 13207
rect 11011 13202 11168 13204
rect 11010 13199 11189 13202
rect 11006 13196 11189 13199
rect 10831 13156 10883 13196
rect 11002 13194 11189 13196
rect 10997 13192 11189 13194
rect 10983 13186 11189 13192
rect 10979 13180 11189 13186
rect 10975 13174 11189 13180
rect 10969 13169 11189 13174
rect 10962 13162 11189 13169
rect 10956 13161 11189 13162
rect 10956 13160 11034 13161
rect 10956 13158 11029 13160
rect 10956 13157 11026 13158
rect 10956 13156 11023 13157
rect 10831 13155 11023 13156
rect 10831 13153 11021 13155
rect 10831 13152 11019 13153
rect 10831 13150 11017 13152
rect 10831 13148 11016 13150
rect 10831 13147 11015 13148
rect 10831 13144 11013 13147
rect 10831 13141 11012 13144
rect 10831 13136 11010 13141
rect 10831 13122 11009 13136
rect 11143 13133 11189 13161
rect 9421 13064 9470 13103
rect 9421 13063 9422 13064
rect 9456 13030 9470 13064
rect 9455 13029 9470 13030
rect 9504 13066 9614 13069
rect 9504 13063 9542 13066
rect 9504 13029 9538 13063
rect 9576 13032 9614 13066
rect 9572 13029 9614 13032
rect 9648 13063 9682 13103
rect 9837 13087 9963 13121
rect 10831 13087 10941 13088
rect 9757 13063 9803 13079
rect 9648 13029 9673 13063
rect 9707 13029 9723 13063
rect 9757 13029 9769 13063
rect 9421 13013 9470 13029
rect 9757 12979 9803 13029
rect 9353 12945 9803 12979
rect 9463 12931 9497 12945
rect 9363 12875 9379 12909
rect 9413 12875 9429 12909
rect 9837 12911 9871 13087
rect 10831 13053 10849 13087
rect 10883 13064 10941 13087
rect 10831 13030 10860 13053
rect 10894 13030 10941 13064
rect 10831 13011 10941 13030
rect 9463 12881 9497 12897
rect 9363 12831 9429 12875
rect 9531 12875 9547 12909
rect 9581 12875 9597 12909
rect 9680 12877 9715 12911
rect 9749 12877 9815 12911
rect 9849 12877 9871 12911
rect 9905 12982 9963 12998
rect 9939 12948 9963 12982
rect 10975 12977 11009 13122
rect 9905 12914 9963 12948
rect 10831 12943 10849 12977
rect 10883 12943 11009 12977
rect 11043 13093 11059 13127
rect 11093 13093 11109 13127
rect 11043 13070 11109 13093
rect 11143 13099 11155 13133
rect 11143 13082 11189 13099
rect 11043 13036 11062 13070
rect 11098 13042 11109 13070
rect 11043 12945 11087 13036
rect 11223 13031 11257 13237
rect 11121 12993 11171 13009
rect 11155 12959 11171 12993
rect 9939 12880 9963 12914
rect 11121 12901 11171 12959
rect 11205 13003 11257 13031
rect 11239 12969 11257 13003
rect 11205 12935 11257 12969
rect 9531 12831 9597 12875
rect 9905 12831 9963 12880
rect 10814 12867 10843 12901
rect 10877 12867 10935 12901
rect 10969 12867 11027 12901
rect 11061 12867 11119 12901
rect 11153 12867 11211 12901
rect 11245 12867 11274 12901
rect 9336 12797 9365 12831
rect 9399 12797 9457 12831
rect 9491 12797 9549 12831
rect 9583 12797 9641 12831
rect 9675 12797 9733 12831
rect 9767 12797 9825 12831
rect 9859 12797 9917 12831
rect 9951 12797 9980 12831
rect 9434 12597 9463 12631
rect 9497 12597 9555 12631
rect 9589 12597 9647 12631
rect 9681 12597 9739 12631
rect 9773 12597 9831 12631
rect 9865 12597 9894 12631
rect 9491 12513 9547 12597
rect 9681 12555 9747 12597
rect 9491 12479 9505 12513
rect 9539 12479 9547 12513
rect 9491 12463 9547 12479
rect 9581 12513 9641 12529
rect 9581 12479 9589 12513
rect 9623 12479 9641 12513
rect 9581 12419 9641 12479
rect 9681 12521 9697 12555
rect 9731 12521 9747 12555
rect 9681 12487 9747 12521
rect 9681 12453 9697 12487
rect 9731 12453 9747 12487
rect 9785 12555 9877 12563
rect 9785 12521 9801 12555
rect 9835 12521 9877 12555
rect 9785 12487 9877 12521
rect 9785 12453 9801 12487
rect 9835 12453 9877 12487
rect 9454 12342 9507 12407
rect 9581 12385 9769 12419
rect 9454 12302 9456 12342
rect 9498 12335 9507 12342
rect 9735 12335 9769 12385
rect 9827 12374 9877 12453
rect 10810 12391 10839 12425
rect 10873 12391 10931 12425
rect 10965 12391 11023 12425
rect 11057 12391 11115 12425
rect 11149 12391 11207 12425
rect 11241 12391 11270 12425
rect 9827 12340 9836 12374
rect 9872 12340 9877 12374
rect 9498 12319 9589 12335
rect 9498 12302 9508 12319
rect 9454 12285 9508 12302
rect 9542 12285 9589 12319
rect 9633 12332 9701 12335
rect 9633 12292 9646 12332
rect 9688 12292 9701 12332
rect 9633 12285 9649 12292
rect 9683 12285 9701 12292
rect 9735 12319 9793 12335
rect 9735 12285 9757 12319
rect 9791 12285 9793 12319
rect 9735 12269 9793 12285
rect 9735 12251 9769 12269
rect 9491 12213 9769 12251
rect 9491 12191 9557 12213
rect 9491 12157 9505 12191
rect 9539 12157 9557 12191
rect 9827 12179 9877 12340
rect 10867 12307 10923 12391
rect 11057 12349 11123 12391
rect 10867 12273 10881 12307
rect 10915 12273 10923 12307
rect 10867 12257 10923 12273
rect 10957 12307 11017 12323
rect 10957 12273 10965 12307
rect 10999 12273 11017 12307
rect 10957 12213 11017 12273
rect 11057 12315 11073 12349
rect 11107 12315 11123 12349
rect 11057 12281 11123 12315
rect 11057 12247 11073 12281
rect 11107 12247 11123 12281
rect 11161 12349 11253 12357
rect 11161 12315 11177 12349
rect 11211 12315 11253 12349
rect 11161 12281 11253 12315
rect 11161 12247 11177 12281
rect 11211 12247 11253 12281
rect 9491 12141 9557 12157
rect 9681 12163 9731 12179
rect 9681 12129 9697 12163
rect 9681 12087 9731 12129
rect 9765 12163 9877 12179
rect 9765 12129 9781 12163
rect 9815 12129 9877 12163
rect 9765 12121 9877 12129
rect 10830 12129 10883 12201
rect 10957 12179 11145 12213
rect 11111 12129 11145 12179
rect 11203 12200 11253 12247
rect 11203 12166 11212 12200
rect 11246 12166 11253 12200
rect 10830 12116 10965 12129
rect 9434 12053 9463 12087
rect 9497 12053 9555 12087
rect 9589 12053 9647 12087
rect 9681 12053 9739 12087
rect 9773 12053 9831 12087
rect 9865 12053 9894 12087
rect 10830 12079 10884 12116
rect 10920 12082 10965 12116
rect 10918 12079 10965 12082
rect 11009 12114 11077 12129
rect 11009 12080 11024 12114
rect 11060 12080 11077 12114
rect 11009 12079 11025 12080
rect 11059 12079 11077 12080
rect 11111 12113 11169 12129
rect 11111 12079 11133 12113
rect 11167 12079 11169 12113
rect 11111 12063 11169 12079
rect 11111 12045 11145 12063
rect 10867 12007 11145 12045
rect 10867 11985 10933 12007
rect 10867 11951 10881 11985
rect 10915 11951 10933 11985
rect 11203 11973 11253 12166
rect 10867 11935 10933 11951
rect 11057 11957 11107 11973
rect 11057 11923 11073 11957
rect 11057 11881 11107 11923
rect 11141 11957 11253 11973
rect 11141 11923 11157 11957
rect 11191 11923 11253 11957
rect 11141 11915 11253 11923
rect 10810 11847 10839 11881
rect 10873 11847 10931 11881
rect 10965 11847 11023 11881
rect 11057 11847 11115 11881
rect 11149 11847 11207 11881
rect 11241 11847 11270 11881
rect 9346 11777 9375 11811
rect 9409 11777 9467 11811
rect 9501 11777 9559 11811
rect 9593 11777 9651 11811
rect 9685 11777 9743 11811
rect 9777 11777 9835 11811
rect 9869 11777 9927 11811
rect 9961 11777 9990 11811
rect 9363 11735 9439 11743
rect 9363 11701 9389 11735
rect 9423 11701 9439 11735
rect 9363 11667 9439 11701
rect 9363 11633 9389 11667
rect 9423 11633 9439 11667
rect 9363 11607 9439 11633
rect 9557 11725 9591 11777
rect 9557 11657 9591 11691
rect 9557 11607 9591 11623
rect 9625 11725 9691 11743
rect 9625 11691 9641 11725
rect 9675 11691 9691 11725
rect 9625 11657 9691 11691
rect 9725 11725 9759 11777
rect 9725 11675 9759 11691
rect 9793 11725 9873 11743
rect 9793 11691 9829 11725
rect 9863 11691 9873 11725
rect 9625 11623 9641 11657
rect 9675 11641 9691 11657
rect 9793 11657 9873 11691
rect 9793 11641 9829 11657
rect 9675 11623 9829 11641
rect 9863 11623 9873 11657
rect 9625 11607 9873 11623
rect 9909 11727 9973 11743
rect 9909 11693 9913 11727
rect 9947 11693 9973 11727
rect 9909 11660 9973 11693
rect 9909 11659 9914 11660
rect 9909 11625 9913 11659
rect 9950 11626 9973 11660
rect 9947 11625 9973 11626
rect 9363 11415 9397 11607
rect 9909 11591 9973 11625
rect 9431 11539 9692 11573
rect 9909 11557 9913 11591
rect 9947 11557 9973 11591
rect 9431 11500 9480 11539
rect 9431 11499 9432 11500
rect 9466 11466 9480 11500
rect 9465 11465 9480 11466
rect 9514 11502 9624 11505
rect 9514 11499 9552 11502
rect 9514 11465 9548 11499
rect 9586 11468 9624 11502
rect 9582 11465 9624 11468
rect 9658 11499 9692 11539
rect 9847 11523 9973 11557
rect 9767 11499 9813 11515
rect 9658 11465 9683 11499
rect 9717 11465 9733 11499
rect 9767 11465 9779 11499
rect 9431 11449 9480 11465
rect 9767 11415 9813 11465
rect 9363 11381 9813 11415
rect 9473 11367 9507 11381
rect 9373 11311 9389 11345
rect 9423 11311 9439 11345
rect 9847 11347 9881 11523
rect 9473 11317 9507 11333
rect 9373 11267 9439 11311
rect 9541 11311 9557 11345
rect 9591 11311 9607 11345
rect 9690 11313 9725 11347
rect 9759 11313 9825 11347
rect 9859 11313 9881 11347
rect 9915 11418 9973 11434
rect 9949 11384 9973 11418
rect 9915 11350 9973 11384
rect 9949 11316 9973 11350
rect 9541 11267 9607 11311
rect 9915 11267 9973 11316
rect 9346 11233 9375 11267
rect 9409 11233 9467 11267
rect 9501 11233 9559 11267
rect 9593 11233 9651 11267
rect 9685 11233 9743 11267
rect 9777 11233 9835 11267
rect 9869 11233 9927 11267
rect 9961 11233 9990 11267
rect 9444 11033 9473 11067
rect 9507 11033 9565 11067
rect 9599 11033 9657 11067
rect 9691 11033 9749 11067
rect 9783 11033 9841 11067
rect 9875 11033 9904 11067
rect 9501 10949 9557 11033
rect 9691 10991 9757 11033
rect 9501 10915 9515 10949
rect 9549 10915 9557 10949
rect 9501 10899 9557 10915
rect 9591 10949 9651 10965
rect 9591 10915 9599 10949
rect 9633 10915 9651 10949
rect 9591 10855 9651 10915
rect 9691 10957 9707 10991
rect 9741 10957 9757 10991
rect 9691 10923 9757 10957
rect 9691 10889 9707 10923
rect 9741 10889 9757 10923
rect 9795 10991 9887 10999
rect 9795 10957 9811 10991
rect 9845 10957 9887 10991
rect 9795 10923 9887 10957
rect 9795 10889 9811 10923
rect 9845 10889 9887 10923
rect 9464 10778 9517 10843
rect 9591 10821 9779 10855
rect 9464 10738 9466 10778
rect 9508 10771 9517 10778
rect 9745 10771 9779 10821
rect 9508 10755 9599 10771
rect 9508 10738 9518 10755
rect 9464 10721 9518 10738
rect 9552 10721 9599 10755
rect 9643 10768 9711 10771
rect 9643 10728 9656 10768
rect 9698 10728 9711 10768
rect 9643 10721 9659 10728
rect 9693 10721 9711 10728
rect 9745 10755 9803 10771
rect 9745 10721 9767 10755
rect 9801 10721 9803 10755
rect 9745 10705 9803 10721
rect 9837 10734 9887 10889
rect 9745 10687 9779 10705
rect 9501 10649 9779 10687
rect 9837 10698 9848 10734
rect 9882 10698 9887 10734
rect 9501 10627 9567 10649
rect 9501 10593 9515 10627
rect 9549 10593 9567 10627
rect 9837 10615 9887 10698
rect 9501 10577 9567 10593
rect 9691 10599 9741 10615
rect 9691 10565 9707 10599
rect 9691 10523 9741 10565
rect 9775 10599 9887 10615
rect 9775 10565 9791 10599
rect 9825 10565 9887 10599
rect 9775 10557 9887 10565
rect 9444 10489 9473 10523
rect 9507 10489 9565 10523
rect 9599 10489 9657 10523
rect 9691 10489 9749 10523
rect 9783 10489 9841 10523
rect 9875 10489 9904 10523
rect 6112 6583 6141 6617
rect 6175 6583 6233 6617
rect 6267 6583 6325 6617
rect 6359 6583 6388 6617
rect 6178 6537 6244 6549
rect 6178 6503 6194 6537
rect 6228 6503 6244 6537
rect 6178 6469 6244 6503
rect 6178 6435 6194 6469
rect 6228 6435 6244 6469
rect 6178 6423 6244 6435
rect 6278 6537 6324 6583
rect 6312 6503 6324 6537
rect 6278 6469 6324 6503
rect 6312 6435 6324 6469
rect 6178 6382 6224 6423
rect 6278 6419 6324 6435
rect 6212 6348 6224 6382
rect 6178 6303 6224 6348
rect 6258 6350 6274 6385
rect 6308 6350 6324 6385
rect 6258 6337 6324 6350
rect 6178 6285 6244 6303
rect 6178 6251 6194 6285
rect 6228 6251 6244 6285
rect 6178 6217 6244 6251
rect 6178 6183 6194 6217
rect 6228 6183 6244 6217
rect 6178 6149 6244 6183
rect 6178 6115 6194 6149
rect 6228 6115 6244 6149
rect 6178 6107 6244 6115
rect 6278 6285 6320 6301
rect 6312 6251 6320 6285
rect 6278 6217 6320 6251
rect 6312 6183 6320 6217
rect 6278 6149 6320 6183
rect 6312 6115 6320 6149
rect 6278 6073 6320 6115
rect 6112 6039 6141 6073
rect 6175 6039 6233 6073
rect 6267 6039 6325 6073
rect 6359 6039 6388 6073
rect 10018 5951 10047 5985
rect 10081 5951 10139 5985
rect 10173 5951 10231 5985
rect 10265 5951 10323 5985
rect 10357 5951 10415 5985
rect 10449 5951 10507 5985
rect 10541 5951 10599 5985
rect 10633 5951 10691 5985
rect 10725 5951 10783 5985
rect 10817 5951 10875 5985
rect 10909 5951 10967 5985
rect 11001 5951 11059 5985
rect 11093 5951 11151 5985
rect 11185 5951 11243 5985
rect 11277 5951 11335 5985
rect 11369 5951 11427 5985
rect 11461 5951 11490 5985
rect 10042 5873 10122 5917
rect 10171 5913 10237 5951
rect 10171 5879 10187 5913
rect 10221 5879 10237 5913
rect 10271 5901 10473 5917
rect 10042 5839 10088 5873
rect 10271 5867 10439 5901
rect 10271 5845 10305 5867
rect 10439 5849 10473 5867
rect 10540 5896 10574 5917
rect 10608 5913 10674 5951
rect 10608 5879 10624 5913
rect 10658 5879 10674 5913
rect 10708 5896 10742 5917
rect 10042 5806 10122 5839
rect 10157 5811 10305 5845
rect 10540 5845 10574 5862
rect 10776 5904 10842 5951
rect 10776 5870 10792 5904
rect 10826 5870 10842 5904
rect 10896 5896 10930 5917
rect 10708 5845 10742 5862
rect 10042 5671 10108 5806
rect 10157 5769 10191 5811
rect 10142 5753 10191 5769
rect 10398 5781 10410 5815
rect 10444 5781 10497 5815
rect 10540 5811 10742 5845
rect 10964 5913 11030 5951
rect 10964 5879 10980 5913
rect 11014 5879 11030 5913
rect 11064 5896 11098 5917
rect 10896 5845 10930 5862
rect 11064 5845 11098 5862
rect 10896 5811 11098 5845
rect 11148 5896 11268 5917
rect 11182 5862 11268 5896
rect 11321 5909 11387 5951
rect 12080 5939 12109 5973
rect 12143 5939 12201 5973
rect 12235 5939 12293 5973
rect 12327 5939 12385 5973
rect 12419 5939 12477 5973
rect 12511 5939 12569 5973
rect 12603 5939 12661 5973
rect 12695 5939 12753 5973
rect 12787 5939 12845 5973
rect 12879 5939 12937 5973
rect 12971 5939 13029 5973
rect 13063 5939 13121 5973
rect 13155 5939 13213 5973
rect 13247 5939 13305 5973
rect 13339 5939 13397 5973
rect 13431 5939 13489 5973
rect 13523 5939 13552 5973
rect 14038 5947 14067 5981
rect 14101 5947 14159 5981
rect 14193 5947 14251 5981
rect 14285 5947 14343 5981
rect 14377 5947 14435 5981
rect 14469 5947 14527 5981
rect 14561 5947 14619 5981
rect 14653 5947 14711 5981
rect 14745 5947 14803 5981
rect 14837 5947 14895 5981
rect 14929 5947 14987 5981
rect 15021 5947 15079 5981
rect 15113 5947 15171 5981
rect 15205 5947 15263 5981
rect 15297 5947 15355 5981
rect 15389 5947 15447 5981
rect 15481 5947 15510 5981
rect 16032 5953 16061 5987
rect 16095 5953 16153 5987
rect 16187 5953 16245 5987
rect 16279 5953 16337 5987
rect 16371 5953 16429 5987
rect 16463 5953 16521 5987
rect 16555 5953 16613 5987
rect 16647 5953 16705 5987
rect 16739 5953 16797 5987
rect 16831 5953 16889 5987
rect 16923 5953 16981 5987
rect 17015 5953 17073 5987
rect 17107 5953 17165 5987
rect 17199 5953 17257 5987
rect 17291 5953 17349 5987
rect 17383 5953 17441 5987
rect 17475 5953 17504 5987
rect 11321 5875 11337 5909
rect 11371 5875 11387 5909
rect 11148 5841 11268 5862
rect 11421 5873 11473 5917
rect 11148 5815 11387 5841
rect 11148 5781 11150 5815
rect 11184 5807 11387 5815
rect 11184 5781 11196 5807
rect 10398 5777 10497 5781
rect 10176 5719 10191 5753
rect 10142 5703 10191 5719
rect 10225 5747 10241 5761
rect 10225 5713 10226 5747
rect 10275 5727 10313 5761
rect 10398 5743 10481 5777
rect 10515 5743 10531 5777
rect 10565 5743 10581 5777
rect 10615 5747 10640 5777
rect 10260 5713 10313 5727
rect 10565 5713 10594 5743
rect 10628 5713 10640 5747
rect 10699 5718 10932 5775
rect 11353 5769 11387 5807
rect 11455 5839 11473 5873
rect 11421 5802 11473 5839
rect 10042 5633 10122 5671
rect 10042 5599 10088 5633
rect 1836 5531 1865 5565
rect 1899 5531 1957 5565
rect 1991 5531 2049 5565
rect 2083 5531 2141 5565
rect 2175 5531 2233 5565
rect 2267 5531 2325 5565
rect 2359 5531 2417 5565
rect 2451 5531 2509 5565
rect 2543 5531 2601 5565
rect 2635 5531 2693 5565
rect 2727 5531 2785 5565
rect 2819 5531 2877 5565
rect 2911 5531 2969 5565
rect 3003 5531 3061 5565
rect 3095 5531 3153 5565
rect 3187 5531 3245 5565
rect 3279 5531 3308 5565
rect 1860 5453 1940 5497
rect 1989 5493 2055 5531
rect 1989 5459 2005 5493
rect 2039 5459 2055 5493
rect 2089 5481 2291 5497
rect 1860 5419 1906 5453
rect 2089 5447 2257 5481
rect 2089 5425 2123 5447
rect 2257 5429 2291 5447
rect 2358 5476 2392 5497
rect 2426 5493 2492 5531
rect 2426 5459 2442 5493
rect 2476 5459 2492 5493
rect 2526 5476 2560 5497
rect 1860 5386 1940 5419
rect 1975 5391 2123 5425
rect 2358 5425 2392 5442
rect 2594 5484 2660 5531
rect 2594 5450 2610 5484
rect 2644 5450 2660 5484
rect 2714 5476 2748 5497
rect 2526 5425 2560 5442
rect 1860 5251 1926 5386
rect 1975 5349 2009 5391
rect 1960 5333 2009 5349
rect 2216 5361 2228 5395
rect 2262 5361 2315 5395
rect 2358 5391 2560 5425
rect 2782 5493 2848 5531
rect 2782 5459 2798 5493
rect 2832 5459 2848 5493
rect 2882 5476 2916 5497
rect 2714 5425 2748 5442
rect 2882 5425 2916 5442
rect 2714 5391 2916 5425
rect 2966 5476 3086 5497
rect 3000 5442 3086 5476
rect 3139 5489 3205 5531
rect 3970 5523 3999 5557
rect 4033 5523 4091 5557
rect 4125 5523 4183 5557
rect 4217 5523 4275 5557
rect 4309 5523 4367 5557
rect 4401 5523 4459 5557
rect 4493 5523 4551 5557
rect 4585 5523 4643 5557
rect 4677 5523 4735 5557
rect 4769 5523 4827 5557
rect 4861 5523 4919 5557
rect 4953 5523 5011 5557
rect 5045 5523 5103 5557
rect 5137 5523 5195 5557
rect 5229 5523 5287 5557
rect 5321 5523 5379 5557
rect 5413 5523 5442 5557
rect 5922 5523 5951 5557
rect 5985 5523 6043 5557
rect 6077 5523 6135 5557
rect 6169 5523 6227 5557
rect 6261 5523 6319 5557
rect 6353 5523 6411 5557
rect 6445 5523 6503 5557
rect 6537 5523 6595 5557
rect 6629 5523 6687 5557
rect 6721 5523 6779 5557
rect 6813 5523 6871 5557
rect 6905 5523 6963 5557
rect 6997 5523 7055 5557
rect 7089 5523 7147 5557
rect 7181 5523 7239 5557
rect 7273 5523 7331 5557
rect 7365 5523 7394 5557
rect 7924 5529 7953 5563
rect 7987 5529 8045 5563
rect 8079 5529 8137 5563
rect 8171 5529 8229 5563
rect 8263 5529 8321 5563
rect 8355 5529 8413 5563
rect 8447 5529 8505 5563
rect 8539 5529 8597 5563
rect 8631 5529 8689 5563
rect 8723 5529 8781 5563
rect 8815 5529 8873 5563
rect 8907 5529 8965 5563
rect 8999 5529 9057 5563
rect 9091 5529 9149 5563
rect 9183 5529 9241 5563
rect 9275 5529 9333 5563
rect 9367 5529 9396 5563
rect 10042 5543 10122 5599
rect 10157 5581 10191 5703
rect 10279 5649 10318 5679
rect 10279 5615 10313 5649
rect 10352 5645 10363 5679
rect 10699 5665 10733 5718
rect 10347 5615 10363 5645
rect 10409 5649 10666 5665
rect 10443 5631 10666 5649
rect 10700 5631 10733 5665
rect 10778 5679 10850 5681
rect 10812 5665 10850 5679
rect 10778 5631 10783 5645
rect 10817 5631 10850 5665
rect 10443 5615 10459 5631
rect 10778 5615 10850 5631
rect 10898 5649 10932 5718
rect 10966 5747 11044 5762
rect 11242 5753 11308 5769
rect 11242 5747 11274 5753
rect 11000 5746 11044 5747
rect 11000 5713 11010 5746
rect 10966 5712 11010 5713
rect 10966 5696 11044 5712
rect 11082 5713 11106 5747
rect 11140 5713 11156 5747
rect 11276 5713 11308 5719
rect 11082 5649 11116 5713
rect 11274 5703 11308 5713
rect 11353 5753 11404 5769
rect 11353 5719 11370 5753
rect 11353 5703 11404 5719
rect 10898 5615 11116 5649
rect 11184 5645 11230 5679
rect 11150 5642 11230 5645
rect 11353 5643 11387 5703
rect 11438 5671 11473 5802
rect 10409 5614 10459 5615
rect 10157 5547 10290 5581
rect 10409 5580 10418 5614
rect 10452 5580 10459 5614
rect 11150 5608 11196 5642
rect 11150 5592 11230 5608
rect 10409 5577 10459 5580
rect 3139 5455 3155 5489
rect 3189 5455 3205 5489
rect 2966 5421 3086 5442
rect 3239 5453 3291 5497
rect 2966 5395 3205 5421
rect 2966 5361 2968 5395
rect 3002 5387 3205 5395
rect 3002 5361 3014 5387
rect 2216 5357 2315 5361
rect 1994 5299 2009 5333
rect 1960 5283 2009 5299
rect 2043 5327 2059 5341
rect 2043 5293 2044 5327
rect 2093 5307 2131 5341
rect 2216 5323 2299 5357
rect 2333 5323 2349 5357
rect 2383 5323 2399 5357
rect 2433 5327 2458 5357
rect 2078 5293 2131 5307
rect 2383 5293 2412 5323
rect 2446 5293 2458 5327
rect 2517 5298 2750 5355
rect 3171 5349 3205 5387
rect 3273 5419 3291 5453
rect 3239 5382 3291 5419
rect 1860 5213 1940 5251
rect 1860 5179 1906 5213
rect 1860 5123 1940 5179
rect 1975 5161 2009 5283
rect 2097 5229 2136 5259
rect 2097 5195 2131 5229
rect 2170 5225 2181 5259
rect 2517 5245 2551 5298
rect 2165 5195 2181 5225
rect 2227 5229 2484 5245
rect 2261 5211 2484 5229
rect 2518 5211 2551 5245
rect 2596 5259 2668 5261
rect 2630 5245 2668 5259
rect 2596 5211 2601 5225
rect 2635 5211 2668 5245
rect 2261 5195 2277 5211
rect 2596 5195 2668 5211
rect 2716 5229 2750 5298
rect 2784 5327 2862 5342
rect 3060 5333 3126 5349
rect 3060 5327 3092 5333
rect 2818 5326 2862 5327
rect 2818 5293 2828 5326
rect 2784 5292 2828 5293
rect 2784 5276 2862 5292
rect 2900 5293 2924 5327
rect 2958 5293 2974 5327
rect 3094 5293 3126 5299
rect 2900 5229 2934 5293
rect 3092 5283 3126 5293
rect 3171 5333 3222 5349
rect 3171 5299 3188 5333
rect 3171 5283 3222 5299
rect 2716 5195 2934 5229
rect 3002 5225 3048 5259
rect 2968 5222 3048 5225
rect 3171 5223 3205 5283
rect 3256 5251 3291 5382
rect 2227 5194 2277 5195
rect 1975 5127 2108 5161
rect 2227 5160 2236 5194
rect 2270 5160 2277 5194
rect 2968 5188 3014 5222
rect 2968 5172 3048 5188
rect 2227 5157 2277 5160
rect 1860 5089 1906 5123
rect 2074 5123 2108 5127
rect 2358 5127 2560 5161
rect 2074 5105 2291 5123
rect 1860 5055 1940 5089
rect 1974 5059 1990 5093
rect 2024 5059 2040 5093
rect 1974 5021 2040 5059
rect 2074 5071 2257 5105
rect 2074 5055 2291 5071
rect 2358 5110 2392 5127
rect 2526 5110 2560 5127
rect 2358 5055 2392 5076
rect 2426 5059 2442 5093
rect 2476 5059 2492 5093
rect 2426 5021 2492 5059
rect 2701 5127 2916 5161
rect 3087 5159 3205 5223
rect 3239 5210 3291 5251
rect 3273 5186 3291 5210
rect 3087 5135 3121 5159
rect 2701 5110 2748 5127
rect 2526 5055 2560 5076
rect 2594 5063 2610 5097
rect 2644 5063 2660 5097
rect 2594 5021 2660 5063
rect 2701 5076 2714 5110
rect 2882 5110 2916 5127
rect 2701 5055 2748 5076
rect 2782 5059 2798 5093
rect 2832 5059 2848 5093
rect 2782 5021 2848 5059
rect 2882 5055 2916 5076
rect 2966 5110 3121 5135
rect 3239 5150 3244 5176
rect 3284 5150 3291 5186
rect 3000 5076 3121 5110
rect 2966 5055 3121 5076
rect 3155 5101 3205 5118
rect 3189 5067 3205 5101
rect 3155 5021 3205 5067
rect 3239 5116 3291 5150
rect 3273 5082 3291 5116
rect 3239 5055 3291 5082
rect 3994 5445 4074 5489
rect 4123 5485 4189 5523
rect 4123 5451 4139 5485
rect 4173 5451 4189 5485
rect 4223 5473 4425 5489
rect 3994 5411 4040 5445
rect 4223 5439 4391 5473
rect 4223 5417 4257 5439
rect 4391 5421 4425 5439
rect 4492 5468 4526 5489
rect 4560 5485 4626 5523
rect 4560 5451 4576 5485
rect 4610 5451 4626 5485
rect 4660 5468 4694 5489
rect 3994 5378 4074 5411
rect 4109 5383 4257 5417
rect 4492 5417 4526 5434
rect 4728 5476 4794 5523
rect 4728 5442 4744 5476
rect 4778 5442 4794 5476
rect 4848 5468 4882 5489
rect 4660 5417 4694 5434
rect 3994 5243 4060 5378
rect 4109 5341 4143 5383
rect 4094 5325 4143 5341
rect 4350 5353 4362 5387
rect 4396 5353 4449 5387
rect 4492 5383 4694 5417
rect 4916 5485 4982 5523
rect 4916 5451 4932 5485
rect 4966 5451 4982 5485
rect 5016 5468 5050 5489
rect 4848 5417 4882 5434
rect 5016 5417 5050 5434
rect 4848 5383 5050 5417
rect 5100 5468 5220 5489
rect 5134 5434 5220 5468
rect 5273 5481 5339 5523
rect 5273 5447 5289 5481
rect 5323 5447 5339 5481
rect 5100 5413 5220 5434
rect 5373 5445 5425 5489
rect 5100 5387 5339 5413
rect 5100 5353 5102 5387
rect 5136 5379 5339 5387
rect 5136 5353 5148 5379
rect 4350 5349 4449 5353
rect 4128 5291 4143 5325
rect 4094 5275 4143 5291
rect 4177 5319 4193 5333
rect 4177 5285 4178 5319
rect 4227 5299 4265 5333
rect 4350 5315 4433 5349
rect 4467 5315 4483 5349
rect 4517 5315 4533 5349
rect 4567 5319 4592 5349
rect 4212 5285 4265 5299
rect 4517 5285 4546 5315
rect 4580 5285 4592 5319
rect 4651 5290 4884 5347
rect 5305 5341 5339 5379
rect 5407 5411 5425 5445
rect 5373 5374 5425 5411
rect 3994 5205 4074 5243
rect 3994 5171 4040 5205
rect 3994 5115 4074 5171
rect 4109 5153 4143 5275
rect 4231 5221 4270 5251
rect 4231 5187 4265 5221
rect 4304 5217 4315 5251
rect 4651 5237 4685 5290
rect 4299 5187 4315 5217
rect 4361 5221 4618 5237
rect 4395 5203 4618 5221
rect 4652 5203 4685 5237
rect 4730 5251 4802 5253
rect 4764 5237 4802 5251
rect 4730 5203 4735 5217
rect 4769 5203 4802 5237
rect 4395 5187 4411 5203
rect 4730 5187 4802 5203
rect 4850 5221 4884 5290
rect 4918 5319 4996 5334
rect 5194 5325 5260 5341
rect 5194 5319 5226 5325
rect 4952 5318 4996 5319
rect 4952 5285 4962 5318
rect 4918 5284 4962 5285
rect 4918 5268 4996 5284
rect 5034 5285 5058 5319
rect 5092 5285 5108 5319
rect 5228 5285 5260 5291
rect 5034 5221 5068 5285
rect 5226 5275 5260 5285
rect 5305 5325 5356 5341
rect 5305 5291 5322 5325
rect 5305 5275 5356 5291
rect 4850 5187 5068 5221
rect 5136 5217 5182 5251
rect 5102 5214 5182 5217
rect 5305 5215 5339 5275
rect 5390 5243 5425 5374
rect 4361 5184 4411 5187
rect 4109 5119 4242 5153
rect 4361 5150 4368 5184
rect 4402 5150 4411 5184
rect 5102 5180 5148 5214
rect 5102 5164 5182 5180
rect 4361 5149 4411 5150
rect 3994 5081 4040 5115
rect 4208 5115 4242 5119
rect 4492 5119 4694 5153
rect 4208 5097 4425 5115
rect 3994 5047 4074 5081
rect 4108 5051 4124 5085
rect 4158 5051 4174 5085
rect 1836 4987 1865 5021
rect 1899 4987 1957 5021
rect 1991 4987 2049 5021
rect 2083 4987 2141 5021
rect 2175 4987 2233 5021
rect 2267 4987 2325 5021
rect 2359 4987 2417 5021
rect 2451 4987 2509 5021
rect 2543 4987 2601 5021
rect 2635 4987 2693 5021
rect 2727 4987 2785 5021
rect 2819 4987 2877 5021
rect 2911 4987 2969 5021
rect 3003 4987 3061 5021
rect 3095 4987 3153 5021
rect 3187 4987 3245 5021
rect 3279 4987 3308 5021
rect 4108 5013 4174 5051
rect 4208 5063 4391 5097
rect 4208 5047 4425 5063
rect 4492 5102 4526 5119
rect 4660 5102 4694 5119
rect 4492 5047 4526 5068
rect 4560 5051 4576 5085
rect 4610 5051 4626 5085
rect 4560 5013 4626 5051
rect 4835 5119 5050 5153
rect 5221 5151 5339 5215
rect 5373 5202 5425 5243
rect 5407 5178 5425 5202
rect 5221 5127 5255 5151
rect 4835 5102 4882 5119
rect 4660 5047 4694 5068
rect 4728 5055 4744 5089
rect 4778 5055 4794 5089
rect 4728 5013 4794 5055
rect 4835 5068 4848 5102
rect 5016 5102 5050 5119
rect 4835 5047 4882 5068
rect 4916 5051 4932 5085
rect 4966 5051 4982 5085
rect 4916 5013 4982 5051
rect 5016 5047 5050 5068
rect 5100 5102 5255 5127
rect 5373 5142 5384 5168
rect 5418 5142 5425 5178
rect 5134 5068 5255 5102
rect 5100 5047 5255 5068
rect 5289 5093 5339 5110
rect 5323 5059 5339 5093
rect 5289 5013 5339 5059
rect 5373 5108 5425 5142
rect 5407 5074 5425 5108
rect 5373 5047 5425 5074
rect 5946 5445 6026 5489
rect 6075 5485 6141 5523
rect 6075 5451 6091 5485
rect 6125 5451 6141 5485
rect 6175 5473 6377 5489
rect 5946 5411 5992 5445
rect 6175 5439 6343 5473
rect 6175 5417 6209 5439
rect 6343 5421 6377 5439
rect 6444 5468 6478 5489
rect 6512 5485 6578 5523
rect 6512 5451 6528 5485
rect 6562 5451 6578 5485
rect 6612 5468 6646 5489
rect 5946 5378 6026 5411
rect 6061 5383 6209 5417
rect 6444 5417 6478 5434
rect 6680 5476 6746 5523
rect 6680 5442 6696 5476
rect 6730 5442 6746 5476
rect 6800 5468 6834 5489
rect 6612 5417 6646 5434
rect 5946 5243 6012 5378
rect 6061 5341 6095 5383
rect 6046 5325 6095 5341
rect 6302 5353 6314 5387
rect 6348 5353 6401 5387
rect 6444 5383 6646 5417
rect 6868 5485 6934 5523
rect 6868 5451 6884 5485
rect 6918 5451 6934 5485
rect 6968 5468 7002 5489
rect 6800 5417 6834 5434
rect 6968 5417 7002 5434
rect 6800 5383 7002 5417
rect 7052 5468 7172 5489
rect 7086 5434 7172 5468
rect 7225 5481 7291 5523
rect 7225 5447 7241 5481
rect 7275 5447 7291 5481
rect 7052 5413 7172 5434
rect 7325 5445 7377 5489
rect 7052 5387 7291 5413
rect 7052 5353 7054 5387
rect 7088 5379 7291 5387
rect 7088 5353 7100 5379
rect 6302 5349 6401 5353
rect 6080 5291 6095 5325
rect 6046 5275 6095 5291
rect 6129 5319 6145 5333
rect 6129 5285 6130 5319
rect 6179 5299 6217 5333
rect 6302 5315 6385 5349
rect 6419 5315 6435 5349
rect 6469 5315 6485 5349
rect 6519 5319 6544 5349
rect 6164 5285 6217 5299
rect 6469 5285 6498 5315
rect 6532 5285 6544 5319
rect 6603 5290 6836 5347
rect 7257 5341 7291 5379
rect 7359 5411 7377 5445
rect 7325 5374 7377 5411
rect 5946 5205 6026 5243
rect 5946 5171 5992 5205
rect 5946 5115 6026 5171
rect 6061 5153 6095 5275
rect 6183 5221 6222 5251
rect 6183 5187 6217 5221
rect 6256 5217 6267 5251
rect 6603 5237 6637 5290
rect 6251 5187 6267 5217
rect 6313 5221 6570 5237
rect 6347 5203 6570 5221
rect 6604 5203 6637 5237
rect 6682 5251 6754 5253
rect 6716 5237 6754 5251
rect 6682 5203 6687 5217
rect 6721 5203 6754 5237
rect 6347 5187 6363 5203
rect 6682 5187 6754 5203
rect 6802 5221 6836 5290
rect 6870 5319 6948 5334
rect 7146 5325 7212 5341
rect 7146 5319 7178 5325
rect 6904 5318 6948 5319
rect 6904 5285 6914 5318
rect 6870 5284 6914 5285
rect 6870 5268 6948 5284
rect 6986 5285 7010 5319
rect 7044 5285 7060 5319
rect 7180 5285 7212 5291
rect 6986 5221 7020 5285
rect 7178 5275 7212 5285
rect 7257 5325 7308 5341
rect 7257 5291 7274 5325
rect 7257 5275 7308 5291
rect 6802 5187 7020 5221
rect 7088 5217 7134 5251
rect 7054 5214 7134 5217
rect 7257 5215 7291 5275
rect 7342 5243 7377 5374
rect 6313 5184 6363 5187
rect 6061 5119 6194 5153
rect 6313 5150 6320 5184
rect 6354 5150 6363 5184
rect 7054 5180 7100 5214
rect 7054 5164 7134 5180
rect 6313 5149 6363 5150
rect 5946 5081 5992 5115
rect 6160 5115 6194 5119
rect 6444 5119 6646 5153
rect 6160 5097 6377 5115
rect 5946 5047 6026 5081
rect 6060 5051 6076 5085
rect 6110 5051 6126 5085
rect 6060 5013 6126 5051
rect 6160 5063 6343 5097
rect 6160 5047 6377 5063
rect 6444 5102 6478 5119
rect 6612 5102 6646 5119
rect 6444 5047 6478 5068
rect 6512 5051 6528 5085
rect 6562 5051 6578 5085
rect 6512 5013 6578 5051
rect 6787 5119 7002 5153
rect 7173 5151 7291 5215
rect 7325 5202 7377 5243
rect 7359 5178 7377 5202
rect 7173 5127 7207 5151
rect 6787 5102 6834 5119
rect 6612 5047 6646 5068
rect 6680 5055 6696 5089
rect 6730 5055 6746 5089
rect 6680 5013 6746 5055
rect 6787 5068 6800 5102
rect 6968 5102 7002 5119
rect 6787 5047 6834 5068
rect 6868 5051 6884 5085
rect 6918 5051 6934 5085
rect 6868 5013 6934 5051
rect 6968 5047 7002 5068
rect 7052 5102 7207 5127
rect 7325 5142 7336 5168
rect 7370 5142 7377 5178
rect 7086 5068 7207 5102
rect 7052 5047 7207 5068
rect 7241 5093 7291 5110
rect 7275 5059 7291 5093
rect 7241 5013 7291 5059
rect 7325 5108 7377 5142
rect 7359 5074 7377 5108
rect 7325 5047 7377 5074
rect 7948 5451 8028 5495
rect 8077 5491 8143 5529
rect 8077 5457 8093 5491
rect 8127 5457 8143 5491
rect 8177 5479 8379 5495
rect 7948 5417 7994 5451
rect 8177 5445 8345 5479
rect 8177 5423 8211 5445
rect 8345 5427 8379 5445
rect 8446 5474 8480 5495
rect 8514 5491 8580 5529
rect 8514 5457 8530 5491
rect 8564 5457 8580 5491
rect 8614 5474 8648 5495
rect 7948 5384 8028 5417
rect 8063 5389 8211 5423
rect 8446 5423 8480 5440
rect 8682 5482 8748 5529
rect 8682 5448 8698 5482
rect 8732 5448 8748 5482
rect 8802 5474 8836 5495
rect 8614 5423 8648 5440
rect 7948 5249 8014 5384
rect 8063 5347 8097 5389
rect 8048 5331 8097 5347
rect 8304 5359 8316 5393
rect 8350 5359 8403 5393
rect 8446 5389 8648 5423
rect 8870 5491 8936 5529
rect 8870 5457 8886 5491
rect 8920 5457 8936 5491
rect 8970 5474 9004 5495
rect 8802 5423 8836 5440
rect 8970 5423 9004 5440
rect 8802 5389 9004 5423
rect 9054 5474 9174 5495
rect 9088 5440 9174 5474
rect 9227 5487 9293 5529
rect 10042 5509 10088 5543
rect 10256 5543 10290 5547
rect 10540 5547 10742 5581
rect 10256 5525 10473 5543
rect 9227 5453 9243 5487
rect 9277 5453 9293 5487
rect 9054 5419 9174 5440
rect 9327 5451 9379 5495
rect 10042 5475 10122 5509
rect 10156 5479 10172 5513
rect 10206 5479 10222 5513
rect 9054 5393 9293 5419
rect 9054 5359 9056 5393
rect 9090 5385 9293 5393
rect 9090 5359 9102 5385
rect 8304 5355 8403 5359
rect 8082 5297 8097 5331
rect 8048 5281 8097 5297
rect 8131 5325 8147 5339
rect 8131 5291 8132 5325
rect 8181 5305 8219 5339
rect 8304 5321 8387 5355
rect 8421 5321 8437 5355
rect 8471 5321 8487 5355
rect 8521 5325 8546 5355
rect 8166 5291 8219 5305
rect 8471 5291 8500 5321
rect 8534 5291 8546 5325
rect 8605 5296 8838 5353
rect 9259 5347 9293 5385
rect 9361 5417 9379 5451
rect 10156 5441 10222 5479
rect 10256 5491 10439 5525
rect 10256 5475 10473 5491
rect 10540 5530 10574 5547
rect 10708 5530 10742 5547
rect 10540 5475 10574 5496
rect 10608 5479 10624 5513
rect 10658 5479 10674 5513
rect 10608 5441 10674 5479
rect 10883 5547 11098 5581
rect 11269 5579 11387 5643
rect 11421 5630 11473 5671
rect 11455 5606 11473 5630
rect 11269 5555 11303 5579
rect 10883 5530 10930 5547
rect 10708 5475 10742 5496
rect 10776 5483 10792 5517
rect 10826 5483 10842 5517
rect 10776 5441 10842 5483
rect 10883 5496 10896 5530
rect 11064 5530 11098 5547
rect 10883 5475 10930 5496
rect 10964 5479 10980 5513
rect 11014 5479 11030 5513
rect 10964 5441 11030 5479
rect 11064 5475 11098 5496
rect 11148 5530 11303 5555
rect 11421 5570 11426 5596
rect 11466 5570 11473 5606
rect 11182 5496 11303 5530
rect 11148 5475 11303 5496
rect 11337 5521 11387 5538
rect 11371 5487 11387 5521
rect 11337 5441 11387 5487
rect 11421 5536 11473 5570
rect 11455 5502 11473 5536
rect 11421 5475 11473 5502
rect 12104 5861 12184 5905
rect 12233 5901 12299 5939
rect 12233 5867 12249 5901
rect 12283 5867 12299 5901
rect 12333 5889 12535 5905
rect 12104 5827 12150 5861
rect 12333 5855 12501 5889
rect 12333 5833 12367 5855
rect 12501 5837 12535 5855
rect 12602 5884 12636 5905
rect 12670 5901 12736 5939
rect 12670 5867 12686 5901
rect 12720 5867 12736 5901
rect 12770 5884 12804 5905
rect 12104 5794 12184 5827
rect 12219 5799 12367 5833
rect 12602 5833 12636 5850
rect 12838 5892 12904 5939
rect 12838 5858 12854 5892
rect 12888 5858 12904 5892
rect 12958 5884 12992 5905
rect 12770 5833 12804 5850
rect 12104 5659 12170 5794
rect 12219 5757 12253 5799
rect 12204 5741 12253 5757
rect 12460 5769 12472 5803
rect 12506 5769 12559 5803
rect 12602 5799 12804 5833
rect 13026 5901 13092 5939
rect 13026 5867 13042 5901
rect 13076 5867 13092 5901
rect 13126 5884 13160 5905
rect 12958 5833 12992 5850
rect 13126 5833 13160 5850
rect 12958 5799 13160 5833
rect 13210 5884 13330 5905
rect 13244 5850 13330 5884
rect 13383 5897 13449 5939
rect 13383 5863 13399 5897
rect 13433 5863 13449 5897
rect 13210 5829 13330 5850
rect 13483 5861 13535 5905
rect 13210 5803 13449 5829
rect 13210 5769 13212 5803
rect 13246 5795 13449 5803
rect 13246 5769 13258 5795
rect 12460 5765 12559 5769
rect 12238 5707 12253 5741
rect 12204 5691 12253 5707
rect 12287 5735 12303 5749
rect 12287 5701 12288 5735
rect 12337 5715 12375 5749
rect 12460 5731 12543 5765
rect 12577 5731 12593 5765
rect 12627 5731 12643 5765
rect 12677 5735 12702 5765
rect 12322 5701 12375 5715
rect 12627 5701 12656 5731
rect 12690 5701 12702 5735
rect 12761 5706 12994 5763
rect 13415 5757 13449 5795
rect 13517 5827 13535 5861
rect 13483 5790 13535 5827
rect 12104 5621 12184 5659
rect 12104 5587 12150 5621
rect 12104 5531 12184 5587
rect 12219 5569 12253 5691
rect 12341 5637 12380 5667
rect 12341 5603 12375 5637
rect 12414 5633 12425 5667
rect 12761 5653 12795 5706
rect 12409 5603 12425 5633
rect 12471 5637 12728 5653
rect 12505 5619 12728 5637
rect 12762 5619 12795 5653
rect 12840 5667 12912 5669
rect 12874 5653 12912 5667
rect 12840 5619 12845 5633
rect 12879 5619 12912 5653
rect 12505 5603 12521 5619
rect 12840 5603 12912 5619
rect 12960 5637 12994 5706
rect 13028 5735 13106 5750
rect 13304 5741 13370 5757
rect 13304 5735 13336 5741
rect 13062 5734 13106 5735
rect 13062 5701 13072 5734
rect 13028 5700 13072 5701
rect 13028 5684 13106 5700
rect 13144 5701 13168 5735
rect 13202 5701 13218 5735
rect 13338 5701 13370 5707
rect 13144 5637 13178 5701
rect 13336 5691 13370 5701
rect 13415 5741 13466 5757
rect 13415 5707 13432 5741
rect 13415 5691 13466 5707
rect 12960 5603 13178 5637
rect 13246 5633 13292 5667
rect 13212 5630 13292 5633
rect 13415 5631 13449 5691
rect 13500 5659 13535 5790
rect 12471 5600 12521 5603
rect 12219 5535 12352 5569
rect 12471 5566 12478 5600
rect 12512 5566 12521 5600
rect 13212 5596 13258 5630
rect 13212 5580 13292 5596
rect 12471 5565 12521 5566
rect 12104 5497 12150 5531
rect 12318 5531 12352 5535
rect 12602 5535 12804 5569
rect 12318 5513 12535 5531
rect 12104 5463 12184 5497
rect 12218 5467 12234 5501
rect 12268 5467 12284 5501
rect 9327 5380 9379 5417
rect 10018 5407 10047 5441
rect 10081 5407 10139 5441
rect 10173 5407 10231 5441
rect 10265 5407 10323 5441
rect 10357 5407 10415 5441
rect 10449 5407 10507 5441
rect 10541 5407 10599 5441
rect 10633 5407 10691 5441
rect 10725 5407 10783 5441
rect 10817 5407 10875 5441
rect 10909 5407 10967 5441
rect 11001 5407 11059 5441
rect 11093 5407 11151 5441
rect 11185 5407 11243 5441
rect 11277 5407 11335 5441
rect 11369 5407 11427 5441
rect 11461 5407 11490 5441
rect 12218 5429 12284 5467
rect 12318 5479 12501 5513
rect 12318 5463 12535 5479
rect 12602 5518 12636 5535
rect 12770 5518 12804 5535
rect 12602 5463 12636 5484
rect 12670 5467 12686 5501
rect 12720 5467 12736 5501
rect 12670 5429 12736 5467
rect 12945 5535 13160 5569
rect 13331 5567 13449 5631
rect 13483 5618 13535 5659
rect 13517 5594 13535 5618
rect 13331 5543 13365 5567
rect 12945 5518 12992 5535
rect 12770 5463 12804 5484
rect 12838 5471 12854 5505
rect 12888 5471 12904 5505
rect 12838 5429 12904 5471
rect 12945 5484 12958 5518
rect 13126 5518 13160 5535
rect 12945 5463 12992 5484
rect 13026 5467 13042 5501
rect 13076 5467 13092 5501
rect 13026 5429 13092 5467
rect 13126 5463 13160 5484
rect 13210 5518 13365 5543
rect 13483 5558 13494 5584
rect 13528 5558 13535 5594
rect 13244 5484 13365 5518
rect 13210 5463 13365 5484
rect 13399 5509 13449 5526
rect 13433 5475 13449 5509
rect 13399 5429 13449 5475
rect 13483 5524 13535 5558
rect 13517 5490 13535 5524
rect 13483 5463 13535 5490
rect 14062 5869 14142 5913
rect 14191 5909 14257 5947
rect 14191 5875 14207 5909
rect 14241 5875 14257 5909
rect 14291 5897 14493 5913
rect 14062 5835 14108 5869
rect 14291 5863 14459 5897
rect 14291 5841 14325 5863
rect 14459 5845 14493 5863
rect 14560 5892 14594 5913
rect 14628 5909 14694 5947
rect 14628 5875 14644 5909
rect 14678 5875 14694 5909
rect 14728 5892 14762 5913
rect 14062 5802 14142 5835
rect 14177 5807 14325 5841
rect 14560 5841 14594 5858
rect 14796 5900 14862 5947
rect 14796 5866 14812 5900
rect 14846 5866 14862 5900
rect 14916 5892 14950 5913
rect 14728 5841 14762 5858
rect 14062 5667 14128 5802
rect 14177 5765 14211 5807
rect 14162 5749 14211 5765
rect 14418 5777 14430 5811
rect 14464 5777 14517 5811
rect 14560 5807 14762 5841
rect 14984 5909 15050 5947
rect 14984 5875 15000 5909
rect 15034 5875 15050 5909
rect 15084 5892 15118 5913
rect 14916 5841 14950 5858
rect 15084 5841 15118 5858
rect 14916 5807 15118 5841
rect 15168 5892 15288 5913
rect 15202 5858 15288 5892
rect 15341 5905 15407 5947
rect 15341 5871 15357 5905
rect 15391 5871 15407 5905
rect 15168 5837 15288 5858
rect 15441 5869 15493 5913
rect 15168 5811 15407 5837
rect 15168 5777 15170 5811
rect 15204 5803 15407 5811
rect 15204 5777 15216 5803
rect 14418 5773 14517 5777
rect 14196 5715 14211 5749
rect 14162 5699 14211 5715
rect 14245 5743 14261 5757
rect 14245 5709 14246 5743
rect 14295 5723 14333 5757
rect 14418 5739 14501 5773
rect 14535 5739 14551 5773
rect 14585 5739 14601 5773
rect 14635 5743 14660 5773
rect 14280 5709 14333 5723
rect 14585 5709 14614 5739
rect 14648 5709 14660 5743
rect 14719 5714 14952 5771
rect 15373 5765 15407 5803
rect 15475 5835 15493 5869
rect 15441 5798 15493 5835
rect 14062 5629 14142 5667
rect 14062 5595 14108 5629
rect 14062 5539 14142 5595
rect 14177 5577 14211 5699
rect 14299 5645 14338 5675
rect 14299 5611 14333 5645
rect 14372 5641 14383 5675
rect 14719 5661 14753 5714
rect 14367 5611 14383 5641
rect 14429 5645 14686 5661
rect 14463 5627 14686 5645
rect 14720 5627 14753 5661
rect 14798 5675 14870 5677
rect 14832 5661 14870 5675
rect 14798 5627 14803 5641
rect 14837 5627 14870 5661
rect 14463 5611 14479 5627
rect 14798 5611 14870 5627
rect 14918 5645 14952 5714
rect 14986 5743 15064 5758
rect 15262 5749 15328 5765
rect 15262 5743 15294 5749
rect 15020 5742 15064 5743
rect 15020 5709 15030 5742
rect 14986 5708 15030 5709
rect 14986 5692 15064 5708
rect 15102 5709 15126 5743
rect 15160 5709 15176 5743
rect 15296 5709 15328 5715
rect 15102 5645 15136 5709
rect 15294 5699 15328 5709
rect 15373 5749 15424 5765
rect 15373 5715 15390 5749
rect 15373 5699 15424 5715
rect 14918 5611 15136 5645
rect 15204 5641 15250 5675
rect 15170 5638 15250 5641
rect 15373 5639 15407 5699
rect 15458 5667 15493 5798
rect 14429 5608 14479 5611
rect 14177 5543 14310 5577
rect 14429 5574 14436 5608
rect 14470 5574 14479 5608
rect 15170 5604 15216 5638
rect 15170 5588 15250 5604
rect 14429 5573 14479 5574
rect 14062 5505 14108 5539
rect 14276 5539 14310 5543
rect 14560 5543 14762 5577
rect 14276 5521 14493 5539
rect 14062 5471 14142 5505
rect 14176 5475 14192 5509
rect 14226 5475 14242 5509
rect 14176 5437 14242 5475
rect 14276 5487 14459 5521
rect 14276 5471 14493 5487
rect 14560 5526 14594 5543
rect 14728 5526 14762 5543
rect 14560 5471 14594 5492
rect 14628 5475 14644 5509
rect 14678 5475 14694 5509
rect 14628 5437 14694 5475
rect 14903 5543 15118 5577
rect 15289 5575 15407 5639
rect 15441 5626 15493 5667
rect 15475 5602 15493 5626
rect 15289 5551 15323 5575
rect 14903 5526 14950 5543
rect 14728 5471 14762 5492
rect 14796 5479 14812 5513
rect 14846 5479 14862 5513
rect 14796 5437 14862 5479
rect 14903 5492 14916 5526
rect 15084 5526 15118 5543
rect 14903 5471 14950 5492
rect 14984 5475 15000 5509
rect 15034 5475 15050 5509
rect 14984 5437 15050 5475
rect 15084 5471 15118 5492
rect 15168 5526 15323 5551
rect 15441 5566 15452 5592
rect 15486 5566 15493 5602
rect 15202 5492 15323 5526
rect 15168 5471 15323 5492
rect 15357 5517 15407 5534
rect 15391 5483 15407 5517
rect 15357 5437 15407 5483
rect 15441 5532 15493 5566
rect 15475 5498 15493 5532
rect 15441 5471 15493 5498
rect 16056 5875 16136 5919
rect 16185 5915 16251 5953
rect 16185 5881 16201 5915
rect 16235 5881 16251 5915
rect 16285 5903 16487 5919
rect 16056 5841 16102 5875
rect 16285 5869 16453 5903
rect 16285 5847 16319 5869
rect 16453 5851 16487 5869
rect 16554 5898 16588 5919
rect 16622 5915 16688 5953
rect 16622 5881 16638 5915
rect 16672 5881 16688 5915
rect 16722 5898 16756 5919
rect 16056 5808 16136 5841
rect 16171 5813 16319 5847
rect 16554 5847 16588 5864
rect 16790 5906 16856 5953
rect 16790 5872 16806 5906
rect 16840 5872 16856 5906
rect 16910 5898 16944 5919
rect 16722 5847 16756 5864
rect 16056 5673 16122 5808
rect 16171 5771 16205 5813
rect 16156 5755 16205 5771
rect 16412 5783 16424 5817
rect 16458 5783 16511 5817
rect 16554 5813 16756 5847
rect 16978 5915 17044 5953
rect 16978 5881 16994 5915
rect 17028 5881 17044 5915
rect 17078 5898 17112 5919
rect 16910 5847 16944 5864
rect 17078 5847 17112 5864
rect 16910 5813 17112 5847
rect 17162 5898 17282 5919
rect 17196 5864 17282 5898
rect 17335 5911 17401 5953
rect 17335 5877 17351 5911
rect 17385 5877 17401 5911
rect 17162 5843 17282 5864
rect 17435 5875 17487 5919
rect 17162 5817 17401 5843
rect 17162 5783 17164 5817
rect 17198 5809 17401 5817
rect 17198 5783 17210 5809
rect 16412 5779 16511 5783
rect 16190 5721 16205 5755
rect 16156 5705 16205 5721
rect 16239 5749 16255 5763
rect 16239 5715 16240 5749
rect 16289 5729 16327 5763
rect 16412 5745 16495 5779
rect 16529 5745 16545 5779
rect 16579 5745 16595 5779
rect 16629 5749 16654 5779
rect 16274 5715 16327 5729
rect 16579 5715 16608 5745
rect 16642 5715 16654 5749
rect 16713 5720 16946 5777
rect 17367 5771 17401 5809
rect 17469 5841 17487 5875
rect 17435 5804 17487 5841
rect 16056 5635 16136 5673
rect 16056 5601 16102 5635
rect 16056 5545 16136 5601
rect 16171 5583 16205 5705
rect 16293 5651 16332 5681
rect 16293 5617 16327 5651
rect 16366 5647 16377 5681
rect 16713 5667 16747 5720
rect 16361 5617 16377 5647
rect 16423 5651 16680 5667
rect 16457 5633 16680 5651
rect 16714 5633 16747 5667
rect 16792 5681 16864 5683
rect 16826 5667 16864 5681
rect 16792 5633 16797 5647
rect 16831 5633 16864 5667
rect 16457 5617 16473 5633
rect 16792 5617 16864 5633
rect 16912 5651 16946 5720
rect 16980 5749 17058 5764
rect 17256 5755 17322 5771
rect 17256 5749 17288 5755
rect 17014 5748 17058 5749
rect 17014 5715 17024 5748
rect 16980 5714 17024 5715
rect 16980 5698 17058 5714
rect 17096 5715 17120 5749
rect 17154 5715 17170 5749
rect 17290 5715 17322 5721
rect 17096 5651 17130 5715
rect 17288 5705 17322 5715
rect 17367 5755 17418 5771
rect 17367 5721 17384 5755
rect 17367 5705 17418 5721
rect 16912 5617 17130 5651
rect 17198 5647 17244 5681
rect 17164 5644 17244 5647
rect 17367 5645 17401 5705
rect 17452 5673 17487 5804
rect 16423 5614 16473 5617
rect 16171 5549 16304 5583
rect 16423 5580 16430 5614
rect 16464 5580 16473 5614
rect 17164 5610 17210 5644
rect 17164 5594 17244 5610
rect 16423 5579 16473 5580
rect 16056 5511 16102 5545
rect 16270 5545 16304 5549
rect 16554 5549 16756 5583
rect 16270 5527 16487 5545
rect 16056 5477 16136 5511
rect 16170 5481 16186 5515
rect 16220 5481 16236 5515
rect 16170 5443 16236 5481
rect 16270 5493 16453 5527
rect 16270 5477 16487 5493
rect 16554 5532 16588 5549
rect 16722 5532 16756 5549
rect 16554 5477 16588 5498
rect 16622 5481 16638 5515
rect 16672 5481 16688 5515
rect 16622 5443 16688 5481
rect 16897 5549 17112 5583
rect 17283 5581 17401 5645
rect 17435 5632 17487 5673
rect 17469 5608 17487 5632
rect 17283 5557 17317 5581
rect 16897 5532 16944 5549
rect 16722 5477 16756 5498
rect 16790 5485 16806 5519
rect 16840 5485 16856 5519
rect 16790 5443 16856 5485
rect 16897 5498 16910 5532
rect 17078 5532 17112 5549
rect 16897 5477 16944 5498
rect 16978 5481 16994 5515
rect 17028 5481 17044 5515
rect 16978 5443 17044 5481
rect 17078 5477 17112 5498
rect 17162 5532 17317 5557
rect 17435 5572 17446 5598
rect 17480 5572 17487 5608
rect 17196 5498 17317 5532
rect 17162 5477 17317 5498
rect 17351 5523 17401 5540
rect 17385 5489 17401 5523
rect 17351 5443 17401 5489
rect 17435 5538 17487 5572
rect 17469 5504 17487 5538
rect 17435 5477 17487 5504
rect 12080 5395 12109 5429
rect 12143 5395 12201 5429
rect 12235 5395 12293 5429
rect 12327 5395 12385 5429
rect 12419 5395 12477 5429
rect 12511 5395 12569 5429
rect 12603 5395 12661 5429
rect 12695 5395 12753 5429
rect 12787 5395 12845 5429
rect 12879 5395 12937 5429
rect 12971 5395 13029 5429
rect 13063 5395 13121 5429
rect 13155 5395 13213 5429
rect 13247 5395 13305 5429
rect 13339 5395 13397 5429
rect 13431 5395 13489 5429
rect 13523 5395 13552 5429
rect 14038 5403 14067 5437
rect 14101 5403 14159 5437
rect 14193 5403 14251 5437
rect 14285 5403 14343 5437
rect 14377 5403 14435 5437
rect 14469 5403 14527 5437
rect 14561 5403 14619 5437
rect 14653 5403 14711 5437
rect 14745 5403 14803 5437
rect 14837 5403 14895 5437
rect 14929 5403 14987 5437
rect 15021 5403 15079 5437
rect 15113 5403 15171 5437
rect 15205 5403 15263 5437
rect 15297 5403 15355 5437
rect 15389 5403 15447 5437
rect 15481 5403 15510 5437
rect 16032 5409 16061 5443
rect 16095 5409 16153 5443
rect 16187 5409 16245 5443
rect 16279 5409 16337 5443
rect 16371 5409 16429 5443
rect 16463 5409 16521 5443
rect 16555 5409 16613 5443
rect 16647 5409 16705 5443
rect 16739 5409 16797 5443
rect 16831 5409 16889 5443
rect 16923 5409 16981 5443
rect 17015 5409 17073 5443
rect 17107 5409 17165 5443
rect 17199 5409 17257 5443
rect 17291 5409 17349 5443
rect 17383 5409 17441 5443
rect 17475 5409 17504 5443
rect 7948 5211 8028 5249
rect 7948 5177 7994 5211
rect 7948 5121 8028 5177
rect 8063 5159 8097 5281
rect 8185 5227 8224 5257
rect 8185 5193 8219 5227
rect 8258 5223 8269 5257
rect 8605 5243 8639 5296
rect 8253 5193 8269 5223
rect 8315 5227 8572 5243
rect 8349 5209 8572 5227
rect 8606 5209 8639 5243
rect 8684 5257 8756 5259
rect 8718 5243 8756 5257
rect 8684 5209 8689 5223
rect 8723 5209 8756 5243
rect 8349 5193 8365 5209
rect 8684 5193 8756 5209
rect 8804 5227 8838 5296
rect 8872 5325 8950 5340
rect 9148 5331 9214 5347
rect 9148 5325 9180 5331
rect 8906 5324 8950 5325
rect 8906 5291 8916 5324
rect 8872 5290 8916 5291
rect 8872 5274 8950 5290
rect 8988 5291 9012 5325
rect 9046 5291 9062 5325
rect 9182 5291 9214 5297
rect 8988 5227 9022 5291
rect 9180 5281 9214 5291
rect 9259 5331 9310 5347
rect 9259 5297 9276 5331
rect 9259 5281 9310 5297
rect 8804 5193 9022 5227
rect 9090 5223 9136 5257
rect 9056 5220 9136 5223
rect 9259 5221 9293 5281
rect 9344 5249 9379 5380
rect 8315 5190 8365 5193
rect 8063 5125 8196 5159
rect 8315 5156 8322 5190
rect 8356 5156 8365 5190
rect 9056 5186 9102 5220
rect 9056 5170 9136 5186
rect 8315 5155 8365 5156
rect 7948 5087 7994 5121
rect 8162 5121 8196 5125
rect 8446 5125 8648 5159
rect 8162 5103 8379 5121
rect 7948 5053 8028 5087
rect 8062 5057 8078 5091
rect 8112 5057 8128 5091
rect 8062 5019 8128 5057
rect 8162 5069 8345 5103
rect 8162 5053 8379 5069
rect 8446 5108 8480 5125
rect 8614 5108 8648 5125
rect 8446 5053 8480 5074
rect 8514 5057 8530 5091
rect 8564 5057 8580 5091
rect 8514 5019 8580 5057
rect 8789 5125 9004 5159
rect 9175 5157 9293 5221
rect 9327 5208 9379 5249
rect 9361 5184 9379 5208
rect 9175 5133 9209 5157
rect 8789 5108 8836 5125
rect 8614 5053 8648 5074
rect 8682 5061 8698 5095
rect 8732 5061 8748 5095
rect 8682 5019 8748 5061
rect 8789 5074 8802 5108
rect 8970 5108 9004 5125
rect 8789 5053 8836 5074
rect 8870 5057 8886 5091
rect 8920 5057 8936 5091
rect 8870 5019 8936 5057
rect 8970 5053 9004 5074
rect 9054 5108 9209 5133
rect 9327 5148 9338 5174
rect 9372 5148 9379 5184
rect 9088 5074 9209 5108
rect 9054 5053 9209 5074
rect 9243 5099 9293 5116
rect 9277 5065 9293 5099
rect 9243 5019 9293 5065
rect 9327 5114 9379 5148
rect 9361 5080 9379 5114
rect 9327 5053 9379 5080
rect 10046 5077 10075 5111
rect 10109 5077 10167 5111
rect 10201 5077 10259 5111
rect 10293 5077 10351 5111
rect 10385 5077 10443 5111
rect 10477 5077 10535 5111
rect 10569 5077 10627 5111
rect 10661 5077 10719 5111
rect 10753 5077 10811 5111
rect 10845 5077 10903 5111
rect 10937 5077 10995 5111
rect 11029 5077 11087 5111
rect 11121 5077 11179 5111
rect 11213 5077 11271 5111
rect 11305 5077 11363 5111
rect 11397 5077 11455 5111
rect 11489 5077 11518 5111
rect 3970 4979 3999 5013
rect 4033 4979 4091 5013
rect 4125 4979 4183 5013
rect 4217 4979 4275 5013
rect 4309 4979 4367 5013
rect 4401 4979 4459 5013
rect 4493 4979 4551 5013
rect 4585 4979 4643 5013
rect 4677 4979 4735 5013
rect 4769 4979 4827 5013
rect 4861 4979 4919 5013
rect 4953 4979 5011 5013
rect 5045 4979 5103 5013
rect 5137 4979 5195 5013
rect 5229 4979 5287 5013
rect 5321 4979 5379 5013
rect 5413 4979 5442 5013
rect 5922 4979 5951 5013
rect 5985 4979 6043 5013
rect 6077 4979 6135 5013
rect 6169 4979 6227 5013
rect 6261 4979 6319 5013
rect 6353 4979 6411 5013
rect 6445 4979 6503 5013
rect 6537 4979 6595 5013
rect 6629 4979 6687 5013
rect 6721 4979 6779 5013
rect 6813 4979 6871 5013
rect 6905 4979 6963 5013
rect 6997 4979 7055 5013
rect 7089 4979 7147 5013
rect 7181 4979 7239 5013
rect 7273 4979 7331 5013
rect 7365 4979 7394 5013
rect 7924 4985 7953 5019
rect 7987 4985 8045 5019
rect 8079 4985 8137 5019
rect 8171 4985 8229 5019
rect 8263 4985 8321 5019
rect 8355 4985 8413 5019
rect 8447 4985 8505 5019
rect 8539 4985 8597 5019
rect 8631 4985 8689 5019
rect 8723 4985 8781 5019
rect 8815 4985 8873 5019
rect 8907 4985 8965 5019
rect 8999 4985 9057 5019
rect 9091 4985 9149 5019
rect 9183 4985 9241 5019
rect 9275 4985 9333 5019
rect 9367 4985 9396 5019
rect 10070 4999 10150 5043
rect 10199 5039 10265 5077
rect 10199 5005 10215 5039
rect 10249 5005 10265 5039
rect 10299 5027 10501 5043
rect 10070 4965 10116 4999
rect 10299 4993 10467 5027
rect 10299 4971 10333 4993
rect 10467 4975 10501 4993
rect 10568 5022 10602 5043
rect 10636 5039 10702 5077
rect 10636 5005 10652 5039
rect 10686 5005 10702 5039
rect 10736 5022 10770 5043
rect 10070 4932 10150 4965
rect 10185 4937 10333 4971
rect 10568 4971 10602 4988
rect 10804 5030 10870 5077
rect 10804 4996 10820 5030
rect 10854 4996 10870 5030
rect 10924 5022 10958 5043
rect 10736 4971 10770 4988
rect 10070 4797 10136 4932
rect 10185 4895 10219 4937
rect 10170 4879 10219 4895
rect 10426 4907 10438 4941
rect 10472 4907 10525 4941
rect 10568 4937 10770 4971
rect 10992 5039 11058 5077
rect 10992 5005 11008 5039
rect 11042 5005 11058 5039
rect 11092 5022 11126 5043
rect 10924 4971 10958 4988
rect 11092 4971 11126 4988
rect 10924 4937 11126 4971
rect 11176 5022 11296 5043
rect 11210 4988 11296 5022
rect 11349 5035 11415 5077
rect 11349 5001 11365 5035
rect 11399 5001 11415 5035
rect 11176 4967 11296 4988
rect 11449 4999 11501 5043
rect 12316 5033 12345 5067
rect 12379 5033 12437 5067
rect 12471 5033 12529 5067
rect 12563 5033 12621 5067
rect 12655 5033 12713 5067
rect 12747 5033 12805 5067
rect 12839 5033 12897 5067
rect 12931 5033 12989 5067
rect 13023 5033 13081 5067
rect 13115 5033 13173 5067
rect 13207 5033 13265 5067
rect 13299 5033 13357 5067
rect 13391 5033 13449 5067
rect 13483 5033 13541 5067
rect 13575 5033 13633 5067
rect 13667 5033 13725 5067
rect 13759 5033 13788 5067
rect 11176 4941 11415 4967
rect 11176 4907 11178 4941
rect 11212 4933 11415 4941
rect 11212 4907 11224 4933
rect 10426 4903 10525 4907
rect 10204 4845 10219 4879
rect 10170 4829 10219 4845
rect 10253 4873 10269 4887
rect 10253 4839 10254 4873
rect 10303 4853 10341 4887
rect 10426 4869 10509 4903
rect 10543 4869 10559 4903
rect 10593 4869 10609 4903
rect 10643 4873 10668 4903
rect 10288 4839 10341 4853
rect 10593 4839 10622 4869
rect 10656 4839 10668 4873
rect 10727 4844 10960 4901
rect 11381 4895 11415 4933
rect 11483 4965 11501 4999
rect 11449 4928 11501 4965
rect 10070 4759 10150 4797
rect 10070 4725 10116 4759
rect 10070 4669 10150 4725
rect 10185 4707 10219 4829
rect 10307 4775 10346 4805
rect 10307 4741 10341 4775
rect 10380 4771 10391 4805
rect 10727 4791 10761 4844
rect 10375 4741 10391 4771
rect 10437 4775 10694 4791
rect 10471 4757 10694 4775
rect 10728 4757 10761 4791
rect 10806 4805 10878 4807
rect 10840 4791 10878 4805
rect 10806 4757 10811 4771
rect 10845 4757 10878 4791
rect 10471 4741 10487 4757
rect 10806 4741 10878 4757
rect 10926 4775 10960 4844
rect 10994 4873 11072 4888
rect 11270 4879 11336 4895
rect 11270 4873 11302 4879
rect 11028 4872 11072 4873
rect 11028 4839 11038 4872
rect 10994 4838 11038 4839
rect 10994 4822 11072 4838
rect 11110 4839 11134 4873
rect 11168 4839 11184 4873
rect 11304 4839 11336 4845
rect 11110 4775 11144 4839
rect 11302 4829 11336 4839
rect 11381 4879 11432 4895
rect 11381 4845 11398 4879
rect 11381 4829 11432 4845
rect 10926 4741 11144 4775
rect 11212 4771 11258 4805
rect 11178 4768 11258 4771
rect 11381 4769 11415 4829
rect 11466 4797 11501 4928
rect 10437 4740 10487 4741
rect 10185 4673 10318 4707
rect 10437 4706 10446 4740
rect 10480 4706 10487 4740
rect 11178 4734 11224 4768
rect 11178 4718 11258 4734
rect 10437 4703 10487 4706
rect 10070 4635 10116 4669
rect 10284 4669 10318 4673
rect 10568 4673 10770 4707
rect 10284 4651 10501 4669
rect 10070 4601 10150 4635
rect 10184 4605 10200 4639
rect 10234 4605 10250 4639
rect 10184 4567 10250 4605
rect 10284 4617 10467 4651
rect 10284 4601 10501 4617
rect 10568 4656 10602 4673
rect 10736 4656 10770 4673
rect 10568 4601 10602 4622
rect 10636 4605 10652 4639
rect 10686 4605 10702 4639
rect 10636 4567 10702 4605
rect 10911 4673 11126 4707
rect 11297 4705 11415 4769
rect 11449 4756 11501 4797
rect 11483 4732 11501 4756
rect 11297 4681 11331 4705
rect 10911 4656 10958 4673
rect 10736 4601 10770 4622
rect 10804 4609 10820 4643
rect 10854 4609 10870 4643
rect 10804 4567 10870 4609
rect 10911 4622 10924 4656
rect 11092 4656 11126 4673
rect 10911 4601 10958 4622
rect 10992 4605 11008 4639
rect 11042 4605 11058 4639
rect 10992 4567 11058 4605
rect 11092 4601 11126 4622
rect 11176 4656 11331 4681
rect 11449 4696 11454 4722
rect 11494 4696 11501 4732
rect 11210 4622 11331 4656
rect 11176 4601 11331 4622
rect 11365 4647 11415 4664
rect 11399 4613 11415 4647
rect 11365 4567 11415 4613
rect 11449 4662 11501 4696
rect 11483 4628 11501 4662
rect 11449 4601 11501 4628
rect 12340 4955 12420 4999
rect 12469 4995 12535 5033
rect 12469 4961 12485 4995
rect 12519 4961 12535 4995
rect 12569 4983 12771 4999
rect 12340 4921 12386 4955
rect 12569 4949 12737 4983
rect 12569 4927 12603 4949
rect 12737 4931 12771 4949
rect 12838 4978 12872 4999
rect 12906 4995 12972 5033
rect 12906 4961 12922 4995
rect 12956 4961 12972 4995
rect 13006 4978 13040 4999
rect 12340 4888 12420 4921
rect 12455 4893 12603 4927
rect 12838 4927 12872 4944
rect 13074 4986 13140 5033
rect 13074 4952 13090 4986
rect 13124 4952 13140 4986
rect 13194 4978 13228 4999
rect 13006 4927 13040 4944
rect 12340 4753 12406 4888
rect 12455 4851 12489 4893
rect 12440 4835 12489 4851
rect 12696 4863 12708 4897
rect 12742 4863 12795 4897
rect 12838 4893 13040 4927
rect 13262 4995 13328 5033
rect 13262 4961 13278 4995
rect 13312 4961 13328 4995
rect 13362 4978 13396 4999
rect 13194 4927 13228 4944
rect 13362 4927 13396 4944
rect 13194 4893 13396 4927
rect 13446 4978 13566 4999
rect 13480 4944 13566 4978
rect 13619 4991 13685 5033
rect 14318 5027 14347 5061
rect 14381 5027 14439 5061
rect 14473 5027 14531 5061
rect 14565 5027 14623 5061
rect 14657 5027 14715 5061
rect 14749 5027 14807 5061
rect 14841 5027 14899 5061
rect 14933 5027 14991 5061
rect 15025 5027 15083 5061
rect 15117 5027 15175 5061
rect 15209 5027 15267 5061
rect 15301 5027 15359 5061
rect 15393 5027 15451 5061
rect 15485 5027 15543 5061
rect 15577 5027 15635 5061
rect 15669 5027 15727 5061
rect 15761 5027 15790 5061
rect 13619 4957 13635 4991
rect 13669 4957 13685 4991
rect 13446 4923 13566 4944
rect 13719 4955 13771 4999
rect 13446 4897 13685 4923
rect 13446 4863 13448 4897
rect 13482 4889 13685 4897
rect 13482 4863 13494 4889
rect 12696 4859 12795 4863
rect 12474 4801 12489 4835
rect 12440 4785 12489 4801
rect 12523 4829 12539 4843
rect 12523 4795 12524 4829
rect 12573 4809 12611 4843
rect 12696 4825 12779 4859
rect 12813 4825 12829 4859
rect 12863 4825 12879 4859
rect 12913 4829 12938 4859
rect 12558 4795 12611 4809
rect 12863 4795 12892 4825
rect 12926 4795 12938 4829
rect 12997 4800 13230 4857
rect 13651 4851 13685 4889
rect 13753 4921 13771 4955
rect 13719 4884 13771 4921
rect 12340 4715 12420 4753
rect 12340 4681 12386 4715
rect 12340 4625 12420 4681
rect 12455 4663 12489 4785
rect 12577 4731 12616 4761
rect 12577 4697 12611 4731
rect 12650 4727 12661 4761
rect 12997 4747 13031 4800
rect 12645 4697 12661 4727
rect 12707 4731 12964 4747
rect 12741 4713 12964 4731
rect 12998 4713 13031 4747
rect 13076 4761 13148 4763
rect 13110 4747 13148 4761
rect 13076 4713 13081 4727
rect 13115 4713 13148 4747
rect 12741 4697 12757 4713
rect 13076 4697 13148 4713
rect 13196 4731 13230 4800
rect 13264 4829 13342 4844
rect 13540 4835 13606 4851
rect 13540 4829 13572 4835
rect 13298 4828 13342 4829
rect 13298 4795 13308 4828
rect 13264 4794 13308 4795
rect 13264 4778 13342 4794
rect 13380 4795 13404 4829
rect 13438 4795 13454 4829
rect 13574 4795 13606 4801
rect 13380 4731 13414 4795
rect 13572 4785 13606 4795
rect 13651 4835 13702 4851
rect 13651 4801 13668 4835
rect 13651 4785 13702 4801
rect 13196 4697 13414 4731
rect 13482 4727 13528 4761
rect 13448 4724 13528 4727
rect 13651 4725 13685 4785
rect 13736 4753 13771 4884
rect 12707 4694 12757 4697
rect 12455 4629 12588 4663
rect 12707 4660 12714 4694
rect 12748 4660 12757 4694
rect 13448 4690 13494 4724
rect 13448 4674 13528 4690
rect 12707 4659 12757 4660
rect 12340 4591 12386 4625
rect 12554 4625 12588 4629
rect 12838 4629 13040 4663
rect 12554 4607 12771 4625
rect 10046 4533 10075 4567
rect 10109 4533 10167 4567
rect 10201 4533 10259 4567
rect 10293 4533 10351 4567
rect 10385 4533 10443 4567
rect 10477 4533 10535 4567
rect 10569 4533 10627 4567
rect 10661 4533 10719 4567
rect 10753 4533 10811 4567
rect 10845 4533 10903 4567
rect 10937 4533 10995 4567
rect 11029 4533 11087 4567
rect 11121 4533 11179 4567
rect 11213 4533 11271 4567
rect 11305 4533 11363 4567
rect 11397 4533 11455 4567
rect 11489 4533 11518 4567
rect 12340 4557 12420 4591
rect 12454 4561 12470 4595
rect 12504 4561 12520 4595
rect 12454 4523 12520 4561
rect 12554 4573 12737 4607
rect 12554 4557 12771 4573
rect 12838 4612 12872 4629
rect 13006 4612 13040 4629
rect 12838 4557 12872 4578
rect 12906 4561 12922 4595
rect 12956 4561 12972 4595
rect 12906 4523 12972 4561
rect 13181 4629 13396 4663
rect 13567 4661 13685 4725
rect 13719 4712 13771 4753
rect 13753 4688 13771 4712
rect 13567 4637 13601 4661
rect 13181 4612 13228 4629
rect 13006 4557 13040 4578
rect 13074 4565 13090 4599
rect 13124 4565 13140 4599
rect 13074 4523 13140 4565
rect 13181 4578 13194 4612
rect 13362 4612 13396 4629
rect 13181 4557 13228 4578
rect 13262 4561 13278 4595
rect 13312 4561 13328 4595
rect 13262 4523 13328 4561
rect 13362 4557 13396 4578
rect 13446 4612 13601 4637
rect 13719 4652 13730 4678
rect 13764 4652 13771 4688
rect 13480 4578 13601 4612
rect 13446 4557 13601 4578
rect 13635 4603 13685 4620
rect 13669 4569 13685 4603
rect 13635 4523 13685 4569
rect 13719 4618 13771 4652
rect 13753 4584 13771 4618
rect 13719 4557 13771 4584
rect 14342 4949 14422 4993
rect 14471 4989 14537 5027
rect 14471 4955 14487 4989
rect 14521 4955 14537 4989
rect 14571 4977 14773 4993
rect 14342 4915 14388 4949
rect 14571 4943 14739 4977
rect 14571 4921 14605 4943
rect 14739 4925 14773 4943
rect 14840 4972 14874 4993
rect 14908 4989 14974 5027
rect 14908 4955 14924 4989
rect 14958 4955 14974 4989
rect 15008 4972 15042 4993
rect 14342 4882 14422 4915
rect 14457 4887 14605 4921
rect 14840 4921 14874 4938
rect 15076 4980 15142 5027
rect 15076 4946 15092 4980
rect 15126 4946 15142 4980
rect 15196 4972 15230 4993
rect 15008 4921 15042 4938
rect 14342 4747 14408 4882
rect 14457 4845 14491 4887
rect 14442 4829 14491 4845
rect 14698 4857 14710 4891
rect 14744 4857 14797 4891
rect 14840 4887 15042 4921
rect 15264 4989 15330 5027
rect 15264 4955 15280 4989
rect 15314 4955 15330 4989
rect 15364 4972 15398 4993
rect 15196 4921 15230 4938
rect 15364 4921 15398 4938
rect 15196 4887 15398 4921
rect 15448 4972 15568 4993
rect 15482 4938 15568 4972
rect 15621 4985 15687 5027
rect 16340 5009 16369 5043
rect 16403 5009 16461 5043
rect 16495 5009 16553 5043
rect 16587 5009 16645 5043
rect 16679 5009 16737 5043
rect 16771 5009 16829 5043
rect 16863 5009 16921 5043
rect 16955 5009 17013 5043
rect 17047 5009 17105 5043
rect 17139 5009 17197 5043
rect 17231 5009 17289 5043
rect 17323 5009 17381 5043
rect 17415 5009 17473 5043
rect 17507 5009 17565 5043
rect 17599 5009 17657 5043
rect 17691 5009 17749 5043
rect 17783 5009 17812 5043
rect 15621 4951 15637 4985
rect 15671 4951 15687 4985
rect 15448 4917 15568 4938
rect 15721 4949 15773 4993
rect 15448 4891 15687 4917
rect 15448 4857 15450 4891
rect 15484 4883 15687 4891
rect 15484 4857 15496 4883
rect 14698 4853 14797 4857
rect 14476 4795 14491 4829
rect 14442 4779 14491 4795
rect 14525 4823 14541 4837
rect 14525 4789 14526 4823
rect 14575 4803 14613 4837
rect 14698 4819 14781 4853
rect 14815 4819 14831 4853
rect 14865 4819 14881 4853
rect 14915 4823 14940 4853
rect 14560 4789 14613 4803
rect 14865 4789 14894 4819
rect 14928 4789 14940 4823
rect 14999 4794 15232 4851
rect 15653 4845 15687 4883
rect 15755 4915 15773 4949
rect 15721 4878 15773 4915
rect 14342 4709 14422 4747
rect 14342 4675 14388 4709
rect 14342 4619 14422 4675
rect 14457 4657 14491 4779
rect 14579 4725 14618 4755
rect 14579 4691 14613 4725
rect 14652 4721 14663 4755
rect 14999 4741 15033 4794
rect 14647 4691 14663 4721
rect 14709 4725 14966 4741
rect 14743 4707 14966 4725
rect 15000 4707 15033 4741
rect 15078 4755 15150 4757
rect 15112 4741 15150 4755
rect 15078 4707 15083 4721
rect 15117 4707 15150 4741
rect 14743 4691 14759 4707
rect 15078 4691 15150 4707
rect 15198 4725 15232 4794
rect 15266 4823 15344 4838
rect 15542 4829 15608 4845
rect 15542 4823 15574 4829
rect 15300 4822 15344 4823
rect 15300 4789 15310 4822
rect 15266 4788 15310 4789
rect 15266 4772 15344 4788
rect 15382 4789 15406 4823
rect 15440 4789 15456 4823
rect 15576 4789 15608 4795
rect 15382 4725 15416 4789
rect 15574 4779 15608 4789
rect 15653 4829 15704 4845
rect 15653 4795 15670 4829
rect 15653 4779 15704 4795
rect 15198 4691 15416 4725
rect 15484 4721 15530 4755
rect 15450 4718 15530 4721
rect 15653 4719 15687 4779
rect 15738 4747 15773 4878
rect 14709 4688 14759 4691
rect 14457 4623 14590 4657
rect 14709 4654 14716 4688
rect 14750 4654 14759 4688
rect 15450 4684 15496 4718
rect 15450 4668 15530 4684
rect 14709 4653 14759 4654
rect 14342 4585 14388 4619
rect 14556 4619 14590 4623
rect 14840 4623 15042 4657
rect 14556 4601 14773 4619
rect 14342 4551 14422 4585
rect 14456 4555 14472 4589
rect 14506 4555 14522 4589
rect 12316 4489 12345 4523
rect 12379 4489 12437 4523
rect 12471 4489 12529 4523
rect 12563 4489 12621 4523
rect 12655 4489 12713 4523
rect 12747 4489 12805 4523
rect 12839 4489 12897 4523
rect 12931 4489 12989 4523
rect 13023 4489 13081 4523
rect 13115 4489 13173 4523
rect 13207 4489 13265 4523
rect 13299 4489 13357 4523
rect 13391 4489 13449 4523
rect 13483 4489 13541 4523
rect 13575 4489 13633 4523
rect 13667 4489 13725 4523
rect 13759 4489 13788 4523
rect 14456 4517 14522 4555
rect 14556 4567 14739 4601
rect 14556 4551 14773 4567
rect 14840 4606 14874 4623
rect 15008 4606 15042 4623
rect 14840 4551 14874 4572
rect 14908 4555 14924 4589
rect 14958 4555 14974 4589
rect 14908 4517 14974 4555
rect 15183 4623 15398 4657
rect 15569 4655 15687 4719
rect 15721 4706 15773 4747
rect 15755 4682 15773 4706
rect 15569 4631 15603 4655
rect 15183 4606 15230 4623
rect 15008 4551 15042 4572
rect 15076 4559 15092 4593
rect 15126 4559 15142 4593
rect 15076 4517 15142 4559
rect 15183 4572 15196 4606
rect 15364 4606 15398 4623
rect 15183 4551 15230 4572
rect 15264 4555 15280 4589
rect 15314 4555 15330 4589
rect 15264 4517 15330 4555
rect 15364 4551 15398 4572
rect 15448 4606 15603 4631
rect 15721 4646 15732 4672
rect 15766 4646 15773 4682
rect 15482 4572 15603 4606
rect 15448 4551 15603 4572
rect 15637 4597 15687 4614
rect 15671 4563 15687 4597
rect 15637 4517 15687 4563
rect 15721 4612 15773 4646
rect 15755 4578 15773 4612
rect 15721 4551 15773 4578
rect 16364 4931 16444 4975
rect 16493 4971 16559 5009
rect 16493 4937 16509 4971
rect 16543 4937 16559 4971
rect 16593 4959 16795 4975
rect 16364 4897 16410 4931
rect 16593 4925 16761 4959
rect 16593 4903 16627 4925
rect 16761 4907 16795 4925
rect 16862 4954 16896 4975
rect 16930 4971 16996 5009
rect 16930 4937 16946 4971
rect 16980 4937 16996 4971
rect 17030 4954 17064 4975
rect 16364 4864 16444 4897
rect 16479 4869 16627 4903
rect 16862 4903 16896 4920
rect 17098 4962 17164 5009
rect 17098 4928 17114 4962
rect 17148 4928 17164 4962
rect 17218 4954 17252 4975
rect 17030 4903 17064 4920
rect 16364 4729 16430 4864
rect 16479 4827 16513 4869
rect 16464 4811 16513 4827
rect 16720 4839 16732 4873
rect 16766 4839 16819 4873
rect 16862 4869 17064 4903
rect 17286 4971 17352 5009
rect 17286 4937 17302 4971
rect 17336 4937 17352 4971
rect 17386 4954 17420 4975
rect 17218 4903 17252 4920
rect 17386 4903 17420 4920
rect 17218 4869 17420 4903
rect 17470 4954 17590 4975
rect 17504 4920 17590 4954
rect 17643 4967 17709 5009
rect 17643 4933 17659 4967
rect 17693 4933 17709 4967
rect 17470 4899 17590 4920
rect 17743 4931 17795 4975
rect 17470 4873 17709 4899
rect 17470 4839 17472 4873
rect 17506 4865 17709 4873
rect 17506 4839 17518 4865
rect 16720 4835 16819 4839
rect 16498 4777 16513 4811
rect 16464 4761 16513 4777
rect 16547 4805 16563 4819
rect 16547 4771 16548 4805
rect 16597 4785 16635 4819
rect 16720 4801 16803 4835
rect 16837 4801 16853 4835
rect 16887 4801 16903 4835
rect 16937 4805 16962 4835
rect 16582 4771 16635 4785
rect 16887 4771 16916 4801
rect 16950 4771 16962 4805
rect 17021 4776 17254 4833
rect 17675 4827 17709 4865
rect 17777 4897 17795 4931
rect 17743 4860 17795 4897
rect 16364 4691 16444 4729
rect 16364 4657 16410 4691
rect 16364 4601 16444 4657
rect 16479 4639 16513 4761
rect 16601 4707 16640 4737
rect 16601 4673 16635 4707
rect 16674 4703 16685 4737
rect 17021 4723 17055 4776
rect 16669 4673 16685 4703
rect 16731 4707 16988 4723
rect 16765 4689 16988 4707
rect 17022 4689 17055 4723
rect 17100 4737 17172 4739
rect 17134 4723 17172 4737
rect 17100 4689 17105 4703
rect 17139 4689 17172 4723
rect 16765 4673 16781 4689
rect 17100 4673 17172 4689
rect 17220 4707 17254 4776
rect 17288 4805 17366 4820
rect 17564 4811 17630 4827
rect 17564 4805 17596 4811
rect 17322 4804 17366 4805
rect 17322 4771 17332 4804
rect 17288 4770 17332 4771
rect 17288 4754 17366 4770
rect 17404 4771 17428 4805
rect 17462 4771 17478 4805
rect 17598 4771 17630 4777
rect 17404 4707 17438 4771
rect 17596 4761 17630 4771
rect 17675 4811 17726 4827
rect 17675 4777 17692 4811
rect 17675 4761 17726 4777
rect 17220 4673 17438 4707
rect 17506 4703 17552 4737
rect 17472 4700 17552 4703
rect 17675 4701 17709 4761
rect 17760 4729 17795 4860
rect 16731 4670 16781 4673
rect 16479 4605 16612 4639
rect 16731 4636 16738 4670
rect 16772 4636 16781 4670
rect 17472 4666 17518 4700
rect 17472 4650 17552 4666
rect 16731 4635 16781 4636
rect 16364 4567 16410 4601
rect 16578 4601 16612 4605
rect 16862 4605 17064 4639
rect 16578 4583 16795 4601
rect 16364 4533 16444 4567
rect 16478 4537 16494 4571
rect 16528 4537 16544 4571
rect 14318 4483 14347 4517
rect 14381 4483 14439 4517
rect 14473 4483 14531 4517
rect 14565 4483 14623 4517
rect 14657 4483 14715 4517
rect 14749 4483 14807 4517
rect 14841 4483 14899 4517
rect 14933 4483 14991 4517
rect 15025 4483 15083 4517
rect 15117 4483 15175 4517
rect 15209 4483 15267 4517
rect 15301 4483 15359 4517
rect 15393 4483 15451 4517
rect 15485 4483 15543 4517
rect 15577 4483 15635 4517
rect 15669 4483 15727 4517
rect 15761 4483 15790 4517
rect 16478 4499 16544 4537
rect 16578 4549 16761 4583
rect 16578 4533 16795 4549
rect 16862 4588 16896 4605
rect 17030 4588 17064 4605
rect 16862 4533 16896 4554
rect 16930 4537 16946 4571
rect 16980 4537 16996 4571
rect 16930 4499 16996 4537
rect 17205 4605 17420 4639
rect 17591 4637 17709 4701
rect 17743 4688 17795 4729
rect 17777 4664 17795 4688
rect 17591 4613 17625 4637
rect 17205 4588 17252 4605
rect 17030 4533 17064 4554
rect 17098 4541 17114 4575
rect 17148 4541 17164 4575
rect 17098 4499 17164 4541
rect 17205 4554 17218 4588
rect 17386 4588 17420 4605
rect 17205 4533 17252 4554
rect 17286 4537 17302 4571
rect 17336 4537 17352 4571
rect 17286 4499 17352 4537
rect 17386 4533 17420 4554
rect 17470 4588 17625 4613
rect 17743 4628 17754 4654
rect 17788 4628 17795 4664
rect 17504 4554 17625 4588
rect 17470 4533 17625 4554
rect 17659 4579 17709 4596
rect 17693 4545 17709 4579
rect 17659 4499 17709 4545
rect 17743 4594 17795 4628
rect 17777 4560 17795 4594
rect 17743 4533 17795 4560
rect 16340 4465 16369 4499
rect 16403 4465 16461 4499
rect 16495 4465 16553 4499
rect 16587 4465 16645 4499
rect 16679 4465 16737 4499
rect 16771 4465 16829 4499
rect 16863 4465 16921 4499
rect 16955 4465 17013 4499
rect 17047 4465 17105 4499
rect 17139 4465 17197 4499
rect 17231 4465 17289 4499
rect 17323 4465 17381 4499
rect 17415 4465 17473 4499
rect 17507 4465 17565 4499
rect 17599 4465 17657 4499
rect 17691 4465 17749 4499
rect 17783 4465 17812 4499
rect 1806 2271 1835 2305
rect 1869 2271 1927 2305
rect 1961 2271 2019 2305
rect 2053 2271 2111 2305
rect 2145 2271 2203 2305
rect 2237 2271 2295 2305
rect 2329 2271 2387 2305
rect 2421 2271 2479 2305
rect 2513 2271 2571 2305
rect 2605 2271 2663 2305
rect 2697 2271 2755 2305
rect 2789 2271 2847 2305
rect 2881 2271 2939 2305
rect 2973 2271 3031 2305
rect 3065 2271 3123 2305
rect 3157 2271 3215 2305
rect 3249 2271 3278 2305
rect 1830 2193 1910 2237
rect 1959 2233 2025 2271
rect 1959 2199 1975 2233
rect 2009 2199 2025 2233
rect 2059 2221 2261 2237
rect 1830 2159 1876 2193
rect 2059 2187 2227 2221
rect 2059 2165 2093 2187
rect 2227 2169 2261 2187
rect 2328 2216 2362 2237
rect 2396 2233 2462 2271
rect 2396 2199 2412 2233
rect 2446 2199 2462 2233
rect 2496 2216 2530 2237
rect 1830 2126 1910 2159
rect 1945 2131 2093 2165
rect 2328 2165 2362 2182
rect 2564 2224 2630 2271
rect 2564 2190 2580 2224
rect 2614 2190 2630 2224
rect 2684 2216 2718 2237
rect 2496 2165 2530 2182
rect 1830 1991 1896 2126
rect 1945 2089 1979 2131
rect 1930 2073 1979 2089
rect 2186 2101 2198 2135
rect 2232 2101 2285 2135
rect 2328 2131 2530 2165
rect 2752 2233 2818 2271
rect 2752 2199 2768 2233
rect 2802 2199 2818 2233
rect 2852 2216 2886 2237
rect 2684 2165 2718 2182
rect 2852 2165 2886 2182
rect 2684 2131 2886 2165
rect 2936 2216 3056 2237
rect 2970 2182 3056 2216
rect 3109 2229 3175 2271
rect 3876 2267 3905 2301
rect 3939 2267 3997 2301
rect 4031 2267 4089 2301
rect 4123 2267 4181 2301
rect 4215 2267 4273 2301
rect 4307 2267 4365 2301
rect 4399 2267 4457 2301
rect 4491 2267 4549 2301
rect 4583 2267 4641 2301
rect 4675 2267 4733 2301
rect 4767 2267 4825 2301
rect 4859 2267 4917 2301
rect 4951 2267 5009 2301
rect 5043 2267 5101 2301
rect 5135 2267 5193 2301
rect 5227 2267 5285 2301
rect 5319 2267 5348 2301
rect 5828 2267 5857 2301
rect 5891 2267 5949 2301
rect 5983 2267 6041 2301
rect 6075 2267 6133 2301
rect 6167 2267 6225 2301
rect 6259 2267 6317 2301
rect 6351 2267 6409 2301
rect 6443 2267 6501 2301
rect 6535 2267 6593 2301
rect 6627 2267 6685 2301
rect 6719 2267 6777 2301
rect 6811 2267 6869 2301
rect 6903 2267 6961 2301
rect 6995 2267 7053 2301
rect 7087 2267 7145 2301
rect 7179 2267 7237 2301
rect 7271 2267 7300 2301
rect 7830 2273 7859 2307
rect 7893 2273 7951 2307
rect 7985 2273 8043 2307
rect 8077 2273 8135 2307
rect 8169 2273 8227 2307
rect 8261 2273 8319 2307
rect 8353 2273 8411 2307
rect 8445 2273 8503 2307
rect 8537 2273 8595 2307
rect 8629 2273 8687 2307
rect 8721 2273 8779 2307
rect 8813 2273 8871 2307
rect 8905 2273 8963 2307
rect 8997 2273 9055 2307
rect 9089 2273 9147 2307
rect 9181 2273 9239 2307
rect 9273 2273 9302 2307
rect 9782 2273 9811 2307
rect 9845 2273 9903 2307
rect 9937 2273 9995 2307
rect 10029 2273 10087 2307
rect 10121 2273 10179 2307
rect 10213 2273 10271 2307
rect 10305 2273 10363 2307
rect 10397 2273 10455 2307
rect 10489 2273 10547 2307
rect 10581 2273 10639 2307
rect 10673 2273 10731 2307
rect 10765 2273 10823 2307
rect 10857 2273 10915 2307
rect 10949 2273 11007 2307
rect 11041 2273 11099 2307
rect 11133 2273 11191 2307
rect 11225 2273 11254 2307
rect 11774 2273 11803 2307
rect 11837 2273 11895 2307
rect 11929 2273 11987 2307
rect 12021 2273 12079 2307
rect 12113 2273 12171 2307
rect 12205 2273 12263 2307
rect 12297 2273 12355 2307
rect 12389 2273 12447 2307
rect 12481 2273 12539 2307
rect 12573 2273 12631 2307
rect 12665 2273 12723 2307
rect 12757 2273 12815 2307
rect 12849 2273 12907 2307
rect 12941 2273 12999 2307
rect 13033 2273 13091 2307
rect 13125 2273 13183 2307
rect 13217 2273 13246 2307
rect 13726 2273 13755 2307
rect 13789 2273 13847 2307
rect 13881 2273 13939 2307
rect 13973 2273 14031 2307
rect 14065 2273 14123 2307
rect 14157 2273 14215 2307
rect 14249 2273 14307 2307
rect 14341 2273 14399 2307
rect 14433 2273 14491 2307
rect 14525 2273 14583 2307
rect 14617 2273 14675 2307
rect 14709 2273 14767 2307
rect 14801 2273 14859 2307
rect 14893 2273 14951 2307
rect 14985 2273 15043 2307
rect 15077 2273 15135 2307
rect 15169 2273 15198 2307
rect 15790 2273 15819 2307
rect 15853 2273 15911 2307
rect 15945 2273 16003 2307
rect 16037 2273 16095 2307
rect 16129 2273 16187 2307
rect 16221 2273 16279 2307
rect 16313 2273 16371 2307
rect 16405 2273 16463 2307
rect 16497 2273 16555 2307
rect 16589 2273 16647 2307
rect 16681 2273 16739 2307
rect 16773 2273 16831 2307
rect 16865 2273 16923 2307
rect 16957 2273 17015 2307
rect 17049 2273 17107 2307
rect 17141 2273 17199 2307
rect 17233 2273 17262 2307
rect 3109 2195 3125 2229
rect 3159 2195 3175 2229
rect 2936 2161 3056 2182
rect 3209 2193 3261 2237
rect 2936 2135 3175 2161
rect 2936 2101 2938 2135
rect 2972 2127 3175 2135
rect 2972 2101 2984 2127
rect 2186 2097 2285 2101
rect 1964 2039 1979 2073
rect 1930 2023 1979 2039
rect 2013 2067 2029 2081
rect 2013 2033 2014 2067
rect 2063 2047 2101 2081
rect 2186 2063 2269 2097
rect 2303 2063 2319 2097
rect 2353 2063 2369 2097
rect 2403 2067 2428 2097
rect 2048 2033 2101 2047
rect 2353 2033 2382 2063
rect 2416 2033 2428 2067
rect 2487 2038 2720 2095
rect 3141 2089 3175 2127
rect 3243 2159 3261 2193
rect 3209 2122 3261 2159
rect 1830 1953 1910 1991
rect 1830 1919 1876 1953
rect 1830 1863 1910 1919
rect 1945 1901 1979 2023
rect 2067 1969 2106 1999
rect 2067 1935 2101 1969
rect 2140 1965 2151 1999
rect 2487 1985 2521 2038
rect 2135 1935 2151 1965
rect 2197 1969 2454 1985
rect 2231 1951 2454 1969
rect 2488 1951 2521 1985
rect 2566 1999 2638 2001
rect 2600 1985 2638 1999
rect 2566 1951 2571 1965
rect 2605 1951 2638 1985
rect 2231 1935 2247 1951
rect 2566 1935 2638 1951
rect 2686 1969 2720 2038
rect 2754 2067 2832 2082
rect 3030 2073 3096 2089
rect 3030 2067 3062 2073
rect 2788 2066 2832 2067
rect 2788 2033 2798 2066
rect 2754 2032 2798 2033
rect 2754 2016 2832 2032
rect 2870 2033 2894 2067
rect 2928 2033 2944 2067
rect 3064 2033 3096 2039
rect 2870 1969 2904 2033
rect 3062 2023 3096 2033
rect 3141 2073 3192 2089
rect 3141 2039 3158 2073
rect 3141 2023 3192 2039
rect 2686 1935 2904 1969
rect 2972 1965 3018 1999
rect 2938 1962 3018 1965
rect 3141 1963 3175 2023
rect 3226 1991 3261 2122
rect 2197 1934 2247 1935
rect 1945 1867 2078 1901
rect 2197 1900 2206 1934
rect 2240 1900 2247 1934
rect 2938 1928 2984 1962
rect 2938 1912 3018 1928
rect 2197 1897 2247 1900
rect 1830 1829 1876 1863
rect 2044 1863 2078 1867
rect 2328 1867 2530 1901
rect 2044 1845 2261 1863
rect 1830 1795 1910 1829
rect 1944 1799 1960 1833
rect 1994 1799 2010 1833
rect 1944 1761 2010 1799
rect 2044 1811 2227 1845
rect 2044 1795 2261 1811
rect 2328 1850 2362 1867
rect 2496 1850 2530 1867
rect 2328 1795 2362 1816
rect 2396 1799 2412 1833
rect 2446 1799 2462 1833
rect 2396 1761 2462 1799
rect 2671 1867 2886 1901
rect 3057 1899 3175 1963
rect 3209 1950 3261 1991
rect 3243 1926 3261 1950
rect 3057 1875 3091 1899
rect 2671 1850 2718 1867
rect 2496 1795 2530 1816
rect 2564 1803 2580 1837
rect 2614 1803 2630 1837
rect 2564 1761 2630 1803
rect 2671 1816 2684 1850
rect 2852 1850 2886 1867
rect 2671 1795 2718 1816
rect 2752 1799 2768 1833
rect 2802 1799 2818 1833
rect 2752 1761 2818 1799
rect 2852 1795 2886 1816
rect 2936 1850 3091 1875
rect 3209 1890 3214 1916
rect 3254 1890 3261 1926
rect 2970 1816 3091 1850
rect 2936 1795 3091 1816
rect 3125 1841 3175 1858
rect 3159 1807 3175 1841
rect 3125 1761 3175 1807
rect 3209 1856 3261 1890
rect 3243 1822 3261 1856
rect 3209 1795 3261 1822
rect 3900 2189 3980 2233
rect 4029 2229 4095 2267
rect 4029 2195 4045 2229
rect 4079 2195 4095 2229
rect 4129 2217 4331 2233
rect 3900 2155 3946 2189
rect 4129 2183 4297 2217
rect 4129 2161 4163 2183
rect 4297 2165 4331 2183
rect 4398 2212 4432 2233
rect 4466 2229 4532 2267
rect 4466 2195 4482 2229
rect 4516 2195 4532 2229
rect 4566 2212 4600 2233
rect 3900 2122 3980 2155
rect 4015 2127 4163 2161
rect 4398 2161 4432 2178
rect 4634 2220 4700 2267
rect 4634 2186 4650 2220
rect 4684 2186 4700 2220
rect 4754 2212 4788 2233
rect 4566 2161 4600 2178
rect 3900 1987 3966 2122
rect 4015 2085 4049 2127
rect 4000 2069 4049 2085
rect 4256 2097 4268 2131
rect 4302 2097 4355 2131
rect 4398 2127 4600 2161
rect 4822 2229 4888 2267
rect 4822 2195 4838 2229
rect 4872 2195 4888 2229
rect 4922 2212 4956 2233
rect 4754 2161 4788 2178
rect 4922 2161 4956 2178
rect 4754 2127 4956 2161
rect 5006 2212 5126 2233
rect 5040 2178 5126 2212
rect 5179 2225 5245 2267
rect 5179 2191 5195 2225
rect 5229 2191 5245 2225
rect 5006 2157 5126 2178
rect 5279 2189 5331 2233
rect 5006 2131 5245 2157
rect 5006 2097 5008 2131
rect 5042 2123 5245 2131
rect 5042 2097 5054 2123
rect 4256 2093 4355 2097
rect 4034 2035 4049 2069
rect 4000 2019 4049 2035
rect 4083 2063 4099 2077
rect 4083 2029 4084 2063
rect 4133 2043 4171 2077
rect 4256 2059 4339 2093
rect 4373 2059 4389 2093
rect 4423 2059 4439 2093
rect 4473 2063 4498 2093
rect 4118 2029 4171 2043
rect 4423 2029 4452 2059
rect 4486 2029 4498 2063
rect 4557 2034 4790 2091
rect 5211 2085 5245 2123
rect 5313 2155 5331 2189
rect 5279 2118 5331 2155
rect 3900 1949 3980 1987
rect 3900 1915 3946 1949
rect 3900 1859 3980 1915
rect 4015 1897 4049 2019
rect 4137 1965 4176 1995
rect 4137 1931 4171 1965
rect 4210 1961 4221 1995
rect 4557 1981 4591 2034
rect 4205 1931 4221 1961
rect 4267 1965 4524 1981
rect 4301 1947 4524 1965
rect 4558 1947 4591 1981
rect 4636 1995 4708 1997
rect 4670 1981 4708 1995
rect 4636 1947 4641 1961
rect 4675 1947 4708 1981
rect 4301 1931 4317 1947
rect 4636 1931 4708 1947
rect 4756 1965 4790 2034
rect 4824 2063 4902 2078
rect 5100 2069 5166 2085
rect 5100 2063 5132 2069
rect 4858 2062 4902 2063
rect 4858 2029 4868 2062
rect 4824 2028 4868 2029
rect 4824 2012 4902 2028
rect 4940 2029 4964 2063
rect 4998 2029 5014 2063
rect 5134 2029 5166 2035
rect 4940 1965 4974 2029
rect 5132 2019 5166 2029
rect 5211 2069 5262 2085
rect 5211 2035 5228 2069
rect 5211 2019 5262 2035
rect 4756 1931 4974 1965
rect 5042 1961 5088 1995
rect 5008 1958 5088 1961
rect 5211 1959 5245 2019
rect 5296 1987 5331 2118
rect 4267 1928 4317 1931
rect 4015 1863 4148 1897
rect 4267 1894 4274 1928
rect 4308 1894 4317 1928
rect 5008 1924 5054 1958
rect 5008 1908 5088 1924
rect 4267 1893 4317 1894
rect 3900 1825 3946 1859
rect 4114 1859 4148 1863
rect 4398 1863 4600 1897
rect 4114 1841 4331 1859
rect 3900 1791 3980 1825
rect 4014 1795 4030 1829
rect 4064 1795 4080 1829
rect 1806 1727 1835 1761
rect 1869 1727 1927 1761
rect 1961 1727 2019 1761
rect 2053 1727 2111 1761
rect 2145 1727 2203 1761
rect 2237 1727 2295 1761
rect 2329 1727 2387 1761
rect 2421 1727 2479 1761
rect 2513 1727 2571 1761
rect 2605 1727 2663 1761
rect 2697 1727 2755 1761
rect 2789 1727 2847 1761
rect 2881 1727 2939 1761
rect 2973 1727 3031 1761
rect 3065 1727 3123 1761
rect 3157 1727 3215 1761
rect 3249 1727 3278 1761
rect 4014 1757 4080 1795
rect 4114 1807 4297 1841
rect 4114 1791 4331 1807
rect 4398 1846 4432 1863
rect 4566 1846 4600 1863
rect 4398 1791 4432 1812
rect 4466 1795 4482 1829
rect 4516 1795 4532 1829
rect 4466 1757 4532 1795
rect 4741 1863 4956 1897
rect 5127 1895 5245 1959
rect 5279 1946 5331 1987
rect 5313 1922 5331 1946
rect 5127 1871 5161 1895
rect 4741 1846 4788 1863
rect 4566 1791 4600 1812
rect 4634 1799 4650 1833
rect 4684 1799 4700 1833
rect 4634 1757 4700 1799
rect 4741 1812 4754 1846
rect 4922 1846 4956 1863
rect 4741 1791 4788 1812
rect 4822 1795 4838 1829
rect 4872 1795 4888 1829
rect 4822 1757 4888 1795
rect 4922 1791 4956 1812
rect 5006 1846 5161 1871
rect 5279 1886 5290 1912
rect 5324 1886 5331 1922
rect 5040 1812 5161 1846
rect 5006 1791 5161 1812
rect 5195 1837 5245 1854
rect 5229 1803 5245 1837
rect 5195 1757 5245 1803
rect 5279 1852 5331 1886
rect 5313 1818 5331 1852
rect 5279 1791 5331 1818
rect 5852 2189 5932 2233
rect 5981 2229 6047 2267
rect 5981 2195 5997 2229
rect 6031 2195 6047 2229
rect 6081 2217 6283 2233
rect 5852 2155 5898 2189
rect 6081 2183 6249 2217
rect 6081 2161 6115 2183
rect 6249 2165 6283 2183
rect 6350 2212 6384 2233
rect 6418 2229 6484 2267
rect 6418 2195 6434 2229
rect 6468 2195 6484 2229
rect 6518 2212 6552 2233
rect 5852 2122 5932 2155
rect 5967 2127 6115 2161
rect 6350 2161 6384 2178
rect 6586 2220 6652 2267
rect 6586 2186 6602 2220
rect 6636 2186 6652 2220
rect 6706 2212 6740 2233
rect 6518 2161 6552 2178
rect 5852 1987 5918 2122
rect 5967 2085 6001 2127
rect 5952 2069 6001 2085
rect 6208 2097 6220 2131
rect 6254 2097 6307 2131
rect 6350 2127 6552 2161
rect 6774 2229 6840 2267
rect 6774 2195 6790 2229
rect 6824 2195 6840 2229
rect 6874 2212 6908 2233
rect 6706 2161 6740 2178
rect 6874 2161 6908 2178
rect 6706 2127 6908 2161
rect 6958 2212 7078 2233
rect 6992 2178 7078 2212
rect 7131 2225 7197 2267
rect 7131 2191 7147 2225
rect 7181 2191 7197 2225
rect 6958 2157 7078 2178
rect 7231 2189 7283 2233
rect 6958 2131 7197 2157
rect 6958 2097 6960 2131
rect 6994 2123 7197 2131
rect 6994 2097 7006 2123
rect 6208 2093 6307 2097
rect 5986 2035 6001 2069
rect 5952 2019 6001 2035
rect 6035 2063 6051 2077
rect 6035 2029 6036 2063
rect 6085 2043 6123 2077
rect 6208 2059 6291 2093
rect 6325 2059 6341 2093
rect 6375 2059 6391 2093
rect 6425 2063 6450 2093
rect 6070 2029 6123 2043
rect 6375 2029 6404 2059
rect 6438 2029 6450 2063
rect 6509 2034 6742 2091
rect 7163 2085 7197 2123
rect 7265 2155 7283 2189
rect 7231 2118 7283 2155
rect 5852 1949 5932 1987
rect 5852 1915 5898 1949
rect 5852 1859 5932 1915
rect 5967 1897 6001 2019
rect 6089 1965 6128 1995
rect 6089 1931 6123 1965
rect 6162 1961 6173 1995
rect 6509 1981 6543 2034
rect 6157 1931 6173 1961
rect 6219 1965 6476 1981
rect 6253 1947 6476 1965
rect 6510 1947 6543 1981
rect 6588 1995 6660 1997
rect 6622 1981 6660 1995
rect 6588 1947 6593 1961
rect 6627 1947 6660 1981
rect 6253 1931 6269 1947
rect 6588 1931 6660 1947
rect 6708 1965 6742 2034
rect 6776 2063 6854 2078
rect 7052 2069 7118 2085
rect 7052 2063 7084 2069
rect 6810 2062 6854 2063
rect 6810 2029 6820 2062
rect 6776 2028 6820 2029
rect 6776 2012 6854 2028
rect 6892 2029 6916 2063
rect 6950 2029 6966 2063
rect 7086 2029 7118 2035
rect 6892 1965 6926 2029
rect 7084 2019 7118 2029
rect 7163 2069 7214 2085
rect 7163 2035 7180 2069
rect 7163 2019 7214 2035
rect 6708 1931 6926 1965
rect 6994 1961 7040 1995
rect 6960 1958 7040 1961
rect 7163 1959 7197 2019
rect 7248 1987 7283 2118
rect 6219 1928 6269 1931
rect 5967 1863 6100 1897
rect 6219 1894 6226 1928
rect 6260 1894 6269 1928
rect 6960 1924 7006 1958
rect 6960 1908 7040 1924
rect 6219 1893 6269 1894
rect 5852 1825 5898 1859
rect 6066 1859 6100 1863
rect 6350 1863 6552 1897
rect 6066 1841 6283 1859
rect 5852 1791 5932 1825
rect 5966 1795 5982 1829
rect 6016 1795 6032 1829
rect 5966 1757 6032 1795
rect 6066 1807 6249 1841
rect 6066 1791 6283 1807
rect 6350 1846 6384 1863
rect 6518 1846 6552 1863
rect 6350 1791 6384 1812
rect 6418 1795 6434 1829
rect 6468 1795 6484 1829
rect 6418 1757 6484 1795
rect 6693 1863 6908 1897
rect 7079 1895 7197 1959
rect 7231 1946 7283 1987
rect 7265 1922 7283 1946
rect 7079 1871 7113 1895
rect 6693 1846 6740 1863
rect 6518 1791 6552 1812
rect 6586 1799 6602 1833
rect 6636 1799 6652 1833
rect 6586 1757 6652 1799
rect 6693 1812 6706 1846
rect 6874 1846 6908 1863
rect 6693 1791 6740 1812
rect 6774 1795 6790 1829
rect 6824 1795 6840 1829
rect 6774 1757 6840 1795
rect 6874 1791 6908 1812
rect 6958 1846 7113 1871
rect 7231 1886 7242 1912
rect 7276 1886 7283 1922
rect 6992 1812 7113 1846
rect 6958 1791 7113 1812
rect 7147 1837 7197 1854
rect 7181 1803 7197 1837
rect 7147 1757 7197 1803
rect 7231 1852 7283 1886
rect 7265 1818 7283 1852
rect 7231 1791 7283 1818
rect 7854 2195 7934 2239
rect 7983 2235 8049 2273
rect 7983 2201 7999 2235
rect 8033 2201 8049 2235
rect 8083 2223 8285 2239
rect 7854 2161 7900 2195
rect 8083 2189 8251 2223
rect 8083 2167 8117 2189
rect 8251 2171 8285 2189
rect 8352 2218 8386 2239
rect 8420 2235 8486 2273
rect 8420 2201 8436 2235
rect 8470 2201 8486 2235
rect 8520 2218 8554 2239
rect 7854 2128 7934 2161
rect 7969 2133 8117 2167
rect 8352 2167 8386 2184
rect 8588 2226 8654 2273
rect 8588 2192 8604 2226
rect 8638 2192 8654 2226
rect 8708 2218 8742 2239
rect 8520 2167 8554 2184
rect 7854 1993 7920 2128
rect 7969 2091 8003 2133
rect 7954 2075 8003 2091
rect 8210 2103 8222 2137
rect 8256 2103 8309 2137
rect 8352 2133 8554 2167
rect 8776 2235 8842 2273
rect 8776 2201 8792 2235
rect 8826 2201 8842 2235
rect 8876 2218 8910 2239
rect 8708 2167 8742 2184
rect 8876 2167 8910 2184
rect 8708 2133 8910 2167
rect 8960 2218 9080 2239
rect 8994 2184 9080 2218
rect 9133 2231 9199 2273
rect 9133 2197 9149 2231
rect 9183 2197 9199 2231
rect 8960 2163 9080 2184
rect 9233 2195 9285 2239
rect 8960 2137 9199 2163
rect 8960 2103 8962 2137
rect 8996 2129 9199 2137
rect 8996 2103 9008 2129
rect 8210 2099 8309 2103
rect 7988 2041 8003 2075
rect 7954 2025 8003 2041
rect 8037 2069 8053 2083
rect 8037 2035 8038 2069
rect 8087 2049 8125 2083
rect 8210 2065 8293 2099
rect 8327 2065 8343 2099
rect 8377 2065 8393 2099
rect 8427 2069 8452 2099
rect 8072 2035 8125 2049
rect 8377 2035 8406 2065
rect 8440 2035 8452 2069
rect 8511 2040 8744 2097
rect 9165 2091 9199 2129
rect 9267 2161 9285 2195
rect 9233 2124 9285 2161
rect 7854 1955 7934 1993
rect 7854 1921 7900 1955
rect 7854 1865 7934 1921
rect 7969 1903 8003 2025
rect 8091 1971 8130 2001
rect 8091 1937 8125 1971
rect 8164 1967 8175 2001
rect 8511 1987 8545 2040
rect 8159 1937 8175 1967
rect 8221 1971 8478 1987
rect 8255 1953 8478 1971
rect 8512 1953 8545 1987
rect 8590 2001 8662 2003
rect 8624 1987 8662 2001
rect 8590 1953 8595 1967
rect 8629 1953 8662 1987
rect 8255 1937 8271 1953
rect 8590 1937 8662 1953
rect 8710 1971 8744 2040
rect 8778 2069 8856 2084
rect 9054 2075 9120 2091
rect 9054 2069 9086 2075
rect 8812 2068 8856 2069
rect 8812 2035 8822 2068
rect 8778 2034 8822 2035
rect 8778 2018 8856 2034
rect 8894 2035 8918 2069
rect 8952 2035 8968 2069
rect 9088 2035 9120 2041
rect 8894 1971 8928 2035
rect 9086 2025 9120 2035
rect 9165 2075 9216 2091
rect 9165 2041 9182 2075
rect 9165 2025 9216 2041
rect 8710 1937 8928 1971
rect 8996 1967 9042 2001
rect 8962 1964 9042 1967
rect 9165 1965 9199 2025
rect 9250 1993 9285 2124
rect 8221 1934 8271 1937
rect 7969 1869 8102 1903
rect 8221 1900 8228 1934
rect 8262 1900 8271 1934
rect 8962 1930 9008 1964
rect 8962 1914 9042 1930
rect 8221 1899 8271 1900
rect 7854 1831 7900 1865
rect 8068 1865 8102 1869
rect 8352 1869 8554 1903
rect 8068 1847 8285 1865
rect 7854 1797 7934 1831
rect 7968 1801 7984 1835
rect 8018 1801 8034 1835
rect 7968 1763 8034 1801
rect 8068 1813 8251 1847
rect 8068 1797 8285 1813
rect 8352 1852 8386 1869
rect 8520 1852 8554 1869
rect 8352 1797 8386 1818
rect 8420 1801 8436 1835
rect 8470 1801 8486 1835
rect 8420 1763 8486 1801
rect 8695 1869 8910 1903
rect 9081 1901 9199 1965
rect 9233 1952 9285 1993
rect 9267 1928 9285 1952
rect 9081 1877 9115 1901
rect 8695 1852 8742 1869
rect 8520 1797 8554 1818
rect 8588 1805 8604 1839
rect 8638 1805 8654 1839
rect 8588 1763 8654 1805
rect 8695 1818 8708 1852
rect 8876 1852 8910 1869
rect 8695 1797 8742 1818
rect 8776 1801 8792 1835
rect 8826 1801 8842 1835
rect 8776 1763 8842 1801
rect 8876 1797 8910 1818
rect 8960 1852 9115 1877
rect 9233 1892 9244 1918
rect 9278 1892 9285 1928
rect 8994 1818 9115 1852
rect 8960 1797 9115 1818
rect 9149 1843 9199 1860
rect 9183 1809 9199 1843
rect 9149 1763 9199 1809
rect 9233 1858 9285 1892
rect 9267 1824 9285 1858
rect 9233 1797 9285 1824
rect 9806 2195 9886 2239
rect 9935 2235 10001 2273
rect 9935 2201 9951 2235
rect 9985 2201 10001 2235
rect 10035 2223 10237 2239
rect 9806 2161 9852 2195
rect 10035 2189 10203 2223
rect 10035 2167 10069 2189
rect 10203 2171 10237 2189
rect 10304 2218 10338 2239
rect 10372 2235 10438 2273
rect 10372 2201 10388 2235
rect 10422 2201 10438 2235
rect 10472 2218 10506 2239
rect 9806 2128 9886 2161
rect 9921 2133 10069 2167
rect 10304 2167 10338 2184
rect 10540 2226 10606 2273
rect 10540 2192 10556 2226
rect 10590 2192 10606 2226
rect 10660 2218 10694 2239
rect 10472 2167 10506 2184
rect 9806 1993 9872 2128
rect 9921 2091 9955 2133
rect 9906 2075 9955 2091
rect 10162 2103 10174 2137
rect 10208 2103 10261 2137
rect 10304 2133 10506 2167
rect 10728 2235 10794 2273
rect 10728 2201 10744 2235
rect 10778 2201 10794 2235
rect 10828 2218 10862 2239
rect 10660 2167 10694 2184
rect 10828 2167 10862 2184
rect 10660 2133 10862 2167
rect 10912 2218 11032 2239
rect 10946 2184 11032 2218
rect 11085 2231 11151 2273
rect 11085 2197 11101 2231
rect 11135 2197 11151 2231
rect 10912 2163 11032 2184
rect 11185 2195 11237 2239
rect 10912 2137 11151 2163
rect 10912 2103 10914 2137
rect 10948 2129 11151 2137
rect 10948 2103 10960 2129
rect 10162 2099 10261 2103
rect 9940 2041 9955 2075
rect 9906 2025 9955 2041
rect 9989 2069 10005 2083
rect 9989 2035 9990 2069
rect 10039 2049 10077 2083
rect 10162 2065 10245 2099
rect 10279 2065 10295 2099
rect 10329 2065 10345 2099
rect 10379 2069 10404 2099
rect 10024 2035 10077 2049
rect 10329 2035 10358 2065
rect 10392 2035 10404 2069
rect 10463 2040 10696 2097
rect 11117 2091 11151 2129
rect 11219 2161 11237 2195
rect 11185 2124 11237 2161
rect 9806 1955 9886 1993
rect 9806 1921 9852 1955
rect 9806 1865 9886 1921
rect 9921 1903 9955 2025
rect 10043 1971 10082 2001
rect 10043 1937 10077 1971
rect 10116 1967 10127 2001
rect 10463 1987 10497 2040
rect 10111 1937 10127 1967
rect 10173 1971 10430 1987
rect 10207 1953 10430 1971
rect 10464 1953 10497 1987
rect 10542 2001 10614 2003
rect 10576 1987 10614 2001
rect 10542 1953 10547 1967
rect 10581 1953 10614 1987
rect 10207 1937 10223 1953
rect 10542 1937 10614 1953
rect 10662 1971 10696 2040
rect 10730 2069 10808 2084
rect 11006 2075 11072 2091
rect 11006 2069 11038 2075
rect 10764 2068 10808 2069
rect 10764 2035 10774 2068
rect 10730 2034 10774 2035
rect 10730 2018 10808 2034
rect 10846 2035 10870 2069
rect 10904 2035 10920 2069
rect 11040 2035 11072 2041
rect 10846 1971 10880 2035
rect 11038 2025 11072 2035
rect 11117 2075 11168 2091
rect 11117 2041 11134 2075
rect 11117 2025 11168 2041
rect 10662 1937 10880 1971
rect 10948 1967 10994 2001
rect 10914 1964 10994 1967
rect 11117 1965 11151 2025
rect 11202 1993 11237 2124
rect 10173 1934 10223 1937
rect 9921 1869 10054 1903
rect 10173 1900 10180 1934
rect 10214 1900 10223 1934
rect 10914 1930 10960 1964
rect 10914 1914 10994 1930
rect 10173 1899 10223 1900
rect 9806 1831 9852 1865
rect 10020 1865 10054 1869
rect 10304 1869 10506 1903
rect 10020 1847 10237 1865
rect 9806 1797 9886 1831
rect 9920 1801 9936 1835
rect 9970 1801 9986 1835
rect 9920 1763 9986 1801
rect 10020 1813 10203 1847
rect 10020 1797 10237 1813
rect 10304 1852 10338 1869
rect 10472 1852 10506 1869
rect 10304 1797 10338 1818
rect 10372 1801 10388 1835
rect 10422 1801 10438 1835
rect 10372 1763 10438 1801
rect 10647 1869 10862 1903
rect 11033 1901 11151 1965
rect 11185 1952 11237 1993
rect 11219 1928 11237 1952
rect 11033 1877 11067 1901
rect 10647 1852 10694 1869
rect 10472 1797 10506 1818
rect 10540 1805 10556 1839
rect 10590 1805 10606 1839
rect 10540 1763 10606 1805
rect 10647 1818 10660 1852
rect 10828 1852 10862 1869
rect 10647 1797 10694 1818
rect 10728 1801 10744 1835
rect 10778 1801 10794 1835
rect 10728 1763 10794 1801
rect 10828 1797 10862 1818
rect 10912 1852 11067 1877
rect 11185 1892 11196 1918
rect 11230 1892 11237 1928
rect 10946 1818 11067 1852
rect 10912 1797 11067 1818
rect 11101 1843 11151 1860
rect 11135 1809 11151 1843
rect 11101 1763 11151 1809
rect 11185 1858 11237 1892
rect 11219 1824 11237 1858
rect 11185 1797 11237 1824
rect 11798 2195 11878 2239
rect 11927 2235 11993 2273
rect 11927 2201 11943 2235
rect 11977 2201 11993 2235
rect 12027 2223 12229 2239
rect 11798 2161 11844 2195
rect 12027 2189 12195 2223
rect 12027 2167 12061 2189
rect 12195 2171 12229 2189
rect 12296 2218 12330 2239
rect 12364 2235 12430 2273
rect 12364 2201 12380 2235
rect 12414 2201 12430 2235
rect 12464 2218 12498 2239
rect 11798 2128 11878 2161
rect 11913 2133 12061 2167
rect 12296 2167 12330 2184
rect 12532 2226 12598 2273
rect 12532 2192 12548 2226
rect 12582 2192 12598 2226
rect 12652 2218 12686 2239
rect 12464 2167 12498 2184
rect 11798 1993 11864 2128
rect 11913 2091 11947 2133
rect 11898 2075 11947 2091
rect 12154 2103 12166 2137
rect 12200 2103 12253 2137
rect 12296 2133 12498 2167
rect 12720 2235 12786 2273
rect 12720 2201 12736 2235
rect 12770 2201 12786 2235
rect 12820 2218 12854 2239
rect 12652 2167 12686 2184
rect 12820 2167 12854 2184
rect 12652 2133 12854 2167
rect 12904 2218 13024 2239
rect 12938 2184 13024 2218
rect 13077 2231 13143 2273
rect 13077 2197 13093 2231
rect 13127 2197 13143 2231
rect 12904 2163 13024 2184
rect 13177 2195 13229 2239
rect 12904 2137 13143 2163
rect 12904 2103 12906 2137
rect 12940 2129 13143 2137
rect 12940 2103 12952 2129
rect 12154 2099 12253 2103
rect 11932 2041 11947 2075
rect 11898 2025 11947 2041
rect 11981 2069 11997 2083
rect 11981 2035 11982 2069
rect 12031 2049 12069 2083
rect 12154 2065 12237 2099
rect 12271 2065 12287 2099
rect 12321 2065 12337 2099
rect 12371 2069 12396 2099
rect 12016 2035 12069 2049
rect 12321 2035 12350 2065
rect 12384 2035 12396 2069
rect 12455 2040 12688 2097
rect 13109 2091 13143 2129
rect 13211 2161 13229 2195
rect 13177 2124 13229 2161
rect 11798 1955 11878 1993
rect 11798 1921 11844 1955
rect 11798 1865 11878 1921
rect 11913 1903 11947 2025
rect 12035 1971 12074 2001
rect 12035 1937 12069 1971
rect 12108 1967 12119 2001
rect 12455 1987 12489 2040
rect 12103 1937 12119 1967
rect 12165 1971 12422 1987
rect 12199 1953 12422 1971
rect 12456 1953 12489 1987
rect 12534 2001 12606 2003
rect 12568 1987 12606 2001
rect 12534 1953 12539 1967
rect 12573 1953 12606 1987
rect 12199 1937 12215 1953
rect 12534 1937 12606 1953
rect 12654 1971 12688 2040
rect 12722 2069 12800 2084
rect 12998 2075 13064 2091
rect 12998 2069 13030 2075
rect 12756 2068 12800 2069
rect 12756 2035 12766 2068
rect 12722 2034 12766 2035
rect 12722 2018 12800 2034
rect 12838 2035 12862 2069
rect 12896 2035 12912 2069
rect 13032 2035 13064 2041
rect 12838 1971 12872 2035
rect 13030 2025 13064 2035
rect 13109 2075 13160 2091
rect 13109 2041 13126 2075
rect 13109 2025 13160 2041
rect 12654 1937 12872 1971
rect 12940 1967 12986 2001
rect 12906 1964 12986 1967
rect 13109 1965 13143 2025
rect 13194 1993 13229 2124
rect 12165 1934 12215 1937
rect 11913 1869 12046 1903
rect 12165 1900 12172 1934
rect 12206 1900 12215 1934
rect 12906 1930 12952 1964
rect 12906 1914 12986 1930
rect 12165 1899 12215 1900
rect 11798 1831 11844 1865
rect 12012 1865 12046 1869
rect 12296 1869 12498 1903
rect 12012 1847 12229 1865
rect 11798 1797 11878 1831
rect 11912 1801 11928 1835
rect 11962 1801 11978 1835
rect 11912 1763 11978 1801
rect 12012 1813 12195 1847
rect 12012 1797 12229 1813
rect 12296 1852 12330 1869
rect 12464 1852 12498 1869
rect 12296 1797 12330 1818
rect 12364 1801 12380 1835
rect 12414 1801 12430 1835
rect 12364 1763 12430 1801
rect 12639 1869 12854 1903
rect 13025 1901 13143 1965
rect 13177 1952 13229 1993
rect 13211 1928 13229 1952
rect 13025 1877 13059 1901
rect 12639 1852 12686 1869
rect 12464 1797 12498 1818
rect 12532 1805 12548 1839
rect 12582 1805 12598 1839
rect 12532 1763 12598 1805
rect 12639 1818 12652 1852
rect 12820 1852 12854 1869
rect 12639 1797 12686 1818
rect 12720 1801 12736 1835
rect 12770 1801 12786 1835
rect 12720 1763 12786 1801
rect 12820 1797 12854 1818
rect 12904 1852 13059 1877
rect 13177 1892 13188 1918
rect 13222 1892 13229 1928
rect 12938 1818 13059 1852
rect 12904 1797 13059 1818
rect 13093 1843 13143 1860
rect 13127 1809 13143 1843
rect 13093 1763 13143 1809
rect 13177 1858 13229 1892
rect 13211 1824 13229 1858
rect 13177 1797 13229 1824
rect 13750 2195 13830 2239
rect 13879 2235 13945 2273
rect 13879 2201 13895 2235
rect 13929 2201 13945 2235
rect 13979 2223 14181 2239
rect 13750 2161 13796 2195
rect 13979 2189 14147 2223
rect 13979 2167 14013 2189
rect 14147 2171 14181 2189
rect 14248 2218 14282 2239
rect 14316 2235 14382 2273
rect 14316 2201 14332 2235
rect 14366 2201 14382 2235
rect 14416 2218 14450 2239
rect 13750 2128 13830 2161
rect 13865 2133 14013 2167
rect 14248 2167 14282 2184
rect 14484 2226 14550 2273
rect 14484 2192 14500 2226
rect 14534 2192 14550 2226
rect 14604 2218 14638 2239
rect 14416 2167 14450 2184
rect 13750 1993 13816 2128
rect 13865 2091 13899 2133
rect 13850 2075 13899 2091
rect 14106 2103 14118 2137
rect 14152 2103 14205 2137
rect 14248 2133 14450 2167
rect 14672 2235 14738 2273
rect 14672 2201 14688 2235
rect 14722 2201 14738 2235
rect 14772 2218 14806 2239
rect 14604 2167 14638 2184
rect 14772 2167 14806 2184
rect 14604 2133 14806 2167
rect 14856 2218 14976 2239
rect 14890 2184 14976 2218
rect 15029 2231 15095 2273
rect 15029 2197 15045 2231
rect 15079 2197 15095 2231
rect 14856 2163 14976 2184
rect 15129 2195 15181 2239
rect 14856 2137 15095 2163
rect 14856 2103 14858 2137
rect 14892 2129 15095 2137
rect 14892 2103 14904 2129
rect 14106 2099 14205 2103
rect 13884 2041 13899 2075
rect 13850 2025 13899 2041
rect 13933 2069 13949 2083
rect 13933 2035 13934 2069
rect 13983 2049 14021 2083
rect 14106 2065 14189 2099
rect 14223 2065 14239 2099
rect 14273 2065 14289 2099
rect 14323 2069 14348 2099
rect 13968 2035 14021 2049
rect 14273 2035 14302 2065
rect 14336 2035 14348 2069
rect 14407 2040 14640 2097
rect 15061 2091 15095 2129
rect 15163 2161 15181 2195
rect 15129 2124 15181 2161
rect 13750 1955 13830 1993
rect 13750 1921 13796 1955
rect 13750 1865 13830 1921
rect 13865 1903 13899 2025
rect 13987 1971 14026 2001
rect 13987 1937 14021 1971
rect 14060 1967 14071 2001
rect 14407 1987 14441 2040
rect 14055 1937 14071 1967
rect 14117 1971 14374 1987
rect 14151 1953 14374 1971
rect 14408 1953 14441 1987
rect 14486 2001 14558 2003
rect 14520 1987 14558 2001
rect 14486 1953 14491 1967
rect 14525 1953 14558 1987
rect 14151 1937 14167 1953
rect 14486 1937 14558 1953
rect 14606 1971 14640 2040
rect 14674 2069 14752 2084
rect 14950 2075 15016 2091
rect 14950 2069 14982 2075
rect 14708 2068 14752 2069
rect 14708 2035 14718 2068
rect 14674 2034 14718 2035
rect 14674 2018 14752 2034
rect 14790 2035 14814 2069
rect 14848 2035 14864 2069
rect 14984 2035 15016 2041
rect 14790 1971 14824 2035
rect 14982 2025 15016 2035
rect 15061 2075 15112 2091
rect 15061 2041 15078 2075
rect 15061 2025 15112 2041
rect 14606 1937 14824 1971
rect 14892 1967 14938 2001
rect 14858 1964 14938 1967
rect 15061 1965 15095 2025
rect 15146 1993 15181 2124
rect 14117 1934 14167 1937
rect 13865 1869 13998 1903
rect 14117 1900 14124 1934
rect 14158 1900 14167 1934
rect 14858 1930 14904 1964
rect 14858 1914 14938 1930
rect 14117 1899 14167 1900
rect 13750 1831 13796 1865
rect 13964 1865 13998 1869
rect 14248 1869 14450 1903
rect 13964 1847 14181 1865
rect 13750 1797 13830 1831
rect 13864 1801 13880 1835
rect 13914 1801 13930 1835
rect 13864 1763 13930 1801
rect 13964 1813 14147 1847
rect 13964 1797 14181 1813
rect 14248 1852 14282 1869
rect 14416 1852 14450 1869
rect 14248 1797 14282 1818
rect 14316 1801 14332 1835
rect 14366 1801 14382 1835
rect 14316 1763 14382 1801
rect 14591 1869 14806 1903
rect 14977 1901 15095 1965
rect 15129 1952 15181 1993
rect 15163 1928 15181 1952
rect 14977 1877 15011 1901
rect 14591 1852 14638 1869
rect 14416 1797 14450 1818
rect 14484 1805 14500 1839
rect 14534 1805 14550 1839
rect 14484 1763 14550 1805
rect 14591 1818 14604 1852
rect 14772 1852 14806 1869
rect 14591 1797 14638 1818
rect 14672 1801 14688 1835
rect 14722 1801 14738 1835
rect 14672 1763 14738 1801
rect 14772 1797 14806 1818
rect 14856 1852 15011 1877
rect 15129 1892 15140 1918
rect 15174 1892 15181 1928
rect 14890 1818 15011 1852
rect 14856 1797 15011 1818
rect 15045 1843 15095 1860
rect 15079 1809 15095 1843
rect 15045 1763 15095 1809
rect 15129 1858 15181 1892
rect 15163 1824 15181 1858
rect 15129 1797 15181 1824
rect 15814 2195 15894 2239
rect 15943 2235 16009 2273
rect 15943 2201 15959 2235
rect 15993 2201 16009 2235
rect 16043 2223 16245 2239
rect 15814 2161 15860 2195
rect 16043 2189 16211 2223
rect 16043 2167 16077 2189
rect 16211 2171 16245 2189
rect 16312 2218 16346 2239
rect 16380 2235 16446 2273
rect 16380 2201 16396 2235
rect 16430 2201 16446 2235
rect 16480 2218 16514 2239
rect 15814 2128 15894 2161
rect 15929 2133 16077 2167
rect 16312 2167 16346 2184
rect 16548 2226 16614 2273
rect 16548 2192 16564 2226
rect 16598 2192 16614 2226
rect 16668 2218 16702 2239
rect 16480 2167 16514 2184
rect 15814 1993 15880 2128
rect 15929 2091 15963 2133
rect 15914 2075 15963 2091
rect 16170 2103 16182 2137
rect 16216 2103 16269 2137
rect 16312 2133 16514 2167
rect 16736 2235 16802 2273
rect 16736 2201 16752 2235
rect 16786 2201 16802 2235
rect 16836 2218 16870 2239
rect 16668 2167 16702 2184
rect 16836 2167 16870 2184
rect 16668 2133 16870 2167
rect 16920 2218 17040 2239
rect 16954 2184 17040 2218
rect 17093 2231 17159 2273
rect 17093 2197 17109 2231
rect 17143 2197 17159 2231
rect 16920 2163 17040 2184
rect 17193 2195 17245 2239
rect 16920 2137 17159 2163
rect 16920 2103 16922 2137
rect 16956 2129 17159 2137
rect 16956 2103 16968 2129
rect 16170 2099 16269 2103
rect 15948 2041 15963 2075
rect 15914 2025 15963 2041
rect 15997 2069 16013 2083
rect 15997 2035 15998 2069
rect 16047 2049 16085 2083
rect 16170 2065 16253 2099
rect 16287 2065 16303 2099
rect 16337 2065 16353 2099
rect 16387 2069 16412 2099
rect 16032 2035 16085 2049
rect 16337 2035 16366 2065
rect 16400 2035 16412 2069
rect 16471 2040 16704 2097
rect 17125 2091 17159 2129
rect 17227 2161 17245 2195
rect 17193 2124 17245 2161
rect 15814 1955 15894 1993
rect 15814 1921 15860 1955
rect 15814 1865 15894 1921
rect 15929 1903 15963 2025
rect 16051 1971 16090 2001
rect 16051 1937 16085 1971
rect 16124 1967 16135 2001
rect 16471 1987 16505 2040
rect 16119 1937 16135 1967
rect 16181 1971 16438 1987
rect 16215 1953 16438 1971
rect 16472 1953 16505 1987
rect 16550 2001 16622 2003
rect 16584 1987 16622 2001
rect 16550 1953 16555 1967
rect 16589 1953 16622 1987
rect 16215 1937 16231 1953
rect 16550 1937 16622 1953
rect 16670 1971 16704 2040
rect 16738 2069 16816 2084
rect 17014 2075 17080 2091
rect 17014 2069 17046 2075
rect 16772 2068 16816 2069
rect 16772 2035 16782 2068
rect 16738 2034 16782 2035
rect 16738 2018 16816 2034
rect 16854 2035 16878 2069
rect 16912 2035 16928 2069
rect 17048 2035 17080 2041
rect 16854 1971 16888 2035
rect 17046 2025 17080 2035
rect 17125 2075 17176 2091
rect 17125 2041 17142 2075
rect 17125 2025 17176 2041
rect 16670 1937 16888 1971
rect 16956 1967 17002 2001
rect 16922 1964 17002 1967
rect 17125 1965 17159 2025
rect 17210 1993 17245 2124
rect 16181 1934 16231 1937
rect 15929 1869 16062 1903
rect 16181 1900 16188 1934
rect 16222 1900 16231 1934
rect 16922 1930 16968 1964
rect 16922 1914 17002 1930
rect 16181 1899 16231 1900
rect 15814 1831 15860 1865
rect 16028 1865 16062 1869
rect 16312 1869 16514 1903
rect 16028 1847 16245 1865
rect 15814 1797 15894 1831
rect 15928 1801 15944 1835
rect 15978 1801 15994 1835
rect 15928 1763 15994 1801
rect 16028 1813 16211 1847
rect 16028 1797 16245 1813
rect 16312 1852 16346 1869
rect 16480 1852 16514 1869
rect 16312 1797 16346 1818
rect 16380 1801 16396 1835
rect 16430 1801 16446 1835
rect 16380 1763 16446 1801
rect 16655 1869 16870 1903
rect 17041 1901 17159 1965
rect 17193 1952 17245 1993
rect 17227 1928 17245 1952
rect 17041 1877 17075 1901
rect 16655 1852 16702 1869
rect 16480 1797 16514 1818
rect 16548 1805 16564 1839
rect 16598 1805 16614 1839
rect 16548 1763 16614 1805
rect 16655 1818 16668 1852
rect 16836 1852 16870 1869
rect 16655 1797 16702 1818
rect 16736 1801 16752 1835
rect 16786 1801 16802 1835
rect 16736 1763 16802 1801
rect 16836 1797 16870 1818
rect 16920 1852 17075 1877
rect 17193 1892 17204 1918
rect 17238 1892 17245 1928
rect 16954 1818 17075 1852
rect 16920 1797 17075 1818
rect 17109 1843 17159 1860
rect 17143 1809 17159 1843
rect 17109 1763 17159 1809
rect 17193 1858 17245 1892
rect 17227 1824 17245 1858
rect 17193 1797 17245 1824
rect 3876 1723 3905 1757
rect 3939 1723 3997 1757
rect 4031 1723 4089 1757
rect 4123 1723 4181 1757
rect 4215 1723 4273 1757
rect 4307 1723 4365 1757
rect 4399 1723 4457 1757
rect 4491 1723 4549 1757
rect 4583 1723 4641 1757
rect 4675 1723 4733 1757
rect 4767 1723 4825 1757
rect 4859 1723 4917 1757
rect 4951 1723 5009 1757
rect 5043 1723 5101 1757
rect 5135 1723 5193 1757
rect 5227 1723 5285 1757
rect 5319 1723 5348 1757
rect 5828 1723 5857 1757
rect 5891 1723 5949 1757
rect 5983 1723 6041 1757
rect 6075 1723 6133 1757
rect 6167 1723 6225 1757
rect 6259 1723 6317 1757
rect 6351 1723 6409 1757
rect 6443 1723 6501 1757
rect 6535 1723 6593 1757
rect 6627 1723 6685 1757
rect 6719 1723 6777 1757
rect 6811 1723 6869 1757
rect 6903 1723 6961 1757
rect 6995 1723 7053 1757
rect 7087 1723 7145 1757
rect 7179 1723 7237 1757
rect 7271 1723 7300 1757
rect 7830 1729 7859 1763
rect 7893 1729 7951 1763
rect 7985 1729 8043 1763
rect 8077 1729 8135 1763
rect 8169 1729 8227 1763
rect 8261 1729 8319 1763
rect 8353 1729 8411 1763
rect 8445 1729 8503 1763
rect 8537 1729 8595 1763
rect 8629 1729 8687 1763
rect 8721 1729 8779 1763
rect 8813 1729 8871 1763
rect 8905 1729 8963 1763
rect 8997 1729 9055 1763
rect 9089 1729 9147 1763
rect 9181 1729 9239 1763
rect 9273 1729 9302 1763
rect 9782 1729 9811 1763
rect 9845 1729 9903 1763
rect 9937 1729 9995 1763
rect 10029 1729 10087 1763
rect 10121 1729 10179 1763
rect 10213 1729 10271 1763
rect 10305 1729 10363 1763
rect 10397 1729 10455 1763
rect 10489 1729 10547 1763
rect 10581 1729 10639 1763
rect 10673 1729 10731 1763
rect 10765 1729 10823 1763
rect 10857 1729 10915 1763
rect 10949 1729 11007 1763
rect 11041 1729 11099 1763
rect 11133 1729 11191 1763
rect 11225 1729 11254 1763
rect 11774 1729 11803 1763
rect 11837 1729 11895 1763
rect 11929 1729 11987 1763
rect 12021 1729 12079 1763
rect 12113 1729 12171 1763
rect 12205 1729 12263 1763
rect 12297 1729 12355 1763
rect 12389 1729 12447 1763
rect 12481 1729 12539 1763
rect 12573 1729 12631 1763
rect 12665 1729 12723 1763
rect 12757 1729 12815 1763
rect 12849 1729 12907 1763
rect 12941 1729 12999 1763
rect 13033 1729 13091 1763
rect 13125 1729 13183 1763
rect 13217 1729 13246 1763
rect 13726 1729 13755 1763
rect 13789 1729 13847 1763
rect 13881 1729 13939 1763
rect 13973 1729 14031 1763
rect 14065 1729 14123 1763
rect 14157 1729 14215 1763
rect 14249 1729 14307 1763
rect 14341 1729 14399 1763
rect 14433 1729 14491 1763
rect 14525 1729 14583 1763
rect 14617 1729 14675 1763
rect 14709 1729 14767 1763
rect 14801 1729 14859 1763
rect 14893 1729 14951 1763
rect 14985 1729 15043 1763
rect 15077 1729 15135 1763
rect 15169 1729 15198 1763
rect 15790 1729 15819 1763
rect 15853 1729 15911 1763
rect 15945 1729 16003 1763
rect 16037 1729 16095 1763
rect 16129 1729 16187 1763
rect 16221 1729 16279 1763
rect 16313 1729 16371 1763
rect 16405 1729 16463 1763
rect 16497 1729 16555 1763
rect 16589 1729 16647 1763
rect 16681 1729 16739 1763
rect 16773 1729 16831 1763
rect 16865 1729 16923 1763
rect 16957 1729 17015 1763
rect 17049 1729 17107 1763
rect 17141 1729 17199 1763
rect 17233 1729 17262 1763
<< viali >>
rect 9496 17532 9532 17568
rect 9596 17536 9632 17572
rect 9363 16573 9397 16607
rect 9455 16573 9489 16607
rect 9547 16573 9581 16607
rect 9639 16573 9673 16607
rect 9731 16573 9765 16607
rect 9823 16573 9857 16607
rect 9915 16573 9949 16607
rect 9910 16387 9944 16394
rect 9910 16356 9935 16387
rect 9935 16356 9944 16387
rect 16416 16366 16452 16400
rect 16502 16354 16540 16388
rect 17184 16358 17222 16392
rect 9420 16295 9454 16296
rect 9420 16262 9453 16295
rect 9453 16262 9454 16295
rect 9540 16295 9574 16298
rect 9540 16264 9570 16295
rect 9570 16264 9574 16295
rect 17278 16350 17312 16384
rect 18048 16362 18082 16396
rect 18150 16358 18186 16392
rect 18672 16356 18708 16390
rect 18758 16344 18796 16378
rect 19440 16348 19478 16382
rect 19534 16340 19568 16374
rect 20304 16352 20338 16386
rect 20406 16348 20442 16382
rect 21436 16350 21472 16384
rect 21522 16338 21560 16372
rect 22204 16342 22242 16376
rect 22298 16334 22332 16368
rect 23068 16346 23102 16380
rect 23170 16342 23206 16376
rect 9363 16029 9397 16063
rect 9455 16029 9489 16063
rect 9547 16029 9581 16063
rect 9639 16029 9673 16063
rect 9731 16029 9765 16063
rect 9823 16029 9857 16063
rect 9915 16029 9949 16063
rect 9461 15829 9495 15863
rect 9553 15829 9587 15863
rect 9645 15829 9679 15863
rect 9737 15829 9771 15863
rect 9829 15829 9863 15863
rect 11503 15719 11537 15753
rect 11595 15719 11629 15753
rect 11687 15719 11721 15753
rect 11779 15719 11813 15753
rect 11871 15719 11905 15753
rect 11963 15719 11997 15753
rect 12055 15719 12089 15753
rect 9454 15534 9496 15574
rect 9644 15551 9686 15564
rect 9644 15524 9647 15551
rect 9647 15524 9681 15551
rect 9681 15524 9686 15551
rect 9836 15460 9872 15494
rect 11498 15368 11534 15404
rect 9461 15285 9495 15319
rect 9553 15285 9587 15319
rect 9645 15285 9679 15319
rect 9737 15285 9771 15319
rect 9829 15285 9863 15319
rect 11670 15407 11685 15438
rect 11685 15407 11704 15438
rect 11670 15402 11704 15407
rect 11768 15280 11802 15314
rect 11864 15348 11898 15384
rect 12056 15402 12090 15436
rect 10645 15219 10679 15253
rect 10737 15219 10771 15253
rect 10829 15219 10863 15253
rect 10921 15219 10955 15253
rect 11013 15219 11047 15253
rect 9373 15009 9407 15043
rect 9465 15009 9499 15043
rect 9557 15009 9591 15043
rect 9649 15009 9683 15043
rect 9741 15009 9775 15043
rect 9833 15009 9867 15043
rect 9925 15009 9959 15043
rect 11503 15175 11537 15209
rect 11595 15175 11629 15209
rect 11687 15175 11721 15209
rect 11779 15175 11813 15209
rect 11871 15175 11905 15209
rect 11963 15175 11997 15209
rect 12055 15175 12089 15209
rect 11010 15143 11017 15152
rect 11017 15143 11050 15152
rect 11010 15116 11050 15143
rect 9922 14925 9945 14934
rect 9945 14925 9956 14934
rect 9922 14900 9956 14925
rect 10690 14941 10724 14942
rect 10690 14908 10724 14941
rect 10830 14941 10866 14942
rect 10830 14908 10831 14941
rect 10831 14908 10865 14941
rect 10865 14908 10866 14941
rect 9430 14731 9464 14732
rect 9430 14698 9463 14731
rect 9463 14698 9464 14731
rect 9550 14731 9584 14734
rect 9550 14700 9580 14731
rect 9580 14700 9584 14731
rect 10645 14675 10679 14709
rect 10737 14675 10771 14709
rect 10829 14675 10863 14709
rect 10921 14675 10955 14709
rect 11013 14675 11047 14709
rect 24150 14616 24186 14650
rect 23530 14546 23568 14580
rect 23672 14528 23708 14562
rect 24556 14554 24592 14588
rect 25364 14562 25400 14598
rect 24456 14518 24492 14552
rect 24712 14528 24746 14562
rect 9373 14465 9407 14499
rect 9465 14465 9499 14499
rect 9557 14465 9591 14499
rect 9649 14465 9683 14499
rect 9741 14465 9775 14499
rect 9833 14465 9867 14499
rect 9925 14465 9959 14499
rect 9471 14265 9505 14299
rect 9563 14265 9597 14299
rect 9655 14265 9689 14299
rect 9747 14265 9781 14299
rect 9839 14265 9873 14299
rect 10719 14253 10753 14287
rect 10811 14253 10845 14287
rect 10903 14253 10937 14287
rect 10995 14253 11029 14287
rect 11087 14253 11121 14287
rect 11179 14253 11213 14287
rect 11271 14253 11305 14287
rect 8212 14036 8254 14076
rect 9464 13970 9506 14010
rect 9654 13987 9696 14000
rect 9654 13960 9657 13987
rect 9657 13960 9691 13987
rect 9691 13960 9696 13987
rect 7752 13904 7792 13938
rect 9844 13854 9880 13888
rect 12617 14237 12651 14271
rect 12709 14237 12743 14271
rect 12801 14237 12835 14271
rect 12893 14237 12927 14271
rect 12985 14237 13019 14271
rect 13077 14237 13111 14271
rect 12762 14136 12798 14170
rect 10716 13975 10750 13980
rect 10716 13946 10721 13975
rect 10721 13946 10750 13975
rect 10886 13850 10920 13884
rect 10984 13890 11018 13924
rect 11078 13941 11103 13974
rect 11103 13941 11114 13974
rect 11078 13936 11114 13941
rect 13078 14062 13103 14080
rect 13103 14062 13120 14080
rect 11260 13853 11265 13856
rect 11265 13853 11298 13856
rect 11689 13879 11723 13913
rect 11781 13879 11815 13913
rect 11873 13879 11907 13913
rect 11965 13879 11999 13913
rect 12057 13879 12091 13913
rect 12618 13925 12623 13942
rect 12623 13925 12657 13942
rect 12657 13925 12658 13942
rect 12618 13908 12658 13925
rect 13078 14040 13120 14062
rect 12746 13959 12796 13964
rect 12746 13925 12749 13959
rect 12749 13925 12783 13959
rect 12783 13925 12796 13959
rect 12746 13922 12796 13925
rect 12918 13959 12956 13960
rect 12918 13925 12925 13959
rect 12925 13925 12956 13959
rect 12918 13924 12956 13925
rect 11260 13819 11298 13853
rect 11260 13818 11265 13819
rect 11265 13818 11298 13819
rect 9471 13721 9505 13755
rect 9563 13721 9597 13755
rect 9655 13721 9689 13755
rect 9747 13721 9781 13755
rect 9839 13721 9873 13755
rect 10719 13709 10753 13743
rect 10811 13709 10845 13743
rect 10903 13709 10937 13743
rect 10995 13709 11029 13743
rect 11087 13709 11121 13743
rect 11179 13709 11213 13743
rect 11271 13709 11305 13743
rect 12028 13735 12039 13768
rect 12039 13735 12062 13768
rect 12028 13734 12062 13735
rect 11700 13524 11734 13558
rect 11878 13601 11912 13608
rect 11878 13574 11896 13601
rect 11896 13574 11912 13601
rect 12617 13693 12651 13727
rect 12709 13693 12743 13727
rect 12801 13693 12835 13727
rect 12893 13693 12927 13727
rect 12985 13693 13019 13727
rect 13077 13693 13111 13727
rect 10843 13411 10877 13445
rect 10935 13411 10969 13445
rect 11027 13411 11061 13445
rect 11119 13411 11153 13445
rect 11211 13411 11245 13445
rect 9365 13341 9399 13375
rect 9457 13341 9491 13375
rect 9549 13341 9583 13375
rect 9641 13341 9675 13375
rect 9733 13341 9767 13375
rect 9825 13341 9859 13375
rect 9917 13341 9951 13375
rect 11012 13326 11021 13338
rect 11021 13326 11048 13338
rect 11012 13302 11048 13326
rect 11689 13335 11723 13369
rect 11781 13335 11815 13369
rect 11873 13335 11907 13369
rect 11965 13335 11999 13369
rect 12057 13335 12091 13369
rect 9914 13223 9948 13224
rect 9914 13190 9937 13223
rect 9937 13190 9948 13223
rect 11208 13253 11239 13282
rect 11239 13253 11246 13282
rect 11208 13244 11246 13253
rect 9422 13063 9456 13064
rect 9422 13030 9455 13063
rect 9455 13030 9456 13063
rect 9542 13063 9576 13066
rect 9542 13032 9572 13063
rect 9572 13032 9576 13063
rect 10860 13053 10883 13064
rect 10883 13053 10894 13064
rect 10860 13030 10894 13053
rect 11062 13036 11098 13070
rect 10843 12867 10877 12901
rect 10935 12867 10969 12901
rect 11027 12867 11061 12901
rect 11119 12867 11153 12901
rect 11211 12867 11245 12901
rect 9365 12797 9399 12831
rect 9457 12797 9491 12831
rect 9549 12797 9583 12831
rect 9641 12797 9675 12831
rect 9733 12797 9767 12831
rect 9825 12797 9859 12831
rect 9917 12797 9951 12831
rect 9463 12597 9497 12631
rect 9555 12597 9589 12631
rect 9647 12597 9681 12631
rect 9739 12597 9773 12631
rect 9831 12597 9865 12631
rect 9456 12302 9498 12342
rect 10839 12391 10873 12425
rect 10931 12391 10965 12425
rect 11023 12391 11057 12425
rect 11115 12391 11149 12425
rect 11207 12391 11241 12425
rect 9836 12340 9872 12374
rect 9646 12319 9688 12332
rect 9646 12292 9649 12319
rect 9649 12292 9683 12319
rect 9683 12292 9688 12319
rect 11212 12166 11246 12200
rect 9463 12053 9497 12087
rect 9555 12053 9589 12087
rect 9647 12053 9681 12087
rect 9739 12053 9773 12087
rect 9831 12053 9865 12087
rect 10884 12113 10920 12116
rect 10884 12082 10918 12113
rect 10918 12082 10920 12113
rect 11024 12113 11060 12114
rect 11024 12080 11025 12113
rect 11025 12080 11059 12113
rect 11059 12080 11060 12113
rect 10839 11847 10873 11881
rect 10931 11847 10965 11881
rect 11023 11847 11057 11881
rect 11115 11847 11149 11881
rect 11207 11847 11241 11881
rect 9375 11777 9409 11811
rect 9467 11777 9501 11811
rect 9559 11777 9593 11811
rect 9651 11777 9685 11811
rect 9743 11777 9777 11811
rect 9835 11777 9869 11811
rect 9927 11777 9961 11811
rect 9914 11659 9950 11660
rect 9914 11626 9947 11659
rect 9947 11626 9950 11659
rect 9432 11499 9466 11500
rect 9432 11466 9465 11499
rect 9465 11466 9466 11499
rect 9552 11499 9586 11502
rect 9552 11468 9582 11499
rect 9582 11468 9586 11499
rect 9375 11233 9409 11267
rect 9467 11233 9501 11267
rect 9559 11233 9593 11267
rect 9651 11233 9685 11267
rect 9743 11233 9777 11267
rect 9835 11233 9869 11267
rect 9927 11233 9961 11267
rect 9473 11033 9507 11067
rect 9565 11033 9599 11067
rect 9657 11033 9691 11067
rect 9749 11033 9783 11067
rect 9841 11033 9875 11067
rect 9466 10738 9508 10778
rect 4982 10694 5016 10730
rect 9656 10755 9698 10768
rect 9656 10728 9659 10755
rect 9659 10728 9693 10755
rect 9693 10728 9698 10755
rect 9848 10698 9882 10734
rect 9473 10489 9507 10523
rect 9565 10489 9599 10523
rect 9657 10489 9691 10523
rect 9749 10489 9783 10523
rect 9841 10489 9875 10523
rect 6141 6583 6175 6617
rect 6233 6583 6267 6617
rect 6325 6583 6359 6617
rect 6178 6348 6212 6382
rect 6274 6351 6308 6384
rect 6274 6350 6308 6351
rect 6141 6039 6175 6073
rect 6233 6039 6267 6073
rect 6325 6039 6359 6073
rect 10047 5951 10081 5985
rect 10139 5951 10173 5985
rect 10231 5951 10265 5985
rect 10323 5951 10357 5985
rect 10415 5951 10449 5985
rect 10507 5951 10541 5985
rect 10599 5951 10633 5985
rect 10691 5951 10725 5985
rect 10783 5951 10817 5985
rect 10875 5951 10909 5985
rect 10967 5951 11001 5985
rect 11059 5951 11093 5985
rect 11151 5951 11185 5985
rect 11243 5951 11277 5985
rect 11335 5951 11369 5985
rect 11427 5951 11461 5985
rect 10410 5781 10444 5815
rect 12109 5939 12143 5973
rect 12201 5939 12235 5973
rect 12293 5939 12327 5973
rect 12385 5939 12419 5973
rect 12477 5939 12511 5973
rect 12569 5939 12603 5973
rect 12661 5939 12695 5973
rect 12753 5939 12787 5973
rect 12845 5939 12879 5973
rect 12937 5939 12971 5973
rect 13029 5939 13063 5973
rect 13121 5939 13155 5973
rect 13213 5939 13247 5973
rect 13305 5939 13339 5973
rect 13397 5939 13431 5973
rect 13489 5939 13523 5973
rect 14067 5947 14101 5981
rect 14159 5947 14193 5981
rect 14251 5947 14285 5981
rect 14343 5947 14377 5981
rect 14435 5947 14469 5981
rect 14527 5947 14561 5981
rect 14619 5947 14653 5981
rect 14711 5947 14745 5981
rect 14803 5947 14837 5981
rect 14895 5947 14929 5981
rect 14987 5947 15021 5981
rect 15079 5947 15113 5981
rect 15171 5947 15205 5981
rect 15263 5947 15297 5981
rect 15355 5947 15389 5981
rect 15447 5947 15481 5981
rect 16061 5953 16095 5987
rect 16153 5953 16187 5987
rect 16245 5953 16279 5987
rect 16337 5953 16371 5987
rect 16429 5953 16463 5987
rect 16521 5953 16555 5987
rect 16613 5953 16647 5987
rect 16705 5953 16739 5987
rect 16797 5953 16831 5987
rect 16889 5953 16923 5987
rect 16981 5953 17015 5987
rect 17073 5953 17107 5987
rect 17165 5953 17199 5987
rect 17257 5953 17291 5987
rect 17349 5953 17383 5987
rect 17441 5953 17475 5987
rect 11150 5781 11184 5815
rect 10226 5727 10241 5747
rect 10241 5727 10260 5747
rect 10594 5743 10615 5747
rect 10615 5743 10628 5747
rect 10226 5713 10260 5727
rect 10594 5713 10628 5743
rect 1865 5531 1899 5565
rect 1957 5531 1991 5565
rect 2049 5531 2083 5565
rect 2141 5531 2175 5565
rect 2233 5531 2267 5565
rect 2325 5531 2359 5565
rect 2417 5531 2451 5565
rect 2509 5531 2543 5565
rect 2601 5531 2635 5565
rect 2693 5531 2727 5565
rect 2785 5531 2819 5565
rect 2877 5531 2911 5565
rect 2969 5531 3003 5565
rect 3061 5531 3095 5565
rect 3153 5531 3187 5565
rect 3245 5531 3279 5565
rect 2228 5361 2262 5395
rect 3999 5523 4033 5557
rect 4091 5523 4125 5557
rect 4183 5523 4217 5557
rect 4275 5523 4309 5557
rect 4367 5523 4401 5557
rect 4459 5523 4493 5557
rect 4551 5523 4585 5557
rect 4643 5523 4677 5557
rect 4735 5523 4769 5557
rect 4827 5523 4861 5557
rect 4919 5523 4953 5557
rect 5011 5523 5045 5557
rect 5103 5523 5137 5557
rect 5195 5523 5229 5557
rect 5287 5523 5321 5557
rect 5379 5523 5413 5557
rect 5951 5523 5985 5557
rect 6043 5523 6077 5557
rect 6135 5523 6169 5557
rect 6227 5523 6261 5557
rect 6319 5523 6353 5557
rect 6411 5523 6445 5557
rect 6503 5523 6537 5557
rect 6595 5523 6629 5557
rect 6687 5523 6721 5557
rect 6779 5523 6813 5557
rect 6871 5523 6905 5557
rect 6963 5523 6997 5557
rect 7055 5523 7089 5557
rect 7147 5523 7181 5557
rect 7239 5523 7273 5557
rect 7331 5523 7365 5557
rect 7953 5529 7987 5563
rect 8045 5529 8079 5563
rect 8137 5529 8171 5563
rect 8229 5529 8263 5563
rect 8321 5529 8355 5563
rect 8413 5529 8447 5563
rect 8505 5529 8539 5563
rect 8597 5529 8631 5563
rect 8689 5529 8723 5563
rect 8781 5529 8815 5563
rect 8873 5529 8907 5563
rect 8965 5529 8999 5563
rect 9057 5529 9091 5563
rect 9149 5529 9183 5563
rect 9241 5529 9275 5563
rect 9333 5529 9367 5563
rect 10318 5649 10352 5679
rect 10318 5645 10347 5649
rect 10347 5645 10352 5649
rect 10778 5665 10812 5679
rect 10778 5645 10783 5665
rect 10783 5645 10812 5665
rect 10966 5713 11000 5747
rect 11242 5719 11274 5747
rect 11274 5719 11276 5747
rect 11242 5713 11276 5719
rect 11150 5645 11184 5679
rect 10418 5580 10452 5614
rect 2968 5361 3002 5395
rect 2044 5307 2059 5327
rect 2059 5307 2078 5327
rect 2412 5323 2433 5327
rect 2433 5323 2446 5327
rect 2044 5293 2078 5307
rect 2412 5293 2446 5323
rect 2136 5229 2170 5259
rect 2136 5225 2165 5229
rect 2165 5225 2170 5229
rect 2596 5245 2630 5259
rect 2596 5225 2601 5245
rect 2601 5225 2630 5245
rect 2784 5293 2818 5327
rect 3060 5299 3092 5327
rect 3092 5299 3094 5327
rect 3060 5293 3094 5299
rect 2968 5225 3002 5259
rect 2236 5160 2270 5194
rect 3244 5176 3273 5186
rect 3273 5176 3284 5186
rect 3244 5150 3284 5176
rect 4362 5353 4396 5387
rect 5102 5353 5136 5387
rect 4178 5299 4193 5319
rect 4193 5299 4212 5319
rect 4546 5315 4567 5319
rect 4567 5315 4580 5319
rect 4178 5285 4212 5299
rect 4546 5285 4580 5315
rect 4270 5221 4304 5251
rect 4270 5217 4299 5221
rect 4299 5217 4304 5221
rect 4730 5237 4764 5251
rect 4730 5217 4735 5237
rect 4735 5217 4764 5237
rect 4918 5285 4952 5319
rect 5194 5291 5226 5319
rect 5226 5291 5228 5319
rect 5194 5285 5228 5291
rect 5102 5217 5136 5251
rect 4368 5150 4402 5184
rect 1865 4987 1899 5021
rect 1957 4987 1991 5021
rect 2049 4987 2083 5021
rect 2141 4987 2175 5021
rect 2233 4987 2267 5021
rect 2325 4987 2359 5021
rect 2417 4987 2451 5021
rect 2509 4987 2543 5021
rect 2601 4987 2635 5021
rect 2693 4987 2727 5021
rect 2785 4987 2819 5021
rect 2877 4987 2911 5021
rect 2969 4987 3003 5021
rect 3061 4987 3095 5021
rect 3153 4987 3187 5021
rect 3245 4987 3279 5021
rect 5384 5168 5407 5178
rect 5407 5168 5418 5178
rect 5384 5142 5418 5168
rect 6314 5353 6348 5387
rect 7054 5353 7088 5387
rect 6130 5299 6145 5319
rect 6145 5299 6164 5319
rect 6498 5315 6519 5319
rect 6519 5315 6532 5319
rect 6130 5285 6164 5299
rect 6498 5285 6532 5315
rect 6222 5221 6256 5251
rect 6222 5217 6251 5221
rect 6251 5217 6256 5221
rect 6682 5237 6716 5251
rect 6682 5217 6687 5237
rect 6687 5217 6716 5237
rect 6870 5285 6904 5319
rect 7146 5291 7178 5319
rect 7178 5291 7180 5319
rect 7146 5285 7180 5291
rect 7054 5217 7088 5251
rect 6320 5150 6354 5184
rect 7336 5168 7359 5178
rect 7359 5168 7370 5178
rect 7336 5142 7370 5168
rect 8316 5359 8350 5393
rect 9056 5359 9090 5393
rect 8132 5305 8147 5325
rect 8147 5305 8166 5325
rect 8500 5321 8521 5325
rect 8521 5321 8534 5325
rect 8132 5291 8166 5305
rect 8500 5291 8534 5321
rect 11426 5596 11455 5606
rect 11455 5596 11466 5606
rect 11426 5570 11466 5596
rect 12472 5769 12506 5803
rect 13212 5769 13246 5803
rect 12288 5715 12303 5735
rect 12303 5715 12322 5735
rect 12656 5731 12677 5735
rect 12677 5731 12690 5735
rect 12288 5701 12322 5715
rect 12656 5701 12690 5731
rect 12380 5637 12414 5667
rect 12380 5633 12409 5637
rect 12409 5633 12414 5637
rect 12840 5653 12874 5667
rect 12840 5633 12845 5653
rect 12845 5633 12874 5653
rect 13028 5701 13062 5735
rect 13304 5707 13336 5735
rect 13336 5707 13338 5735
rect 13304 5701 13338 5707
rect 13212 5633 13246 5667
rect 12478 5566 12512 5600
rect 10047 5407 10081 5441
rect 10139 5407 10173 5441
rect 10231 5407 10265 5441
rect 10323 5407 10357 5441
rect 10415 5407 10449 5441
rect 10507 5407 10541 5441
rect 10599 5407 10633 5441
rect 10691 5407 10725 5441
rect 10783 5407 10817 5441
rect 10875 5407 10909 5441
rect 10967 5407 11001 5441
rect 11059 5407 11093 5441
rect 11151 5407 11185 5441
rect 11243 5407 11277 5441
rect 11335 5407 11369 5441
rect 11427 5407 11461 5441
rect 13494 5584 13517 5594
rect 13517 5584 13528 5594
rect 13494 5558 13528 5584
rect 14430 5777 14464 5811
rect 15170 5777 15204 5811
rect 14246 5723 14261 5743
rect 14261 5723 14280 5743
rect 14614 5739 14635 5743
rect 14635 5739 14648 5743
rect 14246 5709 14280 5723
rect 14614 5709 14648 5739
rect 14338 5645 14372 5675
rect 14338 5641 14367 5645
rect 14367 5641 14372 5645
rect 14798 5661 14832 5675
rect 14798 5641 14803 5661
rect 14803 5641 14832 5661
rect 14986 5709 15020 5743
rect 15262 5715 15294 5743
rect 15294 5715 15296 5743
rect 15262 5709 15296 5715
rect 15170 5641 15204 5675
rect 14436 5574 14470 5608
rect 15452 5592 15475 5602
rect 15475 5592 15486 5602
rect 15452 5566 15486 5592
rect 16424 5783 16458 5817
rect 17164 5783 17198 5817
rect 16240 5729 16255 5749
rect 16255 5729 16274 5749
rect 16608 5745 16629 5749
rect 16629 5745 16642 5749
rect 16240 5715 16274 5729
rect 16608 5715 16642 5745
rect 16332 5651 16366 5681
rect 16332 5647 16361 5651
rect 16361 5647 16366 5651
rect 16792 5667 16826 5681
rect 16792 5647 16797 5667
rect 16797 5647 16826 5667
rect 16980 5715 17014 5749
rect 17256 5721 17288 5749
rect 17288 5721 17290 5749
rect 17256 5715 17290 5721
rect 17164 5647 17198 5681
rect 16430 5580 16464 5614
rect 17446 5598 17469 5608
rect 17469 5598 17480 5608
rect 17446 5572 17480 5598
rect 12109 5395 12143 5429
rect 12201 5395 12235 5429
rect 12293 5395 12327 5429
rect 12385 5395 12419 5429
rect 12477 5395 12511 5429
rect 12569 5395 12603 5429
rect 12661 5395 12695 5429
rect 12753 5395 12787 5429
rect 12845 5395 12879 5429
rect 12937 5395 12971 5429
rect 13029 5395 13063 5429
rect 13121 5395 13155 5429
rect 13213 5395 13247 5429
rect 13305 5395 13339 5429
rect 13397 5395 13431 5429
rect 13489 5395 13523 5429
rect 14067 5403 14101 5437
rect 14159 5403 14193 5437
rect 14251 5403 14285 5437
rect 14343 5403 14377 5437
rect 14435 5403 14469 5437
rect 14527 5403 14561 5437
rect 14619 5403 14653 5437
rect 14711 5403 14745 5437
rect 14803 5403 14837 5437
rect 14895 5403 14929 5437
rect 14987 5403 15021 5437
rect 15079 5403 15113 5437
rect 15171 5403 15205 5437
rect 15263 5403 15297 5437
rect 15355 5403 15389 5437
rect 15447 5403 15481 5437
rect 16061 5409 16095 5443
rect 16153 5409 16187 5443
rect 16245 5409 16279 5443
rect 16337 5409 16371 5443
rect 16429 5409 16463 5443
rect 16521 5409 16555 5443
rect 16613 5409 16647 5443
rect 16705 5409 16739 5443
rect 16797 5409 16831 5443
rect 16889 5409 16923 5443
rect 16981 5409 17015 5443
rect 17073 5409 17107 5443
rect 17165 5409 17199 5443
rect 17257 5409 17291 5443
rect 17349 5409 17383 5443
rect 17441 5409 17475 5443
rect 8224 5227 8258 5257
rect 8224 5223 8253 5227
rect 8253 5223 8258 5227
rect 8684 5243 8718 5257
rect 8684 5223 8689 5243
rect 8689 5223 8718 5243
rect 8872 5291 8906 5325
rect 9148 5297 9180 5325
rect 9180 5297 9182 5325
rect 9148 5291 9182 5297
rect 9056 5223 9090 5257
rect 8322 5156 8356 5190
rect 18608 5188 18642 5222
rect 9338 5174 9361 5184
rect 9361 5174 9372 5184
rect 9338 5148 9372 5174
rect 18690 5160 18724 5194
rect 10075 5077 10109 5111
rect 10167 5077 10201 5111
rect 10259 5077 10293 5111
rect 10351 5077 10385 5111
rect 10443 5077 10477 5111
rect 10535 5077 10569 5111
rect 10627 5077 10661 5111
rect 10719 5077 10753 5111
rect 10811 5077 10845 5111
rect 10903 5077 10937 5111
rect 10995 5077 11029 5111
rect 11087 5077 11121 5111
rect 11179 5077 11213 5111
rect 11271 5077 11305 5111
rect 11363 5077 11397 5111
rect 11455 5077 11489 5111
rect 3999 4979 4033 5013
rect 4091 4979 4125 5013
rect 4183 4979 4217 5013
rect 4275 4979 4309 5013
rect 4367 4979 4401 5013
rect 4459 4979 4493 5013
rect 4551 4979 4585 5013
rect 4643 4979 4677 5013
rect 4735 4979 4769 5013
rect 4827 4979 4861 5013
rect 4919 4979 4953 5013
rect 5011 4979 5045 5013
rect 5103 4979 5137 5013
rect 5195 4979 5229 5013
rect 5287 4979 5321 5013
rect 5379 4979 5413 5013
rect 5951 4979 5985 5013
rect 6043 4979 6077 5013
rect 6135 4979 6169 5013
rect 6227 4979 6261 5013
rect 6319 4979 6353 5013
rect 6411 4979 6445 5013
rect 6503 4979 6537 5013
rect 6595 4979 6629 5013
rect 6687 4979 6721 5013
rect 6779 4979 6813 5013
rect 6871 4979 6905 5013
rect 6963 4979 6997 5013
rect 7055 4979 7089 5013
rect 7147 4979 7181 5013
rect 7239 4979 7273 5013
rect 7331 4979 7365 5013
rect 7953 4985 7987 5019
rect 8045 4985 8079 5019
rect 8137 4985 8171 5019
rect 8229 4985 8263 5019
rect 8321 4985 8355 5019
rect 8413 4985 8447 5019
rect 8505 4985 8539 5019
rect 8597 4985 8631 5019
rect 8689 4985 8723 5019
rect 8781 4985 8815 5019
rect 8873 4985 8907 5019
rect 8965 4985 8999 5019
rect 9057 4985 9091 5019
rect 9149 4985 9183 5019
rect 9241 4985 9275 5019
rect 9333 4985 9367 5019
rect 10438 4907 10472 4941
rect 18432 5070 18470 5108
rect 12345 5033 12379 5067
rect 12437 5033 12471 5067
rect 12529 5033 12563 5067
rect 12621 5033 12655 5067
rect 12713 5033 12747 5067
rect 12805 5033 12839 5067
rect 12897 5033 12931 5067
rect 12989 5033 13023 5067
rect 13081 5033 13115 5067
rect 13173 5033 13207 5067
rect 13265 5033 13299 5067
rect 13357 5033 13391 5067
rect 13449 5033 13483 5067
rect 13541 5033 13575 5067
rect 13633 5033 13667 5067
rect 13725 5033 13759 5067
rect 11178 4907 11212 4941
rect 10254 4853 10269 4873
rect 10269 4853 10288 4873
rect 10622 4869 10643 4873
rect 10643 4869 10656 4873
rect 10254 4839 10288 4853
rect 10622 4839 10656 4869
rect 10346 4775 10380 4805
rect 10346 4771 10375 4775
rect 10375 4771 10380 4775
rect 10806 4791 10840 4805
rect 10806 4771 10811 4791
rect 10811 4771 10840 4791
rect 10994 4839 11028 4873
rect 11270 4845 11302 4873
rect 11302 4845 11304 4873
rect 11270 4839 11304 4845
rect 11178 4771 11212 4805
rect 10446 4706 10480 4740
rect 11454 4722 11483 4732
rect 11483 4722 11494 4732
rect 11454 4696 11494 4722
rect 12708 4863 12742 4897
rect 14347 5027 14381 5061
rect 14439 5027 14473 5061
rect 14531 5027 14565 5061
rect 14623 5027 14657 5061
rect 14715 5027 14749 5061
rect 14807 5027 14841 5061
rect 14899 5027 14933 5061
rect 14991 5027 15025 5061
rect 15083 5027 15117 5061
rect 15175 5027 15209 5061
rect 15267 5027 15301 5061
rect 15359 5027 15393 5061
rect 15451 5027 15485 5061
rect 15543 5027 15577 5061
rect 15635 5027 15669 5061
rect 15727 5027 15761 5061
rect 13448 4863 13482 4897
rect 12524 4809 12539 4829
rect 12539 4809 12558 4829
rect 12892 4825 12913 4829
rect 12913 4825 12926 4829
rect 12524 4795 12558 4809
rect 12892 4795 12926 4825
rect 12616 4731 12650 4761
rect 12616 4727 12645 4731
rect 12645 4727 12650 4731
rect 13076 4747 13110 4761
rect 13076 4727 13081 4747
rect 13081 4727 13110 4747
rect 13264 4795 13298 4829
rect 13540 4801 13572 4829
rect 13572 4801 13574 4829
rect 13540 4795 13574 4801
rect 13448 4727 13482 4761
rect 12714 4660 12748 4694
rect 10075 4533 10109 4567
rect 10167 4533 10201 4567
rect 10259 4533 10293 4567
rect 10351 4533 10385 4567
rect 10443 4533 10477 4567
rect 10535 4533 10569 4567
rect 10627 4533 10661 4567
rect 10719 4533 10753 4567
rect 10811 4533 10845 4567
rect 10903 4533 10937 4567
rect 10995 4533 11029 4567
rect 11087 4533 11121 4567
rect 11179 4533 11213 4567
rect 11271 4533 11305 4567
rect 11363 4533 11397 4567
rect 11455 4533 11489 4567
rect 13730 4678 13753 4688
rect 13753 4678 13764 4688
rect 13730 4652 13764 4678
rect 14710 4857 14744 4891
rect 16369 5009 16403 5043
rect 16461 5009 16495 5043
rect 16553 5009 16587 5043
rect 16645 5009 16679 5043
rect 16737 5009 16771 5043
rect 16829 5009 16863 5043
rect 16921 5009 16955 5043
rect 17013 5009 17047 5043
rect 17105 5009 17139 5043
rect 17197 5009 17231 5043
rect 17289 5009 17323 5043
rect 17381 5009 17415 5043
rect 17473 5009 17507 5043
rect 17565 5009 17599 5043
rect 17657 5009 17691 5043
rect 17749 5009 17783 5043
rect 15450 4857 15484 4891
rect 14526 4803 14541 4823
rect 14541 4803 14560 4823
rect 14894 4819 14915 4823
rect 14915 4819 14928 4823
rect 14526 4789 14560 4803
rect 14894 4789 14928 4819
rect 14618 4725 14652 4755
rect 14618 4721 14647 4725
rect 14647 4721 14652 4725
rect 15078 4741 15112 4755
rect 15078 4721 15083 4741
rect 15083 4721 15112 4741
rect 15266 4789 15300 4823
rect 15542 4795 15574 4823
rect 15574 4795 15576 4823
rect 15542 4789 15576 4795
rect 15450 4721 15484 4755
rect 14716 4654 14750 4688
rect 12345 4489 12379 4523
rect 12437 4489 12471 4523
rect 12529 4489 12563 4523
rect 12621 4489 12655 4523
rect 12713 4489 12747 4523
rect 12805 4489 12839 4523
rect 12897 4489 12931 4523
rect 12989 4489 13023 4523
rect 13081 4489 13115 4523
rect 13173 4489 13207 4523
rect 13265 4489 13299 4523
rect 13357 4489 13391 4523
rect 13449 4489 13483 4523
rect 13541 4489 13575 4523
rect 13633 4489 13667 4523
rect 13725 4489 13759 4523
rect 15732 4672 15755 4682
rect 15755 4672 15766 4682
rect 15732 4646 15766 4672
rect 16732 4839 16766 4873
rect 19064 5004 19102 5042
rect 17472 4839 17506 4873
rect 16548 4785 16563 4805
rect 16563 4785 16582 4805
rect 16916 4801 16937 4805
rect 16937 4801 16950 4805
rect 16548 4771 16582 4785
rect 16916 4771 16950 4801
rect 16640 4707 16674 4737
rect 16640 4703 16669 4707
rect 16669 4703 16674 4707
rect 17100 4723 17134 4737
rect 17100 4703 17105 4723
rect 17105 4703 17134 4723
rect 17288 4771 17322 4805
rect 17564 4777 17596 4805
rect 17596 4777 17598 4805
rect 17564 4771 17598 4777
rect 17472 4703 17506 4737
rect 16738 4636 16772 4670
rect 14347 4483 14381 4517
rect 14439 4483 14473 4517
rect 14531 4483 14565 4517
rect 14623 4483 14657 4517
rect 14715 4483 14749 4517
rect 14807 4483 14841 4517
rect 14899 4483 14933 4517
rect 14991 4483 15025 4517
rect 15083 4483 15117 4517
rect 15175 4483 15209 4517
rect 15267 4483 15301 4517
rect 15359 4483 15393 4517
rect 15451 4483 15485 4517
rect 15543 4483 15577 4517
rect 15635 4483 15669 4517
rect 15727 4483 15761 4517
rect 17754 4654 17777 4664
rect 17777 4654 17788 4664
rect 17754 4628 17788 4654
rect 16369 4465 16403 4499
rect 16461 4465 16495 4499
rect 16553 4465 16587 4499
rect 16645 4465 16679 4499
rect 16737 4465 16771 4499
rect 16829 4465 16863 4499
rect 16921 4465 16955 4499
rect 17013 4465 17047 4499
rect 17105 4465 17139 4499
rect 17197 4465 17231 4499
rect 17289 4465 17323 4499
rect 17381 4465 17415 4499
rect 17473 4465 17507 4499
rect 17565 4465 17599 4499
rect 17657 4465 17691 4499
rect 17749 4465 17783 4499
rect 6148 3088 6182 3122
rect 6244 3090 6278 3124
rect 1835 2271 1869 2305
rect 1927 2271 1961 2305
rect 2019 2271 2053 2305
rect 2111 2271 2145 2305
rect 2203 2271 2237 2305
rect 2295 2271 2329 2305
rect 2387 2271 2421 2305
rect 2479 2271 2513 2305
rect 2571 2271 2605 2305
rect 2663 2271 2697 2305
rect 2755 2271 2789 2305
rect 2847 2271 2881 2305
rect 2939 2271 2973 2305
rect 3031 2271 3065 2305
rect 3123 2271 3157 2305
rect 3215 2271 3249 2305
rect 2198 2101 2232 2135
rect 3905 2267 3939 2301
rect 3997 2267 4031 2301
rect 4089 2267 4123 2301
rect 4181 2267 4215 2301
rect 4273 2267 4307 2301
rect 4365 2267 4399 2301
rect 4457 2267 4491 2301
rect 4549 2267 4583 2301
rect 4641 2267 4675 2301
rect 4733 2267 4767 2301
rect 4825 2267 4859 2301
rect 4917 2267 4951 2301
rect 5009 2267 5043 2301
rect 5101 2267 5135 2301
rect 5193 2267 5227 2301
rect 5285 2267 5319 2301
rect 5857 2267 5891 2301
rect 5949 2267 5983 2301
rect 6041 2267 6075 2301
rect 6133 2267 6167 2301
rect 6225 2267 6259 2301
rect 6317 2267 6351 2301
rect 6409 2267 6443 2301
rect 6501 2267 6535 2301
rect 6593 2267 6627 2301
rect 6685 2267 6719 2301
rect 6777 2267 6811 2301
rect 6869 2267 6903 2301
rect 6961 2267 6995 2301
rect 7053 2267 7087 2301
rect 7145 2267 7179 2301
rect 7237 2267 7271 2301
rect 7859 2273 7893 2307
rect 7951 2273 7985 2307
rect 8043 2273 8077 2307
rect 8135 2273 8169 2307
rect 8227 2273 8261 2307
rect 8319 2273 8353 2307
rect 8411 2273 8445 2307
rect 8503 2273 8537 2307
rect 8595 2273 8629 2307
rect 8687 2273 8721 2307
rect 8779 2273 8813 2307
rect 8871 2273 8905 2307
rect 8963 2273 8997 2307
rect 9055 2273 9089 2307
rect 9147 2273 9181 2307
rect 9239 2273 9273 2307
rect 9811 2273 9845 2307
rect 9903 2273 9937 2307
rect 9995 2273 10029 2307
rect 10087 2273 10121 2307
rect 10179 2273 10213 2307
rect 10271 2273 10305 2307
rect 10363 2273 10397 2307
rect 10455 2273 10489 2307
rect 10547 2273 10581 2307
rect 10639 2273 10673 2307
rect 10731 2273 10765 2307
rect 10823 2273 10857 2307
rect 10915 2273 10949 2307
rect 11007 2273 11041 2307
rect 11099 2273 11133 2307
rect 11191 2273 11225 2307
rect 11803 2273 11837 2307
rect 11895 2273 11929 2307
rect 11987 2273 12021 2307
rect 12079 2273 12113 2307
rect 12171 2273 12205 2307
rect 12263 2273 12297 2307
rect 12355 2273 12389 2307
rect 12447 2273 12481 2307
rect 12539 2273 12573 2307
rect 12631 2273 12665 2307
rect 12723 2273 12757 2307
rect 12815 2273 12849 2307
rect 12907 2273 12941 2307
rect 12999 2273 13033 2307
rect 13091 2273 13125 2307
rect 13183 2273 13217 2307
rect 13755 2273 13789 2307
rect 13847 2273 13881 2307
rect 13939 2273 13973 2307
rect 14031 2273 14065 2307
rect 14123 2273 14157 2307
rect 14215 2273 14249 2307
rect 14307 2273 14341 2307
rect 14399 2273 14433 2307
rect 14491 2273 14525 2307
rect 14583 2273 14617 2307
rect 14675 2273 14709 2307
rect 14767 2273 14801 2307
rect 14859 2273 14893 2307
rect 14951 2273 14985 2307
rect 15043 2273 15077 2307
rect 15135 2273 15169 2307
rect 15819 2273 15853 2307
rect 15911 2273 15945 2307
rect 16003 2273 16037 2307
rect 16095 2273 16129 2307
rect 16187 2273 16221 2307
rect 16279 2273 16313 2307
rect 16371 2273 16405 2307
rect 16463 2273 16497 2307
rect 16555 2273 16589 2307
rect 16647 2273 16681 2307
rect 16739 2273 16773 2307
rect 16831 2273 16865 2307
rect 16923 2273 16957 2307
rect 17015 2273 17049 2307
rect 17107 2273 17141 2307
rect 17199 2273 17233 2307
rect 2938 2101 2972 2135
rect 2014 2047 2029 2067
rect 2029 2047 2048 2067
rect 2382 2063 2403 2067
rect 2403 2063 2416 2067
rect 2014 2033 2048 2047
rect 2382 2033 2416 2063
rect 2106 1969 2140 1999
rect 2106 1965 2135 1969
rect 2135 1965 2140 1969
rect 2566 1985 2600 1999
rect 2566 1965 2571 1985
rect 2571 1965 2600 1985
rect 2754 2033 2788 2067
rect 3030 2039 3062 2067
rect 3062 2039 3064 2067
rect 3030 2033 3064 2039
rect 2938 1965 2972 1999
rect 2206 1900 2240 1934
rect 3214 1916 3243 1926
rect 3243 1916 3254 1926
rect 3214 1890 3254 1916
rect 4268 2097 4302 2131
rect 5008 2097 5042 2131
rect 4084 2043 4099 2063
rect 4099 2043 4118 2063
rect 4452 2059 4473 2063
rect 4473 2059 4486 2063
rect 4084 2029 4118 2043
rect 4452 2029 4486 2059
rect 4176 1965 4210 1995
rect 4176 1961 4205 1965
rect 4205 1961 4210 1965
rect 4636 1981 4670 1995
rect 4636 1961 4641 1981
rect 4641 1961 4670 1981
rect 4824 2029 4858 2063
rect 5100 2035 5132 2063
rect 5132 2035 5134 2063
rect 5100 2029 5134 2035
rect 5008 1961 5042 1995
rect 4274 1894 4308 1928
rect 1835 1727 1869 1761
rect 1927 1727 1961 1761
rect 2019 1727 2053 1761
rect 2111 1727 2145 1761
rect 2203 1727 2237 1761
rect 2295 1727 2329 1761
rect 2387 1727 2421 1761
rect 2479 1727 2513 1761
rect 2571 1727 2605 1761
rect 2663 1727 2697 1761
rect 2755 1727 2789 1761
rect 2847 1727 2881 1761
rect 2939 1727 2973 1761
rect 3031 1727 3065 1761
rect 3123 1727 3157 1761
rect 3215 1727 3249 1761
rect 5290 1912 5313 1922
rect 5313 1912 5324 1922
rect 5290 1886 5324 1912
rect 6220 2097 6254 2131
rect 6960 2097 6994 2131
rect 6036 2043 6051 2063
rect 6051 2043 6070 2063
rect 6404 2059 6425 2063
rect 6425 2059 6438 2063
rect 6036 2029 6070 2043
rect 6404 2029 6438 2059
rect 6128 1965 6162 1995
rect 6128 1961 6157 1965
rect 6157 1961 6162 1965
rect 6588 1981 6622 1995
rect 6588 1961 6593 1981
rect 6593 1961 6622 1981
rect 6776 2029 6810 2063
rect 7052 2035 7084 2063
rect 7084 2035 7086 2063
rect 7052 2029 7086 2035
rect 6960 1961 6994 1995
rect 6226 1894 6260 1928
rect 7242 1912 7265 1922
rect 7265 1912 7276 1922
rect 7242 1886 7276 1912
rect 8222 2103 8256 2137
rect 8962 2103 8996 2137
rect 8038 2049 8053 2069
rect 8053 2049 8072 2069
rect 8406 2065 8427 2069
rect 8427 2065 8440 2069
rect 8038 2035 8072 2049
rect 8406 2035 8440 2065
rect 8130 1971 8164 2001
rect 8130 1967 8159 1971
rect 8159 1967 8164 1971
rect 8590 1987 8624 2001
rect 8590 1967 8595 1987
rect 8595 1967 8624 1987
rect 8778 2035 8812 2069
rect 9054 2041 9086 2069
rect 9086 2041 9088 2069
rect 9054 2035 9088 2041
rect 8962 1967 8996 2001
rect 8228 1900 8262 1934
rect 9244 1918 9267 1928
rect 9267 1918 9278 1928
rect 9244 1892 9278 1918
rect 10174 2103 10208 2137
rect 10914 2103 10948 2137
rect 9990 2049 10005 2069
rect 10005 2049 10024 2069
rect 10358 2065 10379 2069
rect 10379 2065 10392 2069
rect 9990 2035 10024 2049
rect 10358 2035 10392 2065
rect 10082 1971 10116 2001
rect 10082 1967 10111 1971
rect 10111 1967 10116 1971
rect 10542 1987 10576 2001
rect 10542 1967 10547 1987
rect 10547 1967 10576 1987
rect 10730 2035 10764 2069
rect 11006 2041 11038 2069
rect 11038 2041 11040 2069
rect 11006 2035 11040 2041
rect 10914 1967 10948 2001
rect 10180 1900 10214 1934
rect 11196 1918 11219 1928
rect 11219 1918 11230 1928
rect 11196 1892 11230 1918
rect 12166 2103 12200 2137
rect 12906 2103 12940 2137
rect 11982 2049 11997 2069
rect 11997 2049 12016 2069
rect 12350 2065 12371 2069
rect 12371 2065 12384 2069
rect 11982 2035 12016 2049
rect 12350 2035 12384 2065
rect 12074 1971 12108 2001
rect 12074 1967 12103 1971
rect 12103 1967 12108 1971
rect 12534 1987 12568 2001
rect 12534 1967 12539 1987
rect 12539 1967 12568 1987
rect 12722 2035 12756 2069
rect 12998 2041 13030 2069
rect 13030 2041 13032 2069
rect 12998 2035 13032 2041
rect 12906 1967 12940 2001
rect 12172 1900 12206 1934
rect 13188 1918 13211 1928
rect 13211 1918 13222 1928
rect 13188 1892 13222 1918
rect 14118 2103 14152 2137
rect 14858 2103 14892 2137
rect 13934 2049 13949 2069
rect 13949 2049 13968 2069
rect 14302 2065 14323 2069
rect 14323 2065 14336 2069
rect 13934 2035 13968 2049
rect 14302 2035 14336 2065
rect 14026 1971 14060 2001
rect 14026 1967 14055 1971
rect 14055 1967 14060 1971
rect 14486 1987 14520 2001
rect 14486 1967 14491 1987
rect 14491 1967 14520 1987
rect 14674 2035 14708 2069
rect 14950 2041 14982 2069
rect 14982 2041 14984 2069
rect 14950 2035 14984 2041
rect 14858 1967 14892 2001
rect 14124 1900 14158 1934
rect 15140 1918 15163 1928
rect 15163 1918 15174 1928
rect 15140 1892 15174 1918
rect 16182 2103 16216 2137
rect 16922 2103 16956 2137
rect 15998 2049 16013 2069
rect 16013 2049 16032 2069
rect 16366 2065 16387 2069
rect 16387 2065 16400 2069
rect 15998 2035 16032 2049
rect 16366 2035 16400 2065
rect 16090 1971 16124 2001
rect 16090 1967 16119 1971
rect 16119 1967 16124 1971
rect 16550 1987 16584 2001
rect 16550 1967 16555 1987
rect 16555 1967 16584 1987
rect 16738 2035 16772 2069
rect 17014 2041 17046 2069
rect 17046 2041 17048 2069
rect 17014 2035 17048 2041
rect 16922 1967 16956 2001
rect 16188 1900 16222 1934
rect 17204 1918 17227 1928
rect 17227 1918 17238 1928
rect 17204 1892 17238 1918
rect 3905 1723 3939 1757
rect 3997 1723 4031 1757
rect 4089 1723 4123 1757
rect 4181 1723 4215 1757
rect 4273 1723 4307 1757
rect 4365 1723 4399 1757
rect 4457 1723 4491 1757
rect 4549 1723 4583 1757
rect 4641 1723 4675 1757
rect 4733 1723 4767 1757
rect 4825 1723 4859 1757
rect 4917 1723 4951 1757
rect 5009 1723 5043 1757
rect 5101 1723 5135 1757
rect 5193 1723 5227 1757
rect 5285 1723 5319 1757
rect 5857 1723 5891 1757
rect 5949 1723 5983 1757
rect 6041 1723 6075 1757
rect 6133 1723 6167 1757
rect 6225 1723 6259 1757
rect 6317 1723 6351 1757
rect 6409 1723 6443 1757
rect 6501 1723 6535 1757
rect 6593 1723 6627 1757
rect 6685 1723 6719 1757
rect 6777 1723 6811 1757
rect 6869 1723 6903 1757
rect 6961 1723 6995 1757
rect 7053 1723 7087 1757
rect 7145 1723 7179 1757
rect 7237 1723 7271 1757
rect 7859 1729 7893 1763
rect 7951 1729 7985 1763
rect 8043 1729 8077 1763
rect 8135 1729 8169 1763
rect 8227 1729 8261 1763
rect 8319 1729 8353 1763
rect 8411 1729 8445 1763
rect 8503 1729 8537 1763
rect 8595 1729 8629 1763
rect 8687 1729 8721 1763
rect 8779 1729 8813 1763
rect 8871 1729 8905 1763
rect 8963 1729 8997 1763
rect 9055 1729 9089 1763
rect 9147 1729 9181 1763
rect 9239 1729 9273 1763
rect 9811 1729 9845 1763
rect 9903 1729 9937 1763
rect 9995 1729 10029 1763
rect 10087 1729 10121 1763
rect 10179 1729 10213 1763
rect 10271 1729 10305 1763
rect 10363 1729 10397 1763
rect 10455 1729 10489 1763
rect 10547 1729 10581 1763
rect 10639 1729 10673 1763
rect 10731 1729 10765 1763
rect 10823 1729 10857 1763
rect 10915 1729 10949 1763
rect 11007 1729 11041 1763
rect 11099 1729 11133 1763
rect 11191 1729 11225 1763
rect 11803 1729 11837 1763
rect 11895 1729 11929 1763
rect 11987 1729 12021 1763
rect 12079 1729 12113 1763
rect 12171 1729 12205 1763
rect 12263 1729 12297 1763
rect 12355 1729 12389 1763
rect 12447 1729 12481 1763
rect 12539 1729 12573 1763
rect 12631 1729 12665 1763
rect 12723 1729 12757 1763
rect 12815 1729 12849 1763
rect 12907 1729 12941 1763
rect 12999 1729 13033 1763
rect 13091 1729 13125 1763
rect 13183 1729 13217 1763
rect 13755 1729 13789 1763
rect 13847 1729 13881 1763
rect 13939 1729 13973 1763
rect 14031 1729 14065 1763
rect 14123 1729 14157 1763
rect 14215 1729 14249 1763
rect 14307 1729 14341 1763
rect 14399 1729 14433 1763
rect 14491 1729 14525 1763
rect 14583 1729 14617 1763
rect 14675 1729 14709 1763
rect 14767 1729 14801 1763
rect 14859 1729 14893 1763
rect 14951 1729 14985 1763
rect 15043 1729 15077 1763
rect 15135 1729 15169 1763
rect 15819 1729 15853 1763
rect 15911 1729 15945 1763
rect 16003 1729 16037 1763
rect 16095 1729 16129 1763
rect 16187 1729 16221 1763
rect 16279 1729 16313 1763
rect 16371 1729 16405 1763
rect 16463 1729 16497 1763
rect 16555 1729 16589 1763
rect 16647 1729 16681 1763
rect 16739 1729 16773 1763
rect 16831 1729 16865 1763
rect 16923 1729 16957 1763
rect 17015 1729 17049 1763
rect 17107 1729 17141 1763
rect 17199 1729 17233 1763
<< metal1 >>
rect 6603 17576 9539 17587
rect 6603 17504 6646 17576
rect 6722 17568 9539 17576
rect 6722 17532 9496 17568
rect 9532 17532 9539 17568
rect 6722 17504 9539 17532
rect 6603 17497 9539 17504
rect 9573 17572 13733 17587
rect 9573 17536 9596 17572
rect 9632 17536 13733 17572
rect 9573 17497 13733 17536
rect 9045 17054 11482 17055
rect 9036 17042 11482 17054
rect 9036 17041 11414 17042
rect 8787 16986 11414 17041
rect 11474 16986 11482 17042
rect 8787 16977 11482 16986
rect 8787 16964 9497 16977
rect 8787 16963 9000 16964
rect 9160 16963 9497 16964
rect 6578 15408 6682 15424
rect 6578 15356 6608 15408
rect 6660 15356 6682 15408
rect 6578 15342 6682 15356
rect 8787 14096 8865 16963
rect 9334 16628 9978 16638
rect 9334 16607 9456 16628
rect 9508 16607 9978 16628
rect 9334 16573 9363 16607
rect 9397 16573 9455 16607
rect 9508 16574 9547 16607
rect 9489 16573 9547 16574
rect 9581 16573 9639 16607
rect 9673 16573 9731 16607
rect 9765 16573 9823 16607
rect 9857 16573 9915 16607
rect 9949 16573 9978 16607
rect 9334 16542 9978 16573
rect 9412 16296 9472 16542
rect 10812 16410 11014 16442
rect 10812 16408 10872 16410
rect 9898 16394 10872 16408
rect 9898 16356 9910 16394
rect 9944 16356 10872 16394
rect 9898 16344 10872 16356
rect 10942 16408 11014 16410
rect 10942 16344 11125 16408
rect 9898 16342 11125 16344
rect 10812 16316 11014 16342
rect 9412 16262 9420 16296
rect 9454 16262 9472 16296
rect 9412 16242 9472 16262
rect 9502 16298 9612 16312
rect 9502 16264 9540 16298
rect 9574 16264 9612 16298
rect 9502 16256 9612 16264
rect 9536 16094 9567 16256
rect 9334 16078 9978 16094
rect 9334 16063 9842 16078
rect 9900 16063 9978 16078
rect 9334 16029 9363 16063
rect 9397 16029 9455 16063
rect 9489 16029 9547 16063
rect 9581 16029 9639 16063
rect 9673 16029 9731 16063
rect 9765 16029 9823 16063
rect 9900 16029 9915 16063
rect 9949 16029 9978 16063
rect 9334 16024 9842 16029
rect 9900 16024 9978 16029
rect 9334 15998 9978 16024
rect 9432 15878 9892 15894
rect 9432 15863 9612 15878
rect 9674 15863 9892 15878
rect 9432 15829 9461 15863
rect 9495 15829 9553 15863
rect 9587 15829 9612 15863
rect 9679 15829 9737 15863
rect 9771 15829 9829 15863
rect 9863 15829 9892 15863
rect 9432 15818 9612 15829
rect 9674 15818 9892 15829
rect 9432 15798 9892 15818
rect 9440 15574 9516 15590
rect 9642 15574 9696 15798
rect 11059 15637 11125 16342
rect 11474 15772 12118 15784
rect 11474 15753 11578 15772
rect 11646 15753 12118 15772
rect 11474 15719 11503 15753
rect 11537 15719 11578 15753
rect 11646 15719 11687 15753
rect 11721 15719 11779 15753
rect 11813 15719 11871 15753
rect 11905 15719 11963 15753
rect 11997 15719 12055 15753
rect 12089 15719 12118 15753
rect 11474 15710 11578 15719
rect 11646 15710 12118 15719
rect 11474 15688 12118 15710
rect 9440 15534 9454 15574
rect 9496 15534 9516 15574
rect 9440 15518 9516 15534
rect 9632 15564 9700 15574
rect 11059 15571 11913 15637
rect 11657 15568 11723 15571
rect 9632 15524 9644 15564
rect 9686 15524 9700 15564
rect 9450 15350 9504 15518
rect 9632 15512 9700 15524
rect 9824 15506 9910 15514
rect 9824 15494 9842 15506
rect 9824 15460 9836 15494
rect 9824 15452 9842 15460
rect 9896 15452 9910 15506
rect 9824 15440 9910 15452
rect 10060 15462 11722 15520
rect 10060 15456 11723 15462
rect 9632 15350 9700 15352
rect 9432 15336 9892 15350
rect 9432 15319 9764 15336
rect 9832 15319 9892 15336
rect 9432 15285 9461 15319
rect 9495 15285 9553 15319
rect 9587 15285 9645 15319
rect 9679 15285 9737 15319
rect 9863 15285 9892 15319
rect 9432 15274 9764 15285
rect 9832 15274 9892 15285
rect 9432 15254 9892 15274
rect 9344 15056 9988 15074
rect 9344 15043 9448 15056
rect 9514 15043 9988 15056
rect 9344 15009 9373 15043
rect 9407 15009 9448 15043
rect 9514 15009 9557 15043
rect 9591 15009 9649 15043
rect 9683 15009 9741 15043
rect 9775 15009 9833 15043
rect 9867 15009 9925 15043
rect 9959 15009 9988 15043
rect 9344 14990 9448 15009
rect 9514 14990 9988 15009
rect 9344 14978 9988 14990
rect 9422 14732 9482 14978
rect 10060 14946 10124 15456
rect 11657 15438 11723 15456
rect 11444 15412 11548 15428
rect 11444 15360 11474 15412
rect 11526 15404 11548 15412
rect 11534 15368 11548 15404
rect 11657 15402 11670 15438
rect 11704 15402 11723 15438
rect 11657 15394 11723 15402
rect 11526 15360 11548 15368
rect 11444 15346 11548 15360
rect 11847 15384 11913 15571
rect 12044 15444 12100 15448
rect 12044 15436 12266 15444
rect 12044 15402 12056 15436
rect 12090 15402 12266 15436
rect 12044 15394 12266 15402
rect 12044 15390 12100 15394
rect 11847 15348 11864 15384
rect 11898 15348 11913 15384
rect 11756 15318 11814 15334
rect 11214 15314 11814 15318
rect 10616 15268 11076 15284
rect 11214 15280 11768 15314
rect 11802 15280 11814 15314
rect 11214 15274 11814 15280
rect 10616 15253 10996 15268
rect 10616 15219 10645 15253
rect 10679 15219 10737 15253
rect 10771 15219 10829 15253
rect 10863 15219 10921 15253
rect 10955 15219 10996 15253
rect 10616 15206 10996 15219
rect 11064 15206 11076 15268
rect 10616 15188 11076 15206
rect 11216 15160 11296 15274
rect 11756 15268 11814 15274
rect 11847 15270 11913 15348
rect 10970 15152 11296 15160
rect 9906 14934 10124 14946
rect 9906 14900 9922 14934
rect 9956 14900 10124 14934
rect 9906 14882 10124 14900
rect 10156 15084 10886 15136
rect 10970 15116 11010 15152
rect 11050 15116 11296 15152
rect 11474 15222 12118 15240
rect 11474 15209 11980 15222
rect 12048 15209 12118 15222
rect 11474 15175 11503 15209
rect 11537 15175 11595 15209
rect 11629 15175 11687 15209
rect 11721 15175 11779 15209
rect 11813 15175 11871 15209
rect 11905 15175 11963 15209
rect 12048 15175 12055 15209
rect 12089 15175 12118 15209
rect 11474 15160 11980 15175
rect 12048 15160 12118 15175
rect 11474 15144 12118 15160
rect 10970 15102 11296 15116
rect 9422 14698 9430 14732
rect 9464 14698 9482 14732
rect 9422 14678 9482 14698
rect 9512 14734 9622 14748
rect 9512 14700 9550 14734
rect 9584 14700 9622 14734
rect 9512 14692 9622 14700
rect 9546 14530 9577 14692
rect 9344 14512 9988 14530
rect 9344 14499 9878 14512
rect 9944 14499 9988 14512
rect 9344 14465 9373 14499
rect 9407 14465 9465 14499
rect 9499 14465 9557 14499
rect 9591 14465 9649 14499
rect 9683 14465 9741 14499
rect 9775 14465 9833 14499
rect 9867 14465 9878 14499
rect 9959 14465 9988 14499
rect 9344 14446 9878 14465
rect 9944 14446 9988 14465
rect 9344 14434 9988 14446
rect 9442 14318 9902 14330
rect 9442 14299 9548 14318
rect 9620 14299 9902 14318
rect 9442 14265 9471 14299
rect 9505 14265 9548 14299
rect 9620 14265 9655 14299
rect 9689 14265 9747 14299
rect 9781 14265 9839 14299
rect 9873 14265 9902 14299
rect 9442 14248 9548 14265
rect 9620 14248 9902 14265
rect 9442 14234 9902 14248
rect 8182 14076 8865 14096
rect 8182 14036 8212 14076
rect 8254 14036 8865 14076
rect 8182 14018 8865 14036
rect 8602 13990 8638 14018
rect 9450 14010 9526 14028
rect 9654 14010 9700 14234
rect 7636 13974 7742 13976
rect 7636 13938 7806 13974
rect 9450 13970 9464 14010
rect 9506 13970 9526 14010
rect 9450 13954 9526 13970
rect 9642 14000 9710 14010
rect 9642 13960 9654 14000
rect 9696 13960 9710 14000
rect 7636 13936 7752 13938
rect 7636 13882 7652 13936
rect 7704 13904 7752 13936
rect 7792 13904 7806 13938
rect 7704 13882 7806 13904
rect 7636 13856 7806 13882
rect 9458 13786 9512 13954
rect 9642 13948 9710 13960
rect 9832 13904 10004 13918
rect 9832 13888 9896 13904
rect 9832 13854 9844 13888
rect 9880 13854 9896 13888
rect 9832 13842 9896 13854
rect 9956 13842 10004 13904
rect 9832 13824 10004 13842
rect 9442 13774 9902 13786
rect 9442 13755 9750 13774
rect 9822 13755 9902 13774
rect 7640 13738 7734 13754
rect 7640 13676 7656 13738
rect 7724 13676 7734 13738
rect 9442 13721 9471 13755
rect 9505 13721 9563 13755
rect 9597 13721 9655 13755
rect 9689 13721 9747 13755
rect 9822 13721 9839 13755
rect 9873 13721 9902 13755
rect 9442 13704 9750 13721
rect 9822 13704 9902 13721
rect 9442 13690 9902 13704
rect 7640 13656 7734 13676
rect 9336 13388 9980 13406
rect 9336 13375 9442 13388
rect 9514 13375 9980 13388
rect 9336 13341 9365 13375
rect 9399 13341 9442 13375
rect 9514 13341 9549 13375
rect 9583 13341 9641 13375
rect 9675 13341 9733 13375
rect 9767 13341 9825 13375
rect 9859 13341 9917 13375
rect 9951 13341 9980 13375
rect 9336 13322 9442 13341
rect 9514 13322 9980 13341
rect 9336 13310 9980 13322
rect 10156 13370 10208 15084
rect 10834 14960 10886 15084
rect 10636 14955 10772 14956
rect 10428 14942 10772 14955
rect 10428 14908 10690 14942
rect 10724 14908 10772 14942
rect 10428 14882 10772 14908
rect 10806 14942 10886 14960
rect 10806 14908 10830 14942
rect 10866 14908 10886 14942
rect 10806 14894 10886 14908
rect 10428 14877 10711 14882
rect 10428 13975 10506 14877
rect 10616 14720 11076 14740
rect 10616 14709 10660 14720
rect 10728 14709 11076 14720
rect 10616 14675 10645 14709
rect 10728 14675 10737 14709
rect 10771 14675 10829 14709
rect 10863 14675 10921 14709
rect 10955 14675 11013 14709
rect 11047 14675 11076 14709
rect 10616 14658 10660 14675
rect 10728 14658 11076 14675
rect 10616 14644 11076 14658
rect 10690 14298 11334 14318
rect 10690 14287 11216 14298
rect 11284 14287 11334 14298
rect 10690 14253 10719 14287
rect 10753 14253 10811 14287
rect 10845 14253 10903 14287
rect 10937 14253 10995 14287
rect 11029 14253 11087 14287
rect 11121 14253 11179 14287
rect 11213 14253 11216 14287
rect 11305 14253 11334 14287
rect 10690 14236 11216 14253
rect 11284 14236 11334 14253
rect 10690 14222 11334 14236
rect 12213 14181 12263 15394
rect 13643 14697 13733 17497
rect 16187 16853 18657 16863
rect 16187 16847 20570 16853
rect 16187 16833 23479 16847
rect 16187 16367 16217 16833
rect 18512 16823 23479 16833
rect 19995 16817 23479 16823
rect 21207 16806 21237 16817
rect 16400 16400 16466 16420
rect 16400 16367 16416 16400
rect 16187 16366 16416 16367
rect 16452 16366 16466 16400
rect 16187 16337 16466 16366
rect 16496 16392 17234 16412
rect 16496 16388 17184 16392
rect 16496 16354 16502 16388
rect 16540 16358 17184 16388
rect 17222 16358 17234 16392
rect 16540 16354 17234 16358
rect 16496 16338 17234 16354
rect 17264 16396 18106 16418
rect 17264 16384 18048 16396
rect 17264 16350 17278 16384
rect 17312 16362 18048 16384
rect 18082 16362 18106 16396
rect 17312 16350 18106 16362
rect 16400 16336 16466 16337
rect 17264 16328 18106 16350
rect 18138 16392 18200 16416
rect 18138 16358 18150 16392
rect 18186 16390 18200 16392
rect 18656 16390 18722 16410
rect 18186 16388 18314 16390
rect 18656 16388 18672 16390
rect 18186 16358 18672 16388
rect 18138 16356 18672 16358
rect 18708 16356 18722 16390
rect 18138 16348 18722 16356
rect 18194 16342 18722 16348
rect 18512 16327 18722 16342
rect 18752 16382 19490 16402
rect 18752 16378 19440 16382
rect 18752 16344 18758 16378
rect 18796 16348 19440 16378
rect 19478 16348 19490 16382
rect 18796 16344 19490 16348
rect 18752 16328 19490 16344
rect 19520 16386 20362 16408
rect 19520 16374 20304 16386
rect 19520 16340 19534 16374
rect 19568 16352 20304 16374
rect 20338 16352 20362 16386
rect 19568 16340 20362 16352
rect 18656 16326 18722 16327
rect 19520 16318 20362 16340
rect 20394 16392 20456 16406
rect 21418 16392 21486 16404
rect 20394 16384 21486 16392
rect 20394 16382 21436 16384
rect 20394 16348 20406 16382
rect 20442 16350 21436 16382
rect 21472 16350 21486 16384
rect 20442 16348 21486 16350
rect 20394 16338 21486 16348
rect 20440 16336 21486 16338
rect 21418 16320 21486 16336
rect 21516 16376 22254 16396
rect 21516 16372 22204 16376
rect 21516 16338 21522 16372
rect 21560 16342 22204 16372
rect 22242 16342 22254 16376
rect 21560 16338 22254 16342
rect 21516 16322 22254 16338
rect 22284 16380 23126 16402
rect 22284 16368 23068 16380
rect 22284 16334 22298 16368
rect 22332 16346 23068 16368
rect 23102 16346 23126 16380
rect 22332 16334 23126 16346
rect 22284 16312 23126 16334
rect 23158 16376 23220 16400
rect 23158 16342 23170 16376
rect 23206 16374 23220 16376
rect 23449 16374 23479 16817
rect 23206 16344 23479 16374
rect 23206 16342 23220 16344
rect 23158 16332 23220 16342
rect 21575 16086 21605 16182
rect 23373 15607 23403 16344
rect 23372 15606 23403 15607
rect 22975 15577 23403 15606
rect 22975 14749 23005 15577
rect 22975 14719 23731 14749
rect 13643 14607 22797 14697
rect 23701 14614 23731 14719
rect 24138 14714 24198 14726
rect 24138 14662 24144 14714
rect 24196 14662 24198 14714
rect 24138 14650 24198 14662
rect 24138 14616 24150 14650
rect 24186 14616 24198 14650
rect 12588 14288 13140 14302
rect 12588 14271 12782 14288
rect 12850 14271 13140 14288
rect 12588 14237 12617 14271
rect 12651 14237 12709 14271
rect 12743 14237 12782 14271
rect 12850 14237 12893 14271
rect 12927 14237 12985 14271
rect 13019 14237 13077 14271
rect 13111 14237 13140 14271
rect 12588 14226 12782 14237
rect 12850 14226 13140 14237
rect 12588 14206 13140 14226
rect 13643 14182 13733 14607
rect 22618 14599 22797 14607
rect 22618 14580 23581 14599
rect 22618 14546 23530 14580
rect 23568 14546 23581 14580
rect 22618 14509 23581 14546
rect 23644 14562 23732 14614
rect 24138 14578 24198 14616
rect 23644 14528 23672 14562
rect 23708 14528 23732 14562
rect 22618 14508 22736 14509
rect 23644 14490 23732 14528
rect 24444 14564 24510 14620
rect 24444 14512 24452 14564
rect 24504 14512 24510 14564
rect 24444 14502 24510 14512
rect 24550 14588 24604 14620
rect 24550 14578 24556 14588
rect 24592 14578 24604 14588
rect 24550 14526 24552 14578
rect 24550 14502 24604 14526
rect 24684 14562 24770 14618
rect 24684 14536 24712 14562
rect 24746 14536 24770 14562
rect 25348 14598 28230 14610
rect 25348 14562 25364 14598
rect 25400 14562 28230 14598
rect 25348 14546 28230 14562
rect 24684 14484 24698 14536
rect 24750 14484 24770 14536
rect 24684 14434 24770 14484
rect 23850 14318 24212 14334
rect 23850 14258 23992 14318
rect 24054 14258 24212 14318
rect 23850 14240 24212 14258
rect 12213 14176 12264 14181
rect 12213 14170 12940 14176
rect 12213 14136 12762 14170
rect 12798 14136 12940 14170
rect 12213 14129 12940 14136
rect 12256 14128 12940 14129
rect 13470 14132 13733 14182
rect 13470 14100 13732 14132
rect 12312 14034 12980 14094
rect 10689 13980 10767 14033
rect 12312 14022 12386 14034
rect 10689 13975 10716 13980
rect 10428 13946 10716 13975
rect 10750 13946 10767 13980
rect 10428 13897 10767 13946
rect 10156 13360 10242 13370
rect 9414 13064 9474 13310
rect 10156 13308 10164 13360
rect 10226 13308 10242 13360
rect 10156 13300 10242 13308
rect 10156 13232 10208 13300
rect 9902 13224 10208 13232
rect 9902 13190 9914 13224
rect 9948 13190 10208 13224
rect 9902 13180 10208 13190
rect 10428 13089 10506 13897
rect 10868 13894 10938 13940
rect 10868 13842 10878 13894
rect 10930 13842 10938 13894
rect 10868 13802 10938 13842
rect 10966 13934 11034 13990
rect 10966 13882 10976 13934
rect 11028 13882 11034 13934
rect 10966 13804 11034 13882
rect 11068 13974 11140 13992
rect 11068 13936 11078 13974
rect 11114 13936 11140 13974
rect 11068 13890 11140 13936
rect 11068 13834 11074 13890
rect 11126 13834 11140 13890
rect 11660 13922 12120 13944
rect 11660 13913 11694 13922
rect 11762 13913 12120 13922
rect 11660 13879 11689 13913
rect 11762 13879 11781 13913
rect 11815 13879 11873 13913
rect 11907 13879 11965 13913
rect 11999 13879 12057 13913
rect 12091 13879 12120 13913
rect 11068 13808 11140 13834
rect 11246 13856 11532 13876
rect 11246 13818 11260 13856
rect 11298 13818 11532 13856
rect 11660 13860 11694 13879
rect 11762 13860 12120 13879
rect 11660 13848 12120 13860
rect 12312 13934 12384 14022
rect 12702 13984 12842 13996
rect 12502 13978 12608 13980
rect 12502 13942 12672 13978
rect 12502 13940 12618 13942
rect 11246 13802 11532 13818
rect 11451 13789 11532 13802
rect 12312 13790 12382 13934
rect 12502 13886 12518 13940
rect 12570 13908 12618 13940
rect 12658 13908 12672 13942
rect 12570 13886 12672 13908
rect 12702 13908 12732 13984
rect 12812 13962 12842 13984
rect 12908 13976 12980 14034
rect 13048 14080 13732 14100
rect 13048 14040 13078 14080
rect 13120 14040 13732 14080
rect 13048 14022 13732 14040
rect 13468 13996 13732 14022
rect 13468 13994 13504 13996
rect 12812 13908 12840 13962
rect 12886 13960 12980 13976
rect 12886 13924 12918 13960
rect 12956 13924 12980 13960
rect 12886 13908 12980 13924
rect 12702 13894 12840 13908
rect 12502 13860 12672 13886
rect 10690 13758 11334 13774
rect 10690 13743 10728 13758
rect 10796 13743 11334 13758
rect 10690 13709 10719 13743
rect 10796 13709 10811 13743
rect 10845 13709 10903 13743
rect 10937 13709 10995 13743
rect 11029 13709 11087 13743
rect 11121 13709 11179 13743
rect 11213 13709 11271 13743
rect 11305 13709 11334 13743
rect 11451 13715 11929 13789
rect 11986 13768 12382 13790
rect 11986 13734 12028 13768
rect 12062 13734 12382 13768
rect 11986 13718 12382 13734
rect 12506 13742 13140 13758
rect 10690 13696 10728 13709
rect 10796 13696 11334 13709
rect 10690 13678 11334 13696
rect 11855 13608 11929 13715
rect 12506 13680 12522 13742
rect 12590 13727 13140 13742
rect 12590 13693 12617 13727
rect 12651 13693 12709 13727
rect 12743 13693 12801 13727
rect 12835 13693 12893 13727
rect 12927 13693 12985 13727
rect 13019 13693 13077 13727
rect 13111 13693 13140 13727
rect 12590 13680 13140 13693
rect 12506 13662 13140 13680
rect 12506 13660 12600 13662
rect 11410 13558 11759 13581
rect 11410 13524 11700 13558
rect 11734 13524 11759 13558
rect 11410 13507 11759 13524
rect 11855 13574 11878 13608
rect 11912 13574 11929 13608
rect 10814 13454 11274 13476
rect 10814 13445 10850 13454
rect 10918 13445 11274 13454
rect 10814 13411 10843 13445
rect 10918 13411 10935 13445
rect 10969 13411 11027 13445
rect 11061 13411 11119 13445
rect 11153 13411 11211 13445
rect 11245 13411 11274 13445
rect 10814 13394 10850 13411
rect 10918 13394 11274 13411
rect 10814 13380 11274 13394
rect 10986 13342 11084 13348
rect 10986 13290 11006 13342
rect 11060 13290 11084 13342
rect 11410 13302 11484 13507
rect 11855 13493 11929 13574
rect 11660 13382 12120 13400
rect 11660 13369 12002 13382
rect 12070 13369 12120 13382
rect 11660 13335 11689 13369
rect 11723 13335 11781 13369
rect 11815 13335 11873 13369
rect 11907 13335 11965 13369
rect 11999 13335 12002 13369
rect 12091 13335 12120 13369
rect 11660 13320 12002 13335
rect 12070 13320 12120 13335
rect 11660 13304 12120 13320
rect 10986 13272 11084 13290
rect 11198 13282 11484 13302
rect 11198 13244 11208 13282
rect 11246 13244 11484 13282
rect 11198 13228 11484 13244
rect 9414 13030 9422 13064
rect 9456 13030 9474 13064
rect 9414 13010 9474 13030
rect 9504 13066 9614 13080
rect 9504 13032 9542 13066
rect 9576 13032 9614 13066
rect 9504 13024 9614 13032
rect 10428 13064 10947 13089
rect 10428 13030 10860 13064
rect 10894 13030 10947 13064
rect 9538 12862 9569 13024
rect 10428 13011 10947 13030
rect 11042 13086 11124 13158
rect 11042 13032 11062 13086
rect 11114 13032 11124 13086
rect 9336 12848 9980 12862
rect 9336 12831 9856 12848
rect 9928 12831 9980 12848
rect 9336 12797 9365 12831
rect 9399 12797 9457 12831
rect 9491 12797 9549 12831
rect 9583 12797 9641 12831
rect 9675 12797 9733 12831
rect 9767 12797 9825 12831
rect 9951 12797 9980 12831
rect 9336 12782 9856 12797
rect 9928 12782 9980 12797
rect 9336 12766 9980 12782
rect 9434 12646 9894 12662
rect 9434 12631 9500 12646
rect 9574 12631 9894 12646
rect 9434 12597 9463 12631
rect 9497 12597 9500 12631
rect 9589 12597 9647 12631
rect 9681 12597 9739 12631
rect 9773 12597 9831 12631
rect 9865 12597 9894 12631
rect 9434 12580 9500 12597
rect 9574 12580 9894 12597
rect 9434 12566 9894 12580
rect 9442 12342 9518 12368
rect 9642 12342 9692 12566
rect 9826 12394 9976 12408
rect 9826 12374 9872 12394
rect 9442 12302 9456 12342
rect 9498 12302 9518 12342
rect 9442 12286 9518 12302
rect 9634 12332 9702 12342
rect 9634 12292 9646 12332
rect 9688 12292 9702 12332
rect 9826 12340 9836 12374
rect 9826 12326 9872 12340
rect 9934 12326 9976 12394
rect 9826 12310 9976 12326
rect 9456 12118 9508 12286
rect 9634 12280 9702 12292
rect 10428 12125 10506 13011
rect 11042 12974 11124 13032
rect 10814 12920 11274 12932
rect 10814 12901 10862 12920
rect 10930 12901 11274 12920
rect 10814 12867 10843 12901
rect 10930 12867 10935 12901
rect 10969 12867 11027 12901
rect 11061 12867 11119 12901
rect 11153 12867 11211 12901
rect 11245 12867 11274 12901
rect 10814 12860 10862 12867
rect 10930 12860 11274 12867
rect 10814 12836 11274 12860
rect 10810 12436 11270 12456
rect 10810 12425 11146 12436
rect 11214 12425 11270 12436
rect 10810 12391 10839 12425
rect 10873 12391 10931 12425
rect 10965 12391 11023 12425
rect 11057 12391 11115 12425
rect 11241 12391 11270 12425
rect 10810 12374 11146 12391
rect 11214 12374 11270 12391
rect 10810 12360 11270 12374
rect 11200 12212 11268 12222
rect 11200 12160 11206 12212
rect 11258 12160 11268 12212
rect 11200 12154 11268 12160
rect 9434 12104 9894 12118
rect 9434 12087 9772 12104
rect 9846 12087 9894 12104
rect 9434 12053 9463 12087
rect 9497 12053 9555 12087
rect 9589 12053 9647 12087
rect 9681 12053 9739 12087
rect 9865 12053 9894 12087
rect 9434 12038 9772 12053
rect 9846 12038 9894 12053
rect 9434 12022 9894 12038
rect 10428 12116 10961 12125
rect 10428 12082 10884 12116
rect 10920 12082 10961 12116
rect 10428 12047 10961 12082
rect 11008 12122 11078 12130
rect 11008 12070 11016 12122
rect 11068 12070 11078 12122
rect 11008 12064 11078 12070
rect 9346 11824 9990 11842
rect 9346 11811 9426 11824
rect 9506 11811 9990 11824
rect 9346 11777 9375 11811
rect 9409 11777 9426 11811
rect 9506 11777 9559 11811
rect 9593 11777 9651 11811
rect 9685 11777 9743 11811
rect 9777 11777 9835 11811
rect 9869 11777 9927 11811
rect 9961 11777 9990 11811
rect 9346 11760 9426 11777
rect 9506 11760 9990 11777
rect 9346 11746 9990 11760
rect 9424 11500 9484 11746
rect 10428 11674 10506 12047
rect 10810 11896 11270 11912
rect 10810 11881 10868 11896
rect 10936 11881 11270 11896
rect 10810 11847 10839 11881
rect 10965 11847 11023 11881
rect 11057 11847 11115 11881
rect 11149 11847 11207 11881
rect 11241 11847 11270 11881
rect 10810 11834 10868 11847
rect 10936 11834 11270 11847
rect 10810 11816 11270 11834
rect 9908 11660 10506 11674
rect 9908 11626 9914 11660
rect 9950 11626 10506 11660
rect 9908 11596 10506 11626
rect 9424 11466 9432 11500
rect 9466 11466 9484 11500
rect 9424 11446 9484 11466
rect 9514 11502 9624 11516
rect 9514 11468 9552 11502
rect 9586 11468 9624 11502
rect 9514 11460 9624 11468
rect 9548 11298 9579 11460
rect 9346 11282 9990 11298
rect 9346 11267 9860 11282
rect 9940 11267 9990 11282
rect 9346 11233 9375 11267
rect 9409 11233 9467 11267
rect 9501 11233 9559 11267
rect 9593 11233 9651 11267
rect 9685 11233 9743 11267
rect 9777 11233 9835 11267
rect 9961 11233 9990 11267
rect 9346 11218 9860 11233
rect 9940 11218 9990 11233
rect 9346 11202 9990 11218
rect 9444 11078 9904 11098
rect 9444 11067 9492 11078
rect 9572 11067 9904 11078
rect 9444 11033 9473 11067
rect 9599 11033 9657 11067
rect 9691 11033 9749 11067
rect 9783 11033 9841 11067
rect 9875 11033 9904 11067
rect 9444 11014 9492 11033
rect 9572 11014 9904 11033
rect 9444 11002 9904 11014
rect 9452 10778 9528 10790
rect 4970 10732 5202 10762
rect 4970 10730 5054 10732
rect 4970 10694 4982 10730
rect 5016 10694 5054 10730
rect 4970 10676 5054 10694
rect 5108 10676 5202 10732
rect 9452 10738 9466 10778
rect 9508 10738 9528 10778
rect 9452 10722 9528 10738
rect 9642 10768 9714 11002
rect 9642 10734 9656 10768
rect 9644 10728 9656 10734
rect 9698 10734 9714 10768
rect 9836 10736 10068 10766
rect 9836 10734 9920 10736
rect 9698 10728 9712 10734
rect 4970 10652 5202 10676
rect 9472 10554 9522 10722
rect 9644 10712 9712 10728
rect 9836 10698 9848 10734
rect 9882 10698 9920 10734
rect 9836 10680 9920 10698
rect 9974 10680 10068 10736
rect 9836 10656 10068 10680
rect 9644 10554 9712 10558
rect 9444 10544 9904 10554
rect 9444 10523 9770 10544
rect 9850 10523 9904 10544
rect 9444 10489 9473 10523
rect 9507 10489 9565 10523
rect 9599 10489 9657 10523
rect 9691 10489 9749 10523
rect 9875 10489 9904 10523
rect 9444 10480 9770 10489
rect 9850 10480 9904 10489
rect 9444 10458 9904 10480
rect 6112 6638 6388 6648
rect 6112 6617 6226 6638
rect 6282 6617 6388 6638
rect 6112 6583 6141 6617
rect 6175 6583 6226 6617
rect 6282 6583 6325 6617
rect 6359 6583 6388 6617
rect 6112 6580 6226 6583
rect 6282 6580 6388 6583
rect 6112 6552 6388 6580
rect 6134 6390 6228 6398
rect 6134 6338 6168 6390
rect 6220 6338 6228 6390
rect 6262 6396 6328 6398
rect 6262 6344 6268 6396
rect 6320 6344 6328 6396
rect 6262 6338 6328 6344
rect 6134 6332 6228 6338
rect 6112 6088 6388 6104
rect 6112 6073 6170 6088
rect 6226 6073 6388 6088
rect 6112 6039 6141 6073
rect 6226 6039 6233 6073
rect 6267 6039 6325 6073
rect 6359 6039 6388 6073
rect 6112 6030 6170 6039
rect 6226 6030 6388 6039
rect 6112 6008 6388 6030
rect 10018 6002 11490 6016
rect 10018 5985 10406 6002
rect 10464 6000 11490 6002
rect 10464 5985 10774 6000
rect 10832 5985 11490 6000
rect 10018 5951 10047 5985
rect 10081 5951 10139 5985
rect 10173 5951 10231 5985
rect 10265 5951 10323 5985
rect 10357 5951 10406 5985
rect 10464 5951 10507 5985
rect 10541 5951 10599 5985
rect 10633 5951 10691 5985
rect 10725 5951 10774 5985
rect 10832 5951 10875 5985
rect 10909 5951 10967 5985
rect 11001 5951 11059 5985
rect 11093 5951 11151 5985
rect 11185 5951 11243 5985
rect 11277 5951 11335 5985
rect 11369 5951 11427 5985
rect 11461 5951 11490 5985
rect 10018 5940 10406 5951
rect 10464 5940 10774 5951
rect 10018 5936 10774 5940
rect 10832 5936 11490 5951
rect 10018 5920 11490 5936
rect 12080 5986 13552 6004
rect 12080 5973 12796 5986
rect 12852 5973 13552 5986
rect 12080 5939 12109 5973
rect 12143 5939 12201 5973
rect 12235 5939 12293 5973
rect 12327 5939 12385 5973
rect 12419 5939 12477 5973
rect 12511 5939 12569 5973
rect 12603 5939 12661 5973
rect 12695 5939 12753 5973
rect 12787 5939 12796 5973
rect 12879 5939 12937 5973
rect 12971 5939 13029 5973
rect 13063 5939 13121 5973
rect 13155 5939 13213 5973
rect 13247 5939 13305 5973
rect 13339 5939 13397 5973
rect 13431 5939 13489 5973
rect 13523 5939 13552 5973
rect 12080 5928 12796 5939
rect 12852 5928 13552 5939
rect 10214 5747 10272 5753
rect 10214 5713 10226 5747
rect 10260 5744 10272 5747
rect 10300 5744 10328 5920
rect 12080 5908 13552 5928
rect 14038 5994 15510 6012
rect 14038 5981 14754 5994
rect 14810 5981 15510 5994
rect 14038 5947 14067 5981
rect 14101 5947 14159 5981
rect 14193 5947 14251 5981
rect 14285 5947 14343 5981
rect 14377 5947 14435 5981
rect 14469 5947 14527 5981
rect 14561 5947 14619 5981
rect 14653 5947 14711 5981
rect 14745 5947 14754 5981
rect 14837 5947 14895 5981
rect 14929 5947 14987 5981
rect 15021 5947 15079 5981
rect 15113 5947 15171 5981
rect 15205 5947 15263 5981
rect 15297 5947 15355 5981
rect 15389 5947 15447 5981
rect 15481 5947 15510 5981
rect 14038 5936 14754 5947
rect 14810 5936 15510 5947
rect 14038 5916 15510 5936
rect 16032 6000 17504 6018
rect 16032 5987 16748 6000
rect 16804 5987 17504 6000
rect 16032 5953 16061 5987
rect 16095 5953 16153 5987
rect 16187 5953 16245 5987
rect 16279 5953 16337 5987
rect 16371 5953 16429 5987
rect 16463 5953 16521 5987
rect 16555 5953 16613 5987
rect 16647 5953 16705 5987
rect 16739 5953 16748 5987
rect 16831 5953 16889 5987
rect 16923 5953 16981 5987
rect 17015 5953 17073 5987
rect 17107 5953 17165 5987
rect 17199 5953 17257 5987
rect 17291 5953 17349 5987
rect 17383 5953 17441 5987
rect 17475 5953 17504 5987
rect 16032 5942 16748 5953
rect 16804 5942 17504 5953
rect 16032 5922 17504 5942
rect 10398 5815 10456 5821
rect 10398 5781 10410 5815
rect 10444 5812 10456 5815
rect 11138 5815 11196 5821
rect 11138 5812 11150 5815
rect 10444 5784 11150 5812
rect 10444 5781 10456 5784
rect 10398 5775 10456 5781
rect 11138 5781 11150 5784
rect 11184 5781 11196 5815
rect 11138 5775 11196 5781
rect 10582 5747 10640 5753
rect 10582 5744 10594 5747
rect 10260 5716 10594 5744
rect 10260 5713 10272 5716
rect 10214 5707 10272 5713
rect 10582 5713 10594 5716
rect 10628 5744 10640 5747
rect 10954 5747 11012 5753
rect 10954 5744 10966 5747
rect 10628 5716 10966 5744
rect 10628 5713 10640 5716
rect 10582 5707 10640 5713
rect 10954 5713 10966 5716
rect 11000 5744 11012 5747
rect 11230 5747 11288 5753
rect 11230 5744 11242 5747
rect 11000 5716 11242 5744
rect 11000 5713 11012 5716
rect 10954 5707 11012 5713
rect 11230 5713 11242 5716
rect 11276 5713 11288 5747
rect 11230 5707 11288 5713
rect 12276 5735 12334 5741
rect 12276 5701 12288 5735
rect 12322 5732 12334 5735
rect 12362 5732 12390 5908
rect 12460 5803 12518 5809
rect 12460 5769 12472 5803
rect 12506 5800 12518 5803
rect 13200 5803 13258 5809
rect 13200 5800 13212 5803
rect 12506 5772 13212 5800
rect 12506 5769 12518 5772
rect 12460 5763 12518 5769
rect 13200 5769 13212 5772
rect 13246 5769 13258 5803
rect 13200 5763 13258 5769
rect 14234 5743 14292 5749
rect 12644 5735 12702 5741
rect 12644 5732 12656 5735
rect 12322 5704 12656 5732
rect 12322 5701 12334 5704
rect 12276 5695 12334 5701
rect 12644 5701 12656 5704
rect 12690 5732 12702 5735
rect 13016 5735 13074 5741
rect 13016 5732 13028 5735
rect 12690 5704 13028 5732
rect 12690 5701 12702 5704
rect 12644 5695 12702 5701
rect 13016 5701 13028 5704
rect 13062 5732 13074 5735
rect 13292 5735 13350 5741
rect 13292 5732 13304 5735
rect 13062 5704 13304 5732
rect 13062 5701 13074 5704
rect 13016 5695 13074 5701
rect 13292 5701 13304 5704
rect 13338 5701 13350 5735
rect 14234 5709 14246 5743
rect 14280 5740 14292 5743
rect 14320 5740 14348 5916
rect 14418 5811 14476 5817
rect 14418 5777 14430 5811
rect 14464 5808 14476 5811
rect 15158 5811 15216 5817
rect 15158 5808 15170 5811
rect 14464 5780 15170 5808
rect 14464 5777 14476 5780
rect 14418 5771 14476 5777
rect 15158 5777 15170 5780
rect 15204 5777 15216 5811
rect 15158 5771 15216 5777
rect 16228 5749 16286 5755
rect 14602 5743 14660 5749
rect 14602 5740 14614 5743
rect 14280 5712 14614 5740
rect 14280 5709 14292 5712
rect 14234 5703 14292 5709
rect 14602 5709 14614 5712
rect 14648 5740 14660 5743
rect 14974 5743 15032 5749
rect 14974 5740 14986 5743
rect 14648 5712 14986 5740
rect 14648 5709 14660 5712
rect 14602 5703 14660 5709
rect 14974 5709 14986 5712
rect 15020 5740 15032 5743
rect 15250 5743 15308 5749
rect 15250 5740 15262 5743
rect 15020 5712 15262 5740
rect 15020 5709 15032 5712
rect 14974 5703 15032 5709
rect 15250 5709 15262 5712
rect 15296 5709 15308 5743
rect 16228 5715 16240 5749
rect 16274 5746 16286 5749
rect 16314 5746 16342 5922
rect 16412 5817 16470 5823
rect 16412 5783 16424 5817
rect 16458 5814 16470 5817
rect 17152 5817 17210 5823
rect 17152 5814 17164 5817
rect 16458 5786 17164 5814
rect 16458 5783 16470 5786
rect 16412 5777 16470 5783
rect 17152 5783 17164 5786
rect 17198 5783 17210 5817
rect 17152 5777 17210 5783
rect 28166 5774 28230 14546
rect 16596 5749 16654 5755
rect 16596 5746 16608 5749
rect 16274 5718 16608 5746
rect 16274 5715 16286 5718
rect 16228 5709 16286 5715
rect 16596 5715 16608 5718
rect 16642 5746 16654 5749
rect 16968 5749 17026 5755
rect 16968 5746 16980 5749
rect 16642 5718 16980 5746
rect 16642 5715 16654 5718
rect 16596 5709 16654 5715
rect 16968 5715 16980 5718
rect 17014 5746 17026 5749
rect 17244 5749 17302 5755
rect 17244 5746 17256 5749
rect 17014 5718 17256 5746
rect 17014 5715 17026 5718
rect 16968 5709 17026 5715
rect 17244 5715 17256 5718
rect 17290 5715 17302 5749
rect 17244 5709 17302 5715
rect 28166 5710 30432 5774
rect 15250 5703 15308 5709
rect 13292 5695 13350 5701
rect 10306 5679 10364 5685
rect 10306 5645 10318 5679
rect 10352 5676 10364 5679
rect 10766 5679 10824 5685
rect 10766 5676 10778 5679
rect 10352 5648 10778 5676
rect 10352 5645 10364 5648
rect 10306 5639 10364 5645
rect 10766 5645 10778 5648
rect 10812 5676 10824 5679
rect 11138 5679 11196 5685
rect 16320 5681 16378 5687
rect 11138 5676 11150 5679
rect 10812 5648 11150 5676
rect 10812 5645 10824 5648
rect 10766 5639 10824 5645
rect 10404 5618 10470 5620
rect 1836 5578 3308 5596
rect 1836 5565 2564 5578
rect 2620 5565 3308 5578
rect 1836 5531 1865 5565
rect 1899 5531 1957 5565
rect 1991 5531 2049 5565
rect 2083 5531 2141 5565
rect 2175 5531 2233 5565
rect 2267 5531 2325 5565
rect 2359 5531 2417 5565
rect 2451 5531 2509 5565
rect 2543 5531 2564 5565
rect 2635 5531 2693 5565
rect 2727 5531 2785 5565
rect 2819 5531 2877 5565
rect 2911 5531 2969 5565
rect 3003 5531 3061 5565
rect 3095 5531 3153 5565
rect 3187 5531 3245 5565
rect 3279 5531 3308 5565
rect 1836 5520 2564 5531
rect 2620 5520 3308 5531
rect 1836 5500 3308 5520
rect 3970 5570 5442 5588
rect 3970 5557 4686 5570
rect 4742 5557 5442 5570
rect 3970 5523 3999 5557
rect 4033 5523 4091 5557
rect 4125 5523 4183 5557
rect 4217 5523 4275 5557
rect 4309 5523 4367 5557
rect 4401 5523 4459 5557
rect 4493 5523 4551 5557
rect 4585 5523 4643 5557
rect 4677 5523 4686 5557
rect 4769 5523 4827 5557
rect 4861 5523 4919 5557
rect 4953 5523 5011 5557
rect 5045 5523 5103 5557
rect 5137 5523 5195 5557
rect 5229 5523 5287 5557
rect 5321 5523 5379 5557
rect 5413 5523 5442 5557
rect 3970 5512 4686 5523
rect 4742 5512 5442 5523
rect 2032 5327 2090 5333
rect 2032 5293 2044 5327
rect 2078 5324 2090 5327
rect 2118 5324 2146 5500
rect 3970 5492 5442 5512
rect 5922 5570 7394 5588
rect 5922 5557 6638 5570
rect 6694 5557 7394 5570
rect 5922 5523 5951 5557
rect 5985 5523 6043 5557
rect 6077 5523 6135 5557
rect 6169 5523 6227 5557
rect 6261 5523 6319 5557
rect 6353 5523 6411 5557
rect 6445 5523 6503 5557
rect 6537 5523 6595 5557
rect 6629 5523 6638 5557
rect 6721 5523 6779 5557
rect 6813 5523 6871 5557
rect 6905 5523 6963 5557
rect 6997 5523 7055 5557
rect 7089 5523 7147 5557
rect 7181 5523 7239 5557
rect 7273 5523 7331 5557
rect 7365 5523 7394 5557
rect 5922 5512 6638 5523
rect 6694 5512 7394 5523
rect 5922 5492 7394 5512
rect 7924 5576 9396 5594
rect 7924 5563 8640 5576
rect 8696 5563 9396 5576
rect 7924 5529 7953 5563
rect 7987 5529 8045 5563
rect 8079 5529 8137 5563
rect 8171 5529 8229 5563
rect 8263 5529 8321 5563
rect 8355 5529 8413 5563
rect 8447 5529 8505 5563
rect 8539 5529 8597 5563
rect 8631 5529 8640 5563
rect 8723 5529 8781 5563
rect 8815 5529 8873 5563
rect 8907 5529 8965 5563
rect 8999 5529 9057 5563
rect 9091 5529 9149 5563
rect 9183 5529 9241 5563
rect 9275 5529 9333 5563
rect 9367 5529 9396 5563
rect 10404 5566 10410 5618
rect 10462 5566 10470 5618
rect 10404 5562 10470 5566
rect 7924 5518 8640 5529
rect 8696 5518 9396 5529
rect 7924 5498 9396 5518
rect 2216 5395 2274 5401
rect 2216 5361 2228 5395
rect 2262 5392 2274 5395
rect 2956 5395 3014 5401
rect 2956 5392 2968 5395
rect 2262 5364 2968 5392
rect 2262 5361 2274 5364
rect 2216 5355 2274 5361
rect 2956 5361 2968 5364
rect 3002 5361 3014 5395
rect 2956 5355 3014 5361
rect 2400 5327 2458 5333
rect 2400 5324 2412 5327
rect 2078 5296 2412 5324
rect 2078 5293 2090 5296
rect 2032 5287 2090 5293
rect 2400 5293 2412 5296
rect 2446 5324 2458 5327
rect 2772 5327 2830 5333
rect 2772 5324 2784 5327
rect 2446 5296 2784 5324
rect 2446 5293 2458 5296
rect 2400 5287 2458 5293
rect 2772 5293 2784 5296
rect 2818 5324 2830 5327
rect 3048 5327 3106 5333
rect 3048 5324 3060 5327
rect 2818 5296 3060 5324
rect 2818 5293 2830 5296
rect 2772 5287 2830 5293
rect 3048 5293 3060 5296
rect 3094 5293 3106 5327
rect 3048 5287 3106 5293
rect 4166 5319 4224 5325
rect 4166 5285 4178 5319
rect 4212 5316 4224 5319
rect 4252 5316 4280 5492
rect 4350 5387 4408 5393
rect 4350 5353 4362 5387
rect 4396 5384 4408 5387
rect 5090 5387 5148 5393
rect 5090 5384 5102 5387
rect 4396 5356 5102 5384
rect 4396 5353 4408 5356
rect 4350 5347 4408 5353
rect 5090 5353 5102 5356
rect 5136 5353 5148 5387
rect 5090 5347 5148 5353
rect 4534 5319 4592 5325
rect 4534 5316 4546 5319
rect 4212 5288 4546 5316
rect 4212 5285 4224 5288
rect 4166 5279 4224 5285
rect 4534 5285 4546 5288
rect 4580 5316 4592 5319
rect 4906 5319 4964 5325
rect 4906 5316 4918 5319
rect 4580 5288 4918 5316
rect 4580 5285 4592 5288
rect 4534 5279 4592 5285
rect 4906 5285 4918 5288
rect 4952 5316 4964 5319
rect 5182 5319 5240 5325
rect 5182 5316 5194 5319
rect 4952 5288 5194 5316
rect 4952 5285 4964 5288
rect 4906 5279 4964 5285
rect 5182 5285 5194 5288
rect 5228 5285 5240 5319
rect 5182 5279 5240 5285
rect 6118 5319 6176 5325
rect 6118 5285 6130 5319
rect 6164 5316 6176 5319
rect 6204 5316 6232 5492
rect 6302 5387 6360 5393
rect 6302 5353 6314 5387
rect 6348 5384 6360 5387
rect 7042 5387 7100 5393
rect 7042 5384 7054 5387
rect 6348 5356 7054 5384
rect 6348 5353 6360 5356
rect 6302 5347 6360 5353
rect 7042 5353 7054 5356
rect 7088 5353 7100 5387
rect 7042 5347 7100 5353
rect 8120 5325 8178 5331
rect 6486 5319 6544 5325
rect 6486 5316 6498 5319
rect 6164 5288 6498 5316
rect 6164 5285 6176 5288
rect 6118 5279 6176 5285
rect 6486 5285 6498 5288
rect 6532 5316 6544 5319
rect 6858 5319 6916 5325
rect 6858 5316 6870 5319
rect 6532 5288 6870 5316
rect 6532 5285 6544 5288
rect 6486 5279 6544 5285
rect 6858 5285 6870 5288
rect 6904 5316 6916 5319
rect 7134 5319 7192 5325
rect 7134 5316 7146 5319
rect 6904 5288 7146 5316
rect 6904 5285 6916 5288
rect 6858 5279 6916 5285
rect 7134 5285 7146 5288
rect 7180 5285 7192 5319
rect 8120 5291 8132 5325
rect 8166 5322 8178 5325
rect 8206 5322 8234 5498
rect 10860 5472 10888 5648
rect 11138 5645 11150 5648
rect 11184 5645 11196 5679
rect 14326 5675 14384 5681
rect 11138 5639 11196 5645
rect 12368 5667 12426 5673
rect 12368 5633 12380 5667
rect 12414 5664 12426 5667
rect 12828 5667 12886 5673
rect 12828 5664 12840 5667
rect 12414 5636 12840 5664
rect 12414 5633 12426 5636
rect 11412 5606 11472 5630
rect 12368 5627 12426 5633
rect 12828 5633 12840 5636
rect 12874 5664 12886 5667
rect 13200 5667 13258 5673
rect 13200 5664 13212 5667
rect 12874 5636 13212 5664
rect 12874 5633 12886 5636
rect 12828 5627 12886 5633
rect 11412 5570 11426 5606
rect 11466 5604 11472 5606
rect 11466 5596 11818 5604
rect 12464 5600 12524 5606
rect 12464 5596 12478 5600
rect 11466 5570 12478 5596
rect 11412 5566 12478 5570
rect 12512 5566 12524 5600
rect 11412 5554 11472 5566
rect 11804 5562 12524 5566
rect 11896 5558 12524 5562
rect 12464 5544 12524 5558
rect 10018 5452 11490 5472
rect 12922 5460 12950 5636
rect 13200 5633 13212 5636
rect 13246 5633 13258 5667
rect 14326 5641 14338 5675
rect 14372 5672 14384 5675
rect 14786 5675 14844 5681
rect 14786 5672 14798 5675
rect 14372 5644 14798 5672
rect 14372 5641 14384 5644
rect 14326 5635 14384 5641
rect 14786 5641 14798 5644
rect 14832 5672 14844 5675
rect 15158 5675 15216 5681
rect 15158 5672 15170 5675
rect 14832 5644 15170 5672
rect 14832 5641 14844 5644
rect 14786 5635 14844 5641
rect 13200 5627 13258 5633
rect 13482 5594 13534 5612
rect 14422 5608 14482 5614
rect 14422 5604 14436 5608
rect 13480 5558 13494 5594
rect 13528 5558 13588 5594
rect 13854 5574 14436 5604
rect 14470 5574 14482 5608
rect 13854 5566 14482 5574
rect 13480 5556 13588 5558
rect 13482 5546 13534 5556
rect 14422 5552 14482 5566
rect 14880 5468 14908 5644
rect 15158 5641 15170 5644
rect 15204 5641 15216 5675
rect 16320 5647 16332 5681
rect 16366 5678 16378 5681
rect 16780 5681 16838 5687
rect 16780 5678 16792 5681
rect 16366 5650 16792 5678
rect 16366 5647 16378 5650
rect 16320 5641 16378 5647
rect 16780 5647 16792 5650
rect 16826 5678 16838 5681
rect 17152 5681 17210 5687
rect 17152 5678 17164 5681
rect 16826 5650 17164 5678
rect 16826 5647 16838 5650
rect 16780 5641 16838 5647
rect 15158 5635 15216 5641
rect 15440 5602 15492 5620
rect 16416 5614 16476 5620
rect 16416 5610 16430 5614
rect 15848 5606 16430 5610
rect 15524 5602 16430 5606
rect 15438 5566 15452 5602
rect 15486 5580 16430 5602
rect 16464 5580 16476 5614
rect 15486 5572 16476 5580
rect 15486 5566 15884 5572
rect 15438 5564 15884 5566
rect 15440 5554 15492 5564
rect 16416 5558 16476 5572
rect 16874 5474 16902 5650
rect 17152 5647 17164 5650
rect 17198 5647 17210 5681
rect 17152 5641 17210 5647
rect 17434 5608 17486 5626
rect 17432 5572 17446 5608
rect 17480 5596 17540 5608
rect 17480 5572 17822 5596
rect 17432 5570 17822 5572
rect 17434 5564 17822 5570
rect 17434 5560 17514 5564
rect 10018 5441 11214 5452
rect 11270 5441 11490 5452
rect 10018 5407 10047 5441
rect 10081 5407 10139 5441
rect 10173 5407 10231 5441
rect 10265 5407 10323 5441
rect 10357 5407 10415 5441
rect 10449 5407 10507 5441
rect 10541 5407 10599 5441
rect 10633 5407 10691 5441
rect 10725 5407 10783 5441
rect 10817 5407 10875 5441
rect 10909 5407 10967 5441
rect 11001 5407 11059 5441
rect 11093 5407 11151 5441
rect 11185 5407 11214 5441
rect 11277 5407 11335 5441
rect 11369 5407 11427 5441
rect 11461 5407 11490 5441
rect 8304 5393 8362 5399
rect 8304 5359 8316 5393
rect 8350 5390 8362 5393
rect 9044 5393 9102 5399
rect 9044 5390 9056 5393
rect 8350 5362 9056 5390
rect 8350 5359 8362 5362
rect 8304 5353 8362 5359
rect 9044 5359 9056 5362
rect 9090 5359 9102 5393
rect 10018 5394 11214 5407
rect 11270 5394 11490 5407
rect 10018 5376 11490 5394
rect 12080 5440 13552 5460
rect 12080 5429 12800 5440
rect 12856 5429 13552 5440
rect 12080 5395 12109 5429
rect 12143 5395 12201 5429
rect 12235 5395 12293 5429
rect 12327 5395 12385 5429
rect 12419 5395 12477 5429
rect 12511 5395 12569 5429
rect 12603 5395 12661 5429
rect 12695 5395 12753 5429
rect 12787 5395 12800 5429
rect 12879 5395 12937 5429
rect 12971 5395 13029 5429
rect 13063 5395 13121 5429
rect 13155 5395 13213 5429
rect 13247 5395 13305 5429
rect 13339 5395 13397 5429
rect 13431 5395 13489 5429
rect 13523 5395 13552 5429
rect 12080 5382 12800 5395
rect 12856 5382 13552 5395
rect 12080 5364 13552 5382
rect 14038 5448 15510 5468
rect 14038 5437 14758 5448
rect 14814 5437 15510 5448
rect 14038 5403 14067 5437
rect 14101 5403 14159 5437
rect 14193 5403 14251 5437
rect 14285 5403 14343 5437
rect 14377 5403 14435 5437
rect 14469 5403 14527 5437
rect 14561 5403 14619 5437
rect 14653 5403 14711 5437
rect 14745 5403 14758 5437
rect 14837 5403 14895 5437
rect 14929 5403 14987 5437
rect 15021 5403 15079 5437
rect 15113 5403 15171 5437
rect 15205 5403 15263 5437
rect 15297 5403 15355 5437
rect 15389 5403 15447 5437
rect 15481 5403 15510 5437
rect 14038 5390 14758 5403
rect 14814 5390 15510 5403
rect 14038 5372 15510 5390
rect 16032 5454 17504 5474
rect 16032 5443 16752 5454
rect 16808 5443 17504 5454
rect 16032 5409 16061 5443
rect 16095 5409 16153 5443
rect 16187 5409 16245 5443
rect 16279 5409 16337 5443
rect 16371 5409 16429 5443
rect 16463 5409 16521 5443
rect 16555 5409 16613 5443
rect 16647 5409 16705 5443
rect 16739 5409 16752 5443
rect 16831 5409 16889 5443
rect 16923 5409 16981 5443
rect 17015 5409 17073 5443
rect 17107 5409 17165 5443
rect 17199 5409 17257 5443
rect 17291 5409 17349 5443
rect 17383 5409 17441 5443
rect 17475 5409 17504 5443
rect 16032 5396 16752 5409
rect 16808 5396 17504 5409
rect 16032 5378 17504 5396
rect 9044 5353 9102 5359
rect 8488 5325 8546 5331
rect 8488 5322 8500 5325
rect 8166 5294 8500 5322
rect 8166 5291 8178 5294
rect 8120 5285 8178 5291
rect 8488 5291 8500 5294
rect 8534 5322 8546 5325
rect 8860 5325 8918 5331
rect 8860 5322 8872 5325
rect 8534 5294 8872 5322
rect 8534 5291 8546 5294
rect 8488 5285 8546 5291
rect 8860 5291 8872 5294
rect 8906 5322 8918 5325
rect 9136 5325 9194 5331
rect 9136 5322 9148 5325
rect 8906 5294 9148 5322
rect 8906 5291 8918 5294
rect 8860 5285 8918 5291
rect 9136 5291 9148 5294
rect 9182 5291 9194 5325
rect 9136 5285 9194 5291
rect 17790 5302 17822 5564
rect 7134 5279 7192 5285
rect 17790 5270 18732 5302
rect 2124 5259 2182 5265
rect 2124 5225 2136 5259
rect 2170 5256 2182 5259
rect 2584 5259 2642 5265
rect 2584 5256 2596 5259
rect 2170 5228 2596 5256
rect 2170 5225 2182 5228
rect 2124 5219 2182 5225
rect 2584 5225 2596 5228
rect 2630 5256 2642 5259
rect 2956 5259 3014 5265
rect 2956 5256 2968 5259
rect 2630 5228 2968 5256
rect 2630 5225 2642 5228
rect 2584 5219 2642 5225
rect 2222 5198 2288 5200
rect 2222 5146 2228 5198
rect 2280 5146 2288 5198
rect 2222 5142 2288 5146
rect 2678 5052 2706 5228
rect 2956 5225 2968 5228
rect 3002 5225 3014 5259
rect 8212 5257 8270 5263
rect 2956 5219 3014 5225
rect 4258 5251 4316 5257
rect 4258 5217 4270 5251
rect 4304 5248 4316 5251
rect 4718 5251 4776 5257
rect 4718 5248 4730 5251
rect 4304 5220 4730 5248
rect 4304 5217 4316 5220
rect 4258 5211 4316 5217
rect 4718 5217 4730 5220
rect 4764 5248 4776 5251
rect 5090 5251 5148 5257
rect 5090 5248 5102 5251
rect 4764 5220 5102 5248
rect 4764 5217 4776 5220
rect 4718 5211 4776 5217
rect 3230 5186 3290 5210
rect 3230 5150 3244 5186
rect 3284 5184 3290 5186
rect 4354 5184 4414 5190
rect 3284 5180 3837 5184
rect 4354 5180 4368 5184
rect 3284 5150 4368 5180
rect 4402 5150 4414 5184
rect 3230 5146 4414 5150
rect 3230 5134 3290 5146
rect 3636 5142 4414 5146
rect 4354 5128 4414 5142
rect 1836 5040 3308 5052
rect 4812 5044 4840 5220
rect 5090 5217 5102 5220
rect 5136 5217 5148 5251
rect 5090 5211 5148 5217
rect 6210 5251 6268 5257
rect 6210 5217 6222 5251
rect 6256 5248 6268 5251
rect 6670 5251 6728 5257
rect 6670 5248 6682 5251
rect 6256 5220 6682 5248
rect 6256 5217 6268 5220
rect 6210 5211 6268 5217
rect 6670 5217 6682 5220
rect 6716 5248 6728 5251
rect 7042 5251 7100 5257
rect 7042 5248 7054 5251
rect 6716 5220 7054 5248
rect 6716 5217 6728 5220
rect 6670 5211 6728 5217
rect 5372 5178 5424 5196
rect 6306 5184 6366 5190
rect 6306 5180 6320 5184
rect 5612 5178 6320 5180
rect 5370 5142 5384 5178
rect 5418 5150 6320 5178
rect 6354 5150 6366 5184
rect 5418 5142 6366 5150
rect 5370 5140 5659 5142
rect 5372 5130 5424 5140
rect 6306 5128 6366 5142
rect 6764 5044 6792 5220
rect 7042 5217 7054 5220
rect 7088 5217 7100 5251
rect 8212 5223 8224 5257
rect 8258 5254 8270 5257
rect 8672 5257 8730 5263
rect 8672 5254 8684 5257
rect 8258 5226 8684 5254
rect 8258 5223 8270 5226
rect 8212 5217 8270 5223
rect 8672 5223 8684 5226
rect 8718 5254 8730 5257
rect 9044 5257 9102 5263
rect 9044 5254 9056 5257
rect 8718 5226 9056 5254
rect 8718 5223 8730 5226
rect 8672 5217 8730 5223
rect 7042 5211 7100 5217
rect 7324 5178 7376 5196
rect 8308 5190 8368 5196
rect 8308 5186 8322 5190
rect 7550 5178 8322 5186
rect 7322 5142 7336 5178
rect 7370 5156 8322 5178
rect 8356 5156 8368 5190
rect 7370 5148 8368 5156
rect 7370 5142 7611 5148
rect 7322 5140 7611 5142
rect 7324 5130 7376 5140
rect 8308 5134 8368 5148
rect 8766 5050 8794 5226
rect 9044 5223 9056 5226
rect 9090 5223 9102 5257
rect 9044 5217 9102 5223
rect 9906 5210 17524 5242
rect 9326 5184 9378 5202
rect 9906 5184 9938 5210
rect 9324 5148 9338 5184
rect 9372 5148 9938 5184
rect 9324 5146 9938 5148
rect 9326 5136 9378 5146
rect 9762 5144 9938 5146
rect 17492 5146 17524 5210
rect 18598 5222 18648 5242
rect 18598 5188 18608 5222
rect 18642 5188 18648 5222
rect 10046 5120 11518 5142
rect 10046 5111 10188 5120
rect 10244 5111 11518 5120
rect 17492 5114 18178 5146
rect 18598 5134 18648 5188
rect 18678 5194 18732 5270
rect 18678 5160 18690 5194
rect 18724 5160 18732 5194
rect 10046 5077 10075 5111
rect 10109 5077 10167 5111
rect 10244 5077 10259 5111
rect 10293 5077 10351 5111
rect 10385 5077 10443 5111
rect 10477 5077 10535 5111
rect 10569 5077 10627 5111
rect 10661 5077 10719 5111
rect 10753 5077 10811 5111
rect 10845 5077 10903 5111
rect 10937 5077 10995 5111
rect 11029 5077 11087 5111
rect 11121 5077 11179 5111
rect 11213 5077 11271 5111
rect 11305 5077 11363 5111
rect 11397 5077 11455 5111
rect 11489 5077 11518 5111
rect 18146 5102 18178 5114
rect 18426 5108 18480 5120
rect 18250 5102 18432 5108
rect 10046 5062 10188 5077
rect 10244 5062 11518 5077
rect 1836 5021 2584 5040
rect 2640 5021 3308 5040
rect 1836 4987 1865 5021
rect 1899 4987 1957 5021
rect 1991 4987 2049 5021
rect 2083 4987 2141 5021
rect 2175 4987 2233 5021
rect 2267 4987 2325 5021
rect 2359 4987 2417 5021
rect 2451 4987 2509 5021
rect 2543 4987 2584 5021
rect 2640 4987 2693 5021
rect 2727 4987 2785 5021
rect 2819 4987 2877 5021
rect 2911 4987 2969 5021
rect 3003 4987 3061 5021
rect 3095 4987 3153 5021
rect 3187 4987 3245 5021
rect 3279 4987 3308 5021
rect 1836 4982 2584 4987
rect 2640 4982 3308 4987
rect 1836 4956 3308 4982
rect 3970 5024 5442 5044
rect 3970 5013 4690 5024
rect 4746 5013 5442 5024
rect 3970 4979 3999 5013
rect 4033 4979 4091 5013
rect 4125 4979 4183 5013
rect 4217 4979 4275 5013
rect 4309 4979 4367 5013
rect 4401 4979 4459 5013
rect 4493 4979 4551 5013
rect 4585 4979 4643 5013
rect 4677 4979 4690 5013
rect 4769 4979 4827 5013
rect 4861 4979 4919 5013
rect 4953 4979 5011 5013
rect 5045 4979 5103 5013
rect 5137 4979 5195 5013
rect 5229 4979 5287 5013
rect 5321 4979 5379 5013
rect 5413 4979 5442 5013
rect 3970 4966 4690 4979
rect 4746 4966 5442 4979
rect 3970 4948 5442 4966
rect 5922 5024 7394 5044
rect 5922 5013 6642 5024
rect 6698 5013 7394 5024
rect 5922 4979 5951 5013
rect 5985 4979 6043 5013
rect 6077 4979 6135 5013
rect 6169 4979 6227 5013
rect 6261 4979 6319 5013
rect 6353 4979 6411 5013
rect 6445 4979 6503 5013
rect 6537 4979 6595 5013
rect 6629 4979 6642 5013
rect 6721 4979 6779 5013
rect 6813 4979 6871 5013
rect 6905 4979 6963 5013
rect 6997 4979 7055 5013
rect 7089 4979 7147 5013
rect 7181 4979 7239 5013
rect 7273 4979 7331 5013
rect 7365 4979 7394 5013
rect 5922 4966 6642 4979
rect 6698 4966 7394 4979
rect 5922 4948 7394 4966
rect 7924 5030 9396 5050
rect 10046 5046 11518 5062
rect 12316 5080 13788 5098
rect 12316 5067 13032 5080
rect 13088 5067 13788 5080
rect 7924 5019 8644 5030
rect 8700 5019 9396 5030
rect 7924 4985 7953 5019
rect 7987 4985 8045 5019
rect 8079 4985 8137 5019
rect 8171 4985 8229 5019
rect 8263 4985 8321 5019
rect 8355 4985 8413 5019
rect 8447 4985 8505 5019
rect 8539 4985 8597 5019
rect 8631 4985 8644 5019
rect 8723 4985 8781 5019
rect 8815 4985 8873 5019
rect 8907 4985 8965 5019
rect 8999 4985 9057 5019
rect 9091 4985 9149 5019
rect 9183 4985 9241 5019
rect 9275 4985 9333 5019
rect 9367 4985 9396 5019
rect 7924 4972 8644 4985
rect 8700 4972 9396 4985
rect 7924 4954 9396 4972
rect 10242 4873 10300 4879
rect 10242 4839 10254 4873
rect 10288 4870 10300 4873
rect 10328 4870 10356 5046
rect 12316 5033 12345 5067
rect 12379 5033 12437 5067
rect 12471 5033 12529 5067
rect 12563 5033 12621 5067
rect 12655 5033 12713 5067
rect 12747 5033 12805 5067
rect 12839 5033 12897 5067
rect 12931 5033 12989 5067
rect 13023 5033 13032 5067
rect 13115 5033 13173 5067
rect 13207 5033 13265 5067
rect 13299 5033 13357 5067
rect 13391 5033 13449 5067
rect 13483 5033 13541 5067
rect 13575 5033 13633 5067
rect 13667 5033 13725 5067
rect 13759 5033 13788 5067
rect 12316 5022 13032 5033
rect 13088 5022 13788 5033
rect 12316 5002 13788 5022
rect 14318 5074 15790 5092
rect 14318 5061 15034 5074
rect 15090 5061 15790 5074
rect 14318 5027 14347 5061
rect 14381 5027 14439 5061
rect 14473 5027 14531 5061
rect 14565 5027 14623 5061
rect 14657 5027 14715 5061
rect 14749 5027 14807 5061
rect 14841 5027 14899 5061
rect 14933 5027 14991 5061
rect 15025 5027 15034 5061
rect 15117 5027 15175 5061
rect 15209 5027 15267 5061
rect 15301 5027 15359 5061
rect 15393 5027 15451 5061
rect 15485 5027 15543 5061
rect 15577 5027 15635 5061
rect 15669 5027 15727 5061
rect 15761 5027 15790 5061
rect 14318 5016 15034 5027
rect 15090 5016 15790 5027
rect 10426 4941 10484 4947
rect 10426 4907 10438 4941
rect 10472 4938 10484 4941
rect 11166 4941 11224 4947
rect 11166 4938 11178 4941
rect 10472 4910 11178 4938
rect 10472 4907 10484 4910
rect 10426 4901 10484 4907
rect 11166 4907 11178 4910
rect 11212 4907 11224 4941
rect 11166 4901 11224 4907
rect 10610 4873 10668 4879
rect 10610 4870 10622 4873
rect 10288 4842 10622 4870
rect 10288 4839 10300 4842
rect 10242 4833 10300 4839
rect 10610 4839 10622 4842
rect 10656 4870 10668 4873
rect 10982 4873 11040 4879
rect 10982 4870 10994 4873
rect 10656 4842 10994 4870
rect 10656 4839 10668 4842
rect 10610 4833 10668 4839
rect 10982 4839 10994 4842
rect 11028 4870 11040 4873
rect 11258 4873 11316 4879
rect 11258 4870 11270 4873
rect 11028 4842 11270 4870
rect 11028 4839 11040 4842
rect 10982 4833 11040 4839
rect 11258 4839 11270 4842
rect 11304 4839 11316 4873
rect 11258 4833 11316 4839
rect 12512 4829 12570 4835
rect 10334 4805 10392 4811
rect 10334 4771 10346 4805
rect 10380 4802 10392 4805
rect 10794 4805 10852 4811
rect 10794 4802 10806 4805
rect 10380 4774 10806 4802
rect 10380 4771 10392 4774
rect 10334 4765 10392 4771
rect 10794 4771 10806 4774
rect 10840 4802 10852 4805
rect 11166 4805 11224 4811
rect 11166 4802 11178 4805
rect 10840 4774 11178 4802
rect 10840 4771 10852 4774
rect 10794 4765 10852 4771
rect 10432 4744 10498 4746
rect 10432 4692 10438 4744
rect 10490 4692 10498 4744
rect 10432 4688 10498 4692
rect 10888 4598 10916 4774
rect 11166 4771 11178 4774
rect 11212 4771 11224 4805
rect 12512 4795 12524 4829
rect 12558 4826 12570 4829
rect 12598 4826 12626 5002
rect 14318 4996 15790 5016
rect 16340 5056 17812 5074
rect 18146 5070 18432 5102
rect 18470 5070 18572 5108
rect 16340 5043 17056 5056
rect 17112 5043 17812 5056
rect 18426 5054 18480 5070
rect 16340 5009 16369 5043
rect 16403 5009 16461 5043
rect 16495 5009 16553 5043
rect 16587 5009 16645 5043
rect 16679 5009 16737 5043
rect 16771 5009 16829 5043
rect 16863 5009 16921 5043
rect 16955 5009 17013 5043
rect 17047 5009 17056 5043
rect 17139 5009 17197 5043
rect 17231 5009 17289 5043
rect 17323 5009 17381 5043
rect 17415 5009 17473 5043
rect 17507 5009 17565 5043
rect 17599 5009 17657 5043
rect 17691 5009 17749 5043
rect 17783 5009 17812 5043
rect 18608 5024 18640 5134
rect 18678 5114 18732 5160
rect 18678 5110 18716 5114
rect 18250 5023 18640 5024
rect 16340 4998 17056 5009
rect 17112 4998 17812 5009
rect 12696 4897 12754 4903
rect 12696 4863 12708 4897
rect 12742 4894 12754 4897
rect 13436 4897 13494 4903
rect 13436 4894 13448 4897
rect 12742 4866 13448 4894
rect 12742 4863 12754 4866
rect 12696 4857 12754 4863
rect 13436 4863 13448 4866
rect 13482 4863 13494 4897
rect 13436 4857 13494 4863
rect 12880 4829 12938 4835
rect 12880 4826 12892 4829
rect 12558 4798 12892 4826
rect 12558 4795 12570 4798
rect 12512 4789 12570 4795
rect 12880 4795 12892 4798
rect 12926 4826 12938 4829
rect 13252 4829 13310 4835
rect 13252 4826 13264 4829
rect 12926 4798 13264 4826
rect 12926 4795 12938 4798
rect 12880 4789 12938 4795
rect 13252 4795 13264 4798
rect 13298 4826 13310 4829
rect 13528 4829 13586 4835
rect 13528 4826 13540 4829
rect 13298 4798 13540 4826
rect 13298 4795 13310 4798
rect 13252 4789 13310 4795
rect 13528 4795 13540 4798
rect 13574 4795 13586 4829
rect 13528 4789 13586 4795
rect 14514 4823 14572 4829
rect 14514 4789 14526 4823
rect 14560 4820 14572 4823
rect 14600 4820 14628 4996
rect 16340 4978 17812 4998
rect 18169 4992 18640 5023
rect 19046 5050 19112 5098
rect 19046 4998 19056 5050
rect 19108 4998 19112 5050
rect 18169 4985 18277 4992
rect 14698 4891 14756 4897
rect 14698 4857 14710 4891
rect 14744 4888 14756 4891
rect 15438 4891 15496 4897
rect 15438 4888 15450 4891
rect 14744 4860 15450 4888
rect 14744 4857 14756 4860
rect 14698 4851 14756 4857
rect 15438 4857 15450 4860
rect 15484 4857 15496 4891
rect 15438 4851 15496 4857
rect 14882 4823 14940 4829
rect 14882 4820 14894 4823
rect 14560 4792 14894 4820
rect 14560 4789 14572 4792
rect 14514 4783 14572 4789
rect 14882 4789 14894 4792
rect 14928 4820 14940 4823
rect 15254 4823 15312 4829
rect 15254 4820 15266 4823
rect 14928 4792 15266 4820
rect 14928 4789 14940 4792
rect 14882 4783 14940 4789
rect 15254 4789 15266 4792
rect 15300 4820 15312 4823
rect 15530 4823 15588 4829
rect 15530 4820 15542 4823
rect 15300 4792 15542 4820
rect 15300 4789 15312 4792
rect 15254 4783 15312 4789
rect 15530 4789 15542 4792
rect 15576 4789 15588 4823
rect 15530 4783 15588 4789
rect 16536 4805 16594 4811
rect 11166 4765 11224 4771
rect 16536 4771 16548 4805
rect 16582 4802 16594 4805
rect 16622 4802 16650 4978
rect 16720 4873 16778 4879
rect 16720 4839 16732 4873
rect 16766 4870 16778 4873
rect 17460 4873 17518 4879
rect 17460 4870 17472 4873
rect 16766 4842 17472 4870
rect 16766 4839 16778 4842
rect 16720 4833 16778 4839
rect 17460 4839 17472 4842
rect 17506 4839 17518 4873
rect 17460 4833 17518 4839
rect 16904 4805 16962 4811
rect 16904 4802 16916 4805
rect 16582 4774 16916 4802
rect 16582 4771 16594 4774
rect 12604 4761 12662 4767
rect 11440 4732 11500 4756
rect 11440 4696 11454 4732
rect 11494 4730 11500 4732
rect 11494 4712 11818 4730
rect 12604 4727 12616 4761
rect 12650 4758 12662 4761
rect 13064 4761 13122 4767
rect 13064 4758 13076 4761
rect 12650 4730 13076 4758
rect 12650 4727 12662 4730
rect 12604 4721 12662 4727
rect 13064 4727 13076 4730
rect 13110 4758 13122 4761
rect 13436 4761 13494 4767
rect 16536 4765 16594 4771
rect 16904 4771 16916 4774
rect 16950 4802 16962 4805
rect 17276 4805 17334 4811
rect 17276 4802 17288 4805
rect 16950 4774 17288 4802
rect 16950 4771 16962 4774
rect 16904 4765 16962 4771
rect 17276 4771 17288 4774
rect 17322 4802 17334 4805
rect 17552 4805 17610 4811
rect 17552 4802 17564 4805
rect 17322 4774 17564 4802
rect 17322 4771 17334 4774
rect 17276 4765 17334 4771
rect 17552 4771 17564 4774
rect 17598 4771 17610 4805
rect 17552 4765 17610 4771
rect 13436 4758 13448 4761
rect 13110 4730 13448 4758
rect 13110 4727 13122 4730
rect 13064 4721 13122 4727
rect 11494 4696 12102 4712
rect 11440 4692 12102 4696
rect 11440 4680 11500 4692
rect 11774 4690 12102 4692
rect 12700 4694 12760 4700
rect 12700 4690 12714 4694
rect 11774 4660 12714 4690
rect 12748 4660 12760 4694
rect 11774 4652 12760 4660
rect 12700 4638 12760 4652
rect 10046 4580 11518 4598
rect 10046 4567 10788 4580
rect 10844 4567 11518 4580
rect 10046 4533 10075 4567
rect 10109 4533 10167 4567
rect 10201 4533 10259 4567
rect 10293 4533 10351 4567
rect 10385 4566 10443 4567
rect 10477 4566 10535 4567
rect 10385 4533 10440 4566
rect 10492 4533 10535 4566
rect 10569 4533 10627 4567
rect 10661 4533 10719 4567
rect 10753 4533 10788 4567
rect 10845 4533 10903 4567
rect 10937 4533 10995 4567
rect 11029 4533 11087 4567
rect 11121 4533 11179 4567
rect 11213 4533 11271 4567
rect 11305 4533 11363 4567
rect 11397 4533 11455 4567
rect 11489 4533 11518 4567
rect 13158 4554 13186 4730
rect 13436 4727 13448 4730
rect 13482 4727 13494 4761
rect 13436 4721 13494 4727
rect 14606 4755 14664 4761
rect 14606 4721 14618 4755
rect 14652 4752 14664 4755
rect 15066 4755 15124 4761
rect 15066 4752 15078 4755
rect 14652 4724 15078 4752
rect 14652 4721 14664 4724
rect 14606 4715 14664 4721
rect 15066 4721 15078 4724
rect 15112 4752 15124 4755
rect 15438 4755 15496 4761
rect 15438 4752 15450 4755
rect 15112 4724 15450 4752
rect 15112 4721 15124 4724
rect 15066 4715 15124 4721
rect 13718 4688 13770 4706
rect 14702 4688 14762 4694
rect 13716 4652 13730 4688
rect 13764 4684 14105 4688
rect 14702 4684 14716 4688
rect 13764 4654 14716 4684
rect 14750 4654 14762 4688
rect 13764 4652 14762 4654
rect 13716 4650 14762 4652
rect 13718 4640 13770 4650
rect 14082 4646 14762 4650
rect 14702 4632 14762 4646
rect 10046 4512 10440 4533
rect 10492 4522 10788 4533
rect 10844 4522 11518 4533
rect 10492 4512 11518 4522
rect 10046 4502 11518 4512
rect 12316 4534 13788 4554
rect 15160 4548 15188 4724
rect 15438 4721 15450 4724
rect 15484 4721 15496 4755
rect 15438 4715 15496 4721
rect 16628 4737 16686 4743
rect 16628 4703 16640 4737
rect 16674 4734 16686 4737
rect 17088 4737 17146 4743
rect 17088 4734 17100 4737
rect 16674 4706 17100 4734
rect 16674 4703 16686 4706
rect 15720 4682 15772 4700
rect 16628 4697 16686 4703
rect 17088 4703 17100 4706
rect 17134 4734 17146 4737
rect 17460 4737 17518 4743
rect 17460 4734 17472 4737
rect 17134 4706 17472 4734
rect 17134 4703 17146 4706
rect 17088 4697 17146 4703
rect 15718 4646 15732 4682
rect 15766 4666 15870 4682
rect 16724 4670 16784 4676
rect 16724 4666 16738 4670
rect 15766 4646 16738 4666
rect 15718 4644 16738 4646
rect 15720 4634 15772 4644
rect 15845 4636 16738 4644
rect 16772 4636 16784 4670
rect 15845 4628 16784 4636
rect 16724 4614 16784 4628
rect 12316 4523 13036 4534
rect 13092 4523 13788 4534
rect 12316 4489 12345 4523
rect 12379 4489 12437 4523
rect 12471 4489 12529 4523
rect 12563 4489 12621 4523
rect 12655 4489 12713 4523
rect 12747 4489 12805 4523
rect 12839 4489 12897 4523
rect 12931 4489 12989 4523
rect 13023 4489 13036 4523
rect 13115 4489 13173 4523
rect 13207 4489 13265 4523
rect 13299 4489 13357 4523
rect 13391 4489 13449 4523
rect 13483 4489 13541 4523
rect 13575 4489 13633 4523
rect 13667 4489 13725 4523
rect 13759 4489 13788 4523
rect 12316 4476 13036 4489
rect 13092 4476 13788 4489
rect 12316 4458 13788 4476
rect 14318 4528 15790 4548
rect 17182 4530 17210 4706
rect 17460 4703 17472 4706
rect 17506 4703 17518 4737
rect 17460 4697 17518 4703
rect 17742 4664 17794 4682
rect 18169 4664 18207 4985
rect 19046 4944 19112 4998
rect 17740 4628 17754 4664
rect 17788 4628 18207 4664
rect 17740 4626 18207 4628
rect 17742 4616 17794 4626
rect 14318 4517 15038 4528
rect 15094 4517 15790 4528
rect 14318 4483 14347 4517
rect 14381 4483 14439 4517
rect 14473 4483 14531 4517
rect 14565 4483 14623 4517
rect 14657 4483 14715 4517
rect 14749 4483 14807 4517
rect 14841 4483 14899 4517
rect 14933 4483 14991 4517
rect 15025 4483 15038 4517
rect 15117 4483 15175 4517
rect 15209 4483 15267 4517
rect 15301 4483 15359 4517
rect 15393 4483 15451 4517
rect 15485 4483 15543 4517
rect 15577 4483 15635 4517
rect 15669 4483 15727 4517
rect 15761 4483 15790 4517
rect 14318 4470 15038 4483
rect 15094 4470 15790 4483
rect 14318 4452 15790 4470
rect 16340 4510 17812 4530
rect 16340 4499 17060 4510
rect 17116 4499 17812 4510
rect 16340 4465 16369 4499
rect 16403 4465 16461 4499
rect 16495 4465 16553 4499
rect 16587 4465 16645 4499
rect 16679 4465 16737 4499
rect 16771 4465 16829 4499
rect 16863 4465 16921 4499
rect 16955 4465 17013 4499
rect 17047 4465 17060 4499
rect 17139 4465 17197 4499
rect 17231 4465 17289 4499
rect 17323 4465 17381 4499
rect 17415 4465 17473 4499
rect 17507 4465 17565 4499
rect 17599 4465 17657 4499
rect 17691 4465 17749 4499
rect 17783 4465 17812 4499
rect 16340 4452 17060 4465
rect 17116 4452 17812 4465
rect 16340 4434 17812 4452
rect 6104 3130 6198 3138
rect 6104 3078 6138 3130
rect 6190 3078 6198 3130
rect 6232 3136 6298 3138
rect 6232 3084 6238 3136
rect 6290 3084 6298 3136
rect 6232 3078 6298 3084
rect 6104 3072 6198 3078
rect 1806 2318 3278 2336
rect 1806 2305 2604 2318
rect 2660 2305 3278 2318
rect 1806 2271 1835 2305
rect 1869 2271 1927 2305
rect 1961 2271 2019 2305
rect 2053 2271 2111 2305
rect 2145 2271 2203 2305
rect 2237 2271 2295 2305
rect 2329 2271 2387 2305
rect 2421 2271 2479 2305
rect 2513 2271 2571 2305
rect 2660 2271 2663 2305
rect 2697 2271 2755 2305
rect 2789 2271 2847 2305
rect 2881 2271 2939 2305
rect 2973 2271 3031 2305
rect 3065 2271 3123 2305
rect 3157 2271 3215 2305
rect 3249 2271 3278 2305
rect 1806 2260 2604 2271
rect 2660 2260 3278 2271
rect 1806 2240 3278 2260
rect 3876 2314 5348 2332
rect 3876 2301 4592 2314
rect 4648 2301 5348 2314
rect 3876 2267 3905 2301
rect 3939 2267 3997 2301
rect 4031 2267 4089 2301
rect 4123 2267 4181 2301
rect 4215 2267 4273 2301
rect 4307 2267 4365 2301
rect 4399 2267 4457 2301
rect 4491 2267 4549 2301
rect 4583 2267 4592 2301
rect 4675 2267 4733 2301
rect 4767 2267 4825 2301
rect 4859 2267 4917 2301
rect 4951 2267 5009 2301
rect 5043 2267 5101 2301
rect 5135 2267 5193 2301
rect 5227 2267 5285 2301
rect 5319 2267 5348 2301
rect 3876 2256 4592 2267
rect 4648 2256 5348 2267
rect 2002 2067 2060 2073
rect 2002 2033 2014 2067
rect 2048 2064 2060 2067
rect 2088 2064 2116 2240
rect 3876 2236 5348 2256
rect 5828 2314 7300 2332
rect 5828 2301 6544 2314
rect 6600 2301 7300 2314
rect 5828 2267 5857 2301
rect 5891 2267 5949 2301
rect 5983 2267 6041 2301
rect 6075 2267 6133 2301
rect 6167 2267 6225 2301
rect 6259 2267 6317 2301
rect 6351 2267 6409 2301
rect 6443 2267 6501 2301
rect 6535 2267 6544 2301
rect 6627 2267 6685 2301
rect 6719 2267 6777 2301
rect 6811 2267 6869 2301
rect 6903 2267 6961 2301
rect 6995 2267 7053 2301
rect 7087 2267 7145 2301
rect 7179 2267 7237 2301
rect 7271 2267 7300 2301
rect 5828 2256 6544 2267
rect 6600 2256 7300 2267
rect 5828 2236 7300 2256
rect 7830 2320 9302 2338
rect 7830 2307 8546 2320
rect 8602 2307 9302 2320
rect 7830 2273 7859 2307
rect 7893 2273 7951 2307
rect 7985 2273 8043 2307
rect 8077 2273 8135 2307
rect 8169 2273 8227 2307
rect 8261 2273 8319 2307
rect 8353 2273 8411 2307
rect 8445 2273 8503 2307
rect 8537 2273 8546 2307
rect 8629 2273 8687 2307
rect 8721 2273 8779 2307
rect 8813 2273 8871 2307
rect 8905 2273 8963 2307
rect 8997 2273 9055 2307
rect 9089 2273 9147 2307
rect 9181 2273 9239 2307
rect 9273 2273 9302 2307
rect 7830 2262 8546 2273
rect 8602 2262 9302 2273
rect 7830 2242 9302 2262
rect 9782 2320 11254 2338
rect 9782 2307 10498 2320
rect 10554 2307 11254 2320
rect 9782 2273 9811 2307
rect 9845 2273 9903 2307
rect 9937 2273 9995 2307
rect 10029 2273 10087 2307
rect 10121 2273 10179 2307
rect 10213 2273 10271 2307
rect 10305 2273 10363 2307
rect 10397 2273 10455 2307
rect 10489 2273 10498 2307
rect 10581 2273 10639 2307
rect 10673 2273 10731 2307
rect 10765 2273 10823 2307
rect 10857 2273 10915 2307
rect 10949 2273 11007 2307
rect 11041 2273 11099 2307
rect 11133 2273 11191 2307
rect 11225 2273 11254 2307
rect 9782 2262 10498 2273
rect 10554 2262 11254 2273
rect 9782 2242 11254 2262
rect 11774 2320 13246 2338
rect 11774 2307 12490 2320
rect 12546 2307 13246 2320
rect 11774 2273 11803 2307
rect 11837 2273 11895 2307
rect 11929 2273 11987 2307
rect 12021 2273 12079 2307
rect 12113 2273 12171 2307
rect 12205 2273 12263 2307
rect 12297 2273 12355 2307
rect 12389 2273 12447 2307
rect 12481 2273 12490 2307
rect 12573 2273 12631 2307
rect 12665 2273 12723 2307
rect 12757 2273 12815 2307
rect 12849 2273 12907 2307
rect 12941 2273 12999 2307
rect 13033 2273 13091 2307
rect 13125 2273 13183 2307
rect 13217 2273 13246 2307
rect 11774 2262 12490 2273
rect 12546 2262 13246 2273
rect 11774 2242 13246 2262
rect 13726 2320 15198 2338
rect 13726 2307 14442 2320
rect 14498 2307 15198 2320
rect 13726 2273 13755 2307
rect 13789 2273 13847 2307
rect 13881 2273 13939 2307
rect 13973 2273 14031 2307
rect 14065 2273 14123 2307
rect 14157 2273 14215 2307
rect 14249 2273 14307 2307
rect 14341 2273 14399 2307
rect 14433 2273 14442 2307
rect 14525 2273 14583 2307
rect 14617 2273 14675 2307
rect 14709 2273 14767 2307
rect 14801 2273 14859 2307
rect 14893 2273 14951 2307
rect 14985 2273 15043 2307
rect 15077 2273 15135 2307
rect 15169 2273 15198 2307
rect 13726 2262 14442 2273
rect 14498 2262 15198 2273
rect 13726 2242 15198 2262
rect 15790 2320 17262 2338
rect 15790 2307 16506 2320
rect 16562 2307 17262 2320
rect 15790 2273 15819 2307
rect 15853 2273 15911 2307
rect 15945 2273 16003 2307
rect 16037 2273 16095 2307
rect 16129 2273 16187 2307
rect 16221 2273 16279 2307
rect 16313 2273 16371 2307
rect 16405 2273 16463 2307
rect 16497 2273 16506 2307
rect 16589 2273 16647 2307
rect 16681 2273 16739 2307
rect 16773 2273 16831 2307
rect 16865 2273 16923 2307
rect 16957 2273 17015 2307
rect 17049 2273 17107 2307
rect 17141 2273 17199 2307
rect 17233 2273 17262 2307
rect 15790 2262 16506 2273
rect 16562 2262 17262 2273
rect 15790 2242 17262 2262
rect 2186 2135 2244 2141
rect 2186 2101 2198 2135
rect 2232 2132 2244 2135
rect 2926 2135 2984 2141
rect 2926 2132 2938 2135
rect 2232 2104 2938 2132
rect 2232 2101 2244 2104
rect 2186 2095 2244 2101
rect 2926 2101 2938 2104
rect 2972 2101 2984 2135
rect 2926 2095 2984 2101
rect 2370 2067 2428 2073
rect 2370 2064 2382 2067
rect 2048 2036 2382 2064
rect 2048 2033 2060 2036
rect 2002 2027 2060 2033
rect 2370 2033 2382 2036
rect 2416 2064 2428 2067
rect 2742 2067 2800 2073
rect 2742 2064 2754 2067
rect 2416 2036 2754 2064
rect 2416 2033 2428 2036
rect 2370 2027 2428 2033
rect 2742 2033 2754 2036
rect 2788 2064 2800 2067
rect 3018 2067 3076 2073
rect 3018 2064 3030 2067
rect 2788 2036 3030 2064
rect 2788 2033 2800 2036
rect 2742 2027 2800 2033
rect 3018 2033 3030 2036
rect 3064 2033 3076 2067
rect 3018 2027 3076 2033
rect 4072 2063 4130 2069
rect 4072 2029 4084 2063
rect 4118 2060 4130 2063
rect 4158 2060 4186 2236
rect 4256 2131 4314 2137
rect 4256 2097 4268 2131
rect 4302 2128 4314 2131
rect 4996 2131 5054 2137
rect 4996 2128 5008 2131
rect 4302 2100 5008 2128
rect 4302 2097 4314 2100
rect 4256 2091 4314 2097
rect 4996 2097 5008 2100
rect 5042 2097 5054 2131
rect 4996 2091 5054 2097
rect 4440 2063 4498 2069
rect 4440 2060 4452 2063
rect 4118 2032 4452 2060
rect 4118 2029 4130 2032
rect 4072 2023 4130 2029
rect 4440 2029 4452 2032
rect 4486 2060 4498 2063
rect 4812 2063 4870 2069
rect 4812 2060 4824 2063
rect 4486 2032 4824 2060
rect 4486 2029 4498 2032
rect 4440 2023 4498 2029
rect 4812 2029 4824 2032
rect 4858 2060 4870 2063
rect 5088 2063 5146 2069
rect 5088 2060 5100 2063
rect 4858 2032 5100 2060
rect 4858 2029 4870 2032
rect 4812 2023 4870 2029
rect 5088 2029 5100 2032
rect 5134 2029 5146 2063
rect 5088 2023 5146 2029
rect 6024 2063 6082 2069
rect 6024 2029 6036 2063
rect 6070 2060 6082 2063
rect 6110 2060 6138 2236
rect 6208 2131 6266 2137
rect 6208 2097 6220 2131
rect 6254 2128 6266 2131
rect 6948 2131 7006 2137
rect 6948 2128 6960 2131
rect 6254 2100 6960 2128
rect 6254 2097 6266 2100
rect 6208 2091 6266 2097
rect 6948 2097 6960 2100
rect 6994 2097 7006 2131
rect 6948 2091 7006 2097
rect 8026 2069 8084 2075
rect 6392 2063 6450 2069
rect 6392 2060 6404 2063
rect 6070 2032 6404 2060
rect 6070 2029 6082 2032
rect 6024 2023 6082 2029
rect 6392 2029 6404 2032
rect 6438 2060 6450 2063
rect 6764 2063 6822 2069
rect 6764 2060 6776 2063
rect 6438 2032 6776 2060
rect 6438 2029 6450 2032
rect 6392 2023 6450 2029
rect 6764 2029 6776 2032
rect 6810 2060 6822 2063
rect 7040 2063 7098 2069
rect 7040 2060 7052 2063
rect 6810 2032 7052 2060
rect 6810 2029 6822 2032
rect 6764 2023 6822 2029
rect 7040 2029 7052 2032
rect 7086 2029 7098 2063
rect 8026 2035 8038 2069
rect 8072 2066 8084 2069
rect 8112 2066 8140 2242
rect 8210 2137 8268 2143
rect 8210 2103 8222 2137
rect 8256 2134 8268 2137
rect 8950 2137 9008 2143
rect 8950 2134 8962 2137
rect 8256 2106 8962 2134
rect 8256 2103 8268 2106
rect 8210 2097 8268 2103
rect 8950 2103 8962 2106
rect 8996 2103 9008 2137
rect 8950 2097 9008 2103
rect 8394 2069 8452 2075
rect 8394 2066 8406 2069
rect 8072 2038 8406 2066
rect 8072 2035 8084 2038
rect 8026 2029 8084 2035
rect 8394 2035 8406 2038
rect 8440 2066 8452 2069
rect 8766 2069 8824 2075
rect 8766 2066 8778 2069
rect 8440 2038 8778 2066
rect 8440 2035 8452 2038
rect 8394 2029 8452 2035
rect 8766 2035 8778 2038
rect 8812 2066 8824 2069
rect 9042 2069 9100 2075
rect 9042 2066 9054 2069
rect 8812 2038 9054 2066
rect 8812 2035 8824 2038
rect 8766 2029 8824 2035
rect 9042 2035 9054 2038
rect 9088 2035 9100 2069
rect 9042 2029 9100 2035
rect 9978 2069 10036 2075
rect 9978 2035 9990 2069
rect 10024 2066 10036 2069
rect 10064 2066 10092 2242
rect 10162 2137 10220 2143
rect 10162 2103 10174 2137
rect 10208 2134 10220 2137
rect 10902 2137 10960 2143
rect 10902 2134 10914 2137
rect 10208 2106 10914 2134
rect 10208 2103 10220 2106
rect 10162 2097 10220 2103
rect 10902 2103 10914 2106
rect 10948 2103 10960 2137
rect 10902 2097 10960 2103
rect 10346 2069 10404 2075
rect 10346 2066 10358 2069
rect 10024 2038 10358 2066
rect 10024 2035 10036 2038
rect 9978 2029 10036 2035
rect 10346 2035 10358 2038
rect 10392 2066 10404 2069
rect 10718 2069 10776 2075
rect 10718 2066 10730 2069
rect 10392 2038 10730 2066
rect 10392 2035 10404 2038
rect 10346 2029 10404 2035
rect 10718 2035 10730 2038
rect 10764 2066 10776 2069
rect 10994 2069 11052 2075
rect 10994 2066 11006 2069
rect 10764 2038 11006 2066
rect 10764 2035 10776 2038
rect 10718 2029 10776 2035
rect 10994 2035 11006 2038
rect 11040 2035 11052 2069
rect 10994 2029 11052 2035
rect 11970 2069 12028 2075
rect 11970 2035 11982 2069
rect 12016 2066 12028 2069
rect 12056 2066 12084 2242
rect 12154 2137 12212 2143
rect 12154 2103 12166 2137
rect 12200 2134 12212 2137
rect 12894 2137 12952 2143
rect 12894 2134 12906 2137
rect 12200 2106 12906 2134
rect 12200 2103 12212 2106
rect 12154 2097 12212 2103
rect 12894 2103 12906 2106
rect 12940 2103 12952 2137
rect 12894 2097 12952 2103
rect 12338 2069 12396 2075
rect 12338 2066 12350 2069
rect 12016 2038 12350 2066
rect 12016 2035 12028 2038
rect 11970 2029 12028 2035
rect 12338 2035 12350 2038
rect 12384 2066 12396 2069
rect 12710 2069 12768 2075
rect 12710 2066 12722 2069
rect 12384 2038 12722 2066
rect 12384 2035 12396 2038
rect 12338 2029 12396 2035
rect 12710 2035 12722 2038
rect 12756 2066 12768 2069
rect 12986 2069 13044 2075
rect 12986 2066 12998 2069
rect 12756 2038 12998 2066
rect 12756 2035 12768 2038
rect 12710 2029 12768 2035
rect 12986 2035 12998 2038
rect 13032 2035 13044 2069
rect 12986 2029 13044 2035
rect 13922 2069 13980 2075
rect 13922 2035 13934 2069
rect 13968 2066 13980 2069
rect 14008 2066 14036 2242
rect 14106 2137 14164 2143
rect 14106 2103 14118 2137
rect 14152 2134 14164 2137
rect 14846 2137 14904 2143
rect 14846 2134 14858 2137
rect 14152 2106 14858 2134
rect 14152 2103 14164 2106
rect 14106 2097 14164 2103
rect 14846 2103 14858 2106
rect 14892 2103 14904 2137
rect 14846 2097 14904 2103
rect 14290 2069 14348 2075
rect 14290 2066 14302 2069
rect 13968 2038 14302 2066
rect 13968 2035 13980 2038
rect 13922 2029 13980 2035
rect 14290 2035 14302 2038
rect 14336 2066 14348 2069
rect 14662 2069 14720 2075
rect 14662 2066 14674 2069
rect 14336 2038 14674 2066
rect 14336 2035 14348 2038
rect 14290 2029 14348 2035
rect 14662 2035 14674 2038
rect 14708 2066 14720 2069
rect 14938 2069 14996 2075
rect 14938 2066 14950 2069
rect 14708 2038 14950 2066
rect 14708 2035 14720 2038
rect 14662 2029 14720 2035
rect 14938 2035 14950 2038
rect 14984 2035 14996 2069
rect 14938 2029 14996 2035
rect 15986 2069 16044 2075
rect 15986 2035 15998 2069
rect 16032 2066 16044 2069
rect 16072 2066 16100 2242
rect 16170 2137 16228 2143
rect 16170 2103 16182 2137
rect 16216 2134 16228 2137
rect 16910 2137 16968 2143
rect 16910 2134 16922 2137
rect 16216 2106 16922 2134
rect 16216 2103 16228 2106
rect 16170 2097 16228 2103
rect 16910 2103 16922 2106
rect 16956 2103 16968 2137
rect 16910 2097 16968 2103
rect 16354 2069 16412 2075
rect 16354 2066 16366 2069
rect 16032 2038 16366 2066
rect 16032 2035 16044 2038
rect 15986 2029 16044 2035
rect 16354 2035 16366 2038
rect 16400 2066 16412 2069
rect 16726 2069 16784 2075
rect 16726 2066 16738 2069
rect 16400 2038 16738 2066
rect 16400 2035 16412 2038
rect 16354 2029 16412 2035
rect 16726 2035 16738 2038
rect 16772 2066 16784 2069
rect 17002 2069 17060 2075
rect 17002 2066 17014 2069
rect 16772 2038 17014 2066
rect 16772 2035 16784 2038
rect 16726 2029 16784 2035
rect 17002 2035 17014 2038
rect 17048 2035 17060 2069
rect 17002 2029 17060 2035
rect 7040 2023 7098 2029
rect 2094 1999 2152 2005
rect 2094 1965 2106 1999
rect 2140 1996 2152 1999
rect 2554 1999 2612 2005
rect 2554 1996 2566 1999
rect 2140 1968 2566 1996
rect 2140 1965 2152 1968
rect 2094 1959 2152 1965
rect 2554 1965 2566 1968
rect 2600 1996 2612 1999
rect 2926 1999 2984 2005
rect 8118 2001 8176 2007
rect 2926 1996 2938 1999
rect 2600 1968 2938 1996
rect 2600 1965 2612 1968
rect 2554 1959 2612 1965
rect 2192 1938 2258 1940
rect 2192 1886 2198 1938
rect 2250 1886 2258 1938
rect 2192 1882 2258 1886
rect 2648 1792 2676 1968
rect 2926 1965 2938 1968
rect 2972 1965 2984 1999
rect 2926 1959 2984 1965
rect 4164 1995 4222 2001
rect 4164 1961 4176 1995
rect 4210 1992 4222 1995
rect 4624 1995 4682 2001
rect 4624 1992 4636 1995
rect 4210 1964 4636 1992
rect 4210 1961 4222 1964
rect 4164 1955 4222 1961
rect 4624 1961 4636 1964
rect 4670 1992 4682 1995
rect 4996 1995 5054 2001
rect 4996 1992 5008 1995
rect 4670 1964 5008 1992
rect 4670 1961 4682 1964
rect 4624 1955 4682 1961
rect 3200 1926 3260 1950
rect 3200 1890 3214 1926
rect 3254 1924 3260 1926
rect 4260 1928 4320 1934
rect 4260 1924 4274 1928
rect 3254 1894 4274 1924
rect 4308 1894 4320 1928
rect 3254 1890 4320 1894
rect 3200 1886 4320 1890
rect 3200 1874 3260 1886
rect 4260 1872 4320 1886
rect 1806 1778 3278 1792
rect 4718 1788 4746 1964
rect 4996 1961 5008 1964
rect 5042 1961 5054 1995
rect 4996 1955 5054 1961
rect 6116 1995 6174 2001
rect 6116 1961 6128 1995
rect 6162 1992 6174 1995
rect 6576 1995 6634 2001
rect 6576 1992 6588 1995
rect 6162 1964 6588 1992
rect 6162 1961 6174 1964
rect 6116 1955 6174 1961
rect 6576 1961 6588 1964
rect 6622 1992 6634 1995
rect 6948 1995 7006 2001
rect 6948 1992 6960 1995
rect 6622 1964 6960 1992
rect 6622 1961 6634 1964
rect 6576 1955 6634 1961
rect 5278 1922 5330 1940
rect 6212 1928 6272 1934
rect 6212 1924 6226 1928
rect 5518 1922 6226 1924
rect 5276 1886 5290 1922
rect 5324 1894 6226 1922
rect 6260 1894 6272 1928
rect 5324 1886 6272 1894
rect 5276 1884 5565 1886
rect 5278 1874 5330 1884
rect 6212 1872 6272 1886
rect 6670 1788 6698 1964
rect 6948 1961 6960 1964
rect 6994 1961 7006 1995
rect 8118 1967 8130 2001
rect 8164 1998 8176 2001
rect 8578 2001 8636 2007
rect 8578 1998 8590 2001
rect 8164 1970 8590 1998
rect 8164 1967 8176 1970
rect 8118 1961 8176 1967
rect 8578 1967 8590 1970
rect 8624 1998 8636 2001
rect 8950 2001 9008 2007
rect 8950 1998 8962 2001
rect 8624 1970 8962 1998
rect 8624 1967 8636 1970
rect 8578 1961 8636 1967
rect 6948 1955 7006 1961
rect 7230 1922 7282 1940
rect 8214 1934 8274 1940
rect 8214 1930 8228 1934
rect 7456 1922 8228 1930
rect 7228 1886 7242 1922
rect 7276 1900 8228 1922
rect 8262 1900 8274 1934
rect 7276 1892 8274 1900
rect 7276 1886 7517 1892
rect 7228 1884 7517 1886
rect 7230 1874 7282 1884
rect 8214 1878 8274 1892
rect 8672 1794 8700 1970
rect 8950 1967 8962 1970
rect 8996 1967 9008 2001
rect 8950 1961 9008 1967
rect 10070 2001 10128 2007
rect 10070 1967 10082 2001
rect 10116 1998 10128 2001
rect 10530 2001 10588 2007
rect 10530 1998 10542 2001
rect 10116 1970 10542 1998
rect 10116 1967 10128 1970
rect 10070 1961 10128 1967
rect 10530 1967 10542 1970
rect 10576 1998 10588 2001
rect 10902 2001 10960 2007
rect 10902 1998 10914 2001
rect 10576 1970 10914 1998
rect 10576 1967 10588 1970
rect 10530 1961 10588 1967
rect 9232 1928 9284 1946
rect 10166 1934 10226 1940
rect 10166 1930 10180 1934
rect 9472 1928 10180 1930
rect 9230 1892 9244 1928
rect 9278 1900 10180 1928
rect 10214 1900 10226 1934
rect 9278 1892 10226 1900
rect 9230 1890 9519 1892
rect 9232 1880 9284 1890
rect 10166 1878 10226 1892
rect 10624 1794 10652 1970
rect 10902 1967 10914 1970
rect 10948 1967 10960 2001
rect 10902 1961 10960 1967
rect 12062 2001 12120 2007
rect 12062 1967 12074 2001
rect 12108 1998 12120 2001
rect 12522 2001 12580 2007
rect 12522 1998 12534 2001
rect 12108 1970 12534 1998
rect 12108 1967 12120 1970
rect 12062 1961 12120 1967
rect 12522 1967 12534 1970
rect 12568 1998 12580 2001
rect 12894 2001 12952 2007
rect 12894 1998 12906 2001
rect 12568 1970 12906 1998
rect 12568 1967 12580 1970
rect 12522 1961 12580 1967
rect 11184 1928 11236 1946
rect 12158 1934 12218 1940
rect 12158 1930 12172 1934
rect 11317 1928 12172 1930
rect 11182 1892 11196 1928
rect 11230 1900 12172 1928
rect 12206 1900 12218 1934
rect 11230 1892 12218 1900
rect 11182 1890 11382 1892
rect 11184 1880 11236 1890
rect 12158 1878 12218 1892
rect 12616 1794 12644 1970
rect 12894 1967 12906 1970
rect 12940 1967 12952 2001
rect 12894 1961 12952 1967
rect 14014 2001 14072 2007
rect 14014 1967 14026 2001
rect 14060 1998 14072 2001
rect 14474 2001 14532 2007
rect 14474 1998 14486 2001
rect 14060 1970 14486 1998
rect 14060 1967 14072 1970
rect 14014 1961 14072 1967
rect 14474 1967 14486 1970
rect 14520 1998 14532 2001
rect 14846 2001 14904 2007
rect 14846 1998 14858 2001
rect 14520 1970 14858 1998
rect 14520 1967 14532 1970
rect 14474 1961 14532 1967
rect 13176 1928 13228 1946
rect 14110 1934 14170 1940
rect 14110 1930 14124 1934
rect 13416 1928 14124 1930
rect 13174 1892 13188 1928
rect 13222 1900 14124 1928
rect 14158 1900 14170 1934
rect 13222 1892 14170 1900
rect 13174 1890 13463 1892
rect 13176 1880 13228 1890
rect 14110 1878 14170 1892
rect 14568 1794 14596 1970
rect 14846 1967 14858 1970
rect 14892 1967 14904 2001
rect 14846 1961 14904 1967
rect 16078 2001 16136 2007
rect 16078 1967 16090 2001
rect 16124 1998 16136 2001
rect 16538 2001 16596 2007
rect 16538 1998 16550 2001
rect 16124 1970 16550 1998
rect 16124 1967 16136 1970
rect 16078 1961 16136 1967
rect 16538 1967 16550 1970
rect 16584 1998 16596 2001
rect 16910 2001 16968 2007
rect 16910 1998 16922 2001
rect 16584 1970 16922 1998
rect 16584 1967 16596 1970
rect 16538 1961 16596 1967
rect 15128 1928 15180 1946
rect 16174 1934 16234 1940
rect 16174 1930 16188 1934
rect 15538 1928 16188 1930
rect 15126 1892 15140 1928
rect 15174 1900 16188 1928
rect 16222 1900 16234 1934
rect 15174 1892 16234 1900
rect 15126 1890 15575 1892
rect 15128 1880 15180 1890
rect 16174 1878 16234 1892
rect 16632 1794 16660 1970
rect 16910 1967 16922 1970
rect 16956 1967 16968 2001
rect 16910 1961 16968 1967
rect 17192 1928 17244 1946
rect 17362 1930 17488 1982
rect 17362 1928 17402 1930
rect 17190 1892 17204 1928
rect 17238 1892 17402 1928
rect 17190 1890 17402 1892
rect 17192 1880 17244 1890
rect 17362 1876 17402 1890
rect 17454 1876 17488 1930
rect 17362 1828 17488 1876
rect 1806 1761 2604 1778
rect 2656 1761 3278 1778
rect 1806 1727 1835 1761
rect 1869 1727 1927 1761
rect 1961 1727 2019 1761
rect 2053 1727 2111 1761
rect 2145 1727 2203 1761
rect 2237 1727 2295 1761
rect 2329 1727 2387 1761
rect 2421 1727 2479 1761
rect 2513 1727 2571 1761
rect 2656 1727 2663 1761
rect 2697 1727 2755 1761
rect 2789 1727 2847 1761
rect 2881 1727 2939 1761
rect 2973 1727 3031 1761
rect 3065 1727 3123 1761
rect 3157 1727 3215 1761
rect 3249 1727 3278 1761
rect 1806 1720 2604 1727
rect 2656 1720 3278 1727
rect 1806 1696 3278 1720
rect 3876 1768 5348 1788
rect 3876 1757 4596 1768
rect 4652 1757 5348 1768
rect 3876 1723 3905 1757
rect 3939 1723 3997 1757
rect 4031 1723 4089 1757
rect 4123 1723 4181 1757
rect 4215 1723 4273 1757
rect 4307 1723 4365 1757
rect 4399 1723 4457 1757
rect 4491 1723 4549 1757
rect 4583 1723 4596 1757
rect 4675 1723 4733 1757
rect 4767 1723 4825 1757
rect 4859 1723 4917 1757
rect 4951 1723 5009 1757
rect 5043 1723 5101 1757
rect 5135 1723 5193 1757
rect 5227 1723 5285 1757
rect 5319 1723 5348 1757
rect 3876 1710 4596 1723
rect 4652 1710 5348 1723
rect 3876 1692 5348 1710
rect 5828 1768 7300 1788
rect 5828 1757 6548 1768
rect 6604 1757 7300 1768
rect 5828 1723 5857 1757
rect 5891 1723 5949 1757
rect 5983 1723 6041 1757
rect 6075 1723 6133 1757
rect 6167 1723 6225 1757
rect 6259 1723 6317 1757
rect 6351 1723 6409 1757
rect 6443 1723 6501 1757
rect 6535 1723 6548 1757
rect 6627 1723 6685 1757
rect 6719 1723 6777 1757
rect 6811 1723 6869 1757
rect 6903 1723 6961 1757
rect 6995 1723 7053 1757
rect 7087 1723 7145 1757
rect 7179 1723 7237 1757
rect 7271 1723 7300 1757
rect 5828 1710 6548 1723
rect 6604 1710 7300 1723
rect 5828 1692 7300 1710
rect 7830 1774 9302 1794
rect 7830 1763 8550 1774
rect 8606 1763 9302 1774
rect 7830 1729 7859 1763
rect 7893 1729 7951 1763
rect 7985 1729 8043 1763
rect 8077 1729 8135 1763
rect 8169 1729 8227 1763
rect 8261 1729 8319 1763
rect 8353 1729 8411 1763
rect 8445 1729 8503 1763
rect 8537 1729 8550 1763
rect 8629 1729 8687 1763
rect 8721 1729 8779 1763
rect 8813 1729 8871 1763
rect 8905 1729 8963 1763
rect 8997 1729 9055 1763
rect 9089 1729 9147 1763
rect 9181 1729 9239 1763
rect 9273 1729 9302 1763
rect 7830 1716 8550 1729
rect 8606 1716 9302 1729
rect 7830 1698 9302 1716
rect 9782 1774 11254 1794
rect 9782 1763 10502 1774
rect 10558 1763 11254 1774
rect 9782 1729 9811 1763
rect 9845 1729 9903 1763
rect 9937 1729 9995 1763
rect 10029 1729 10087 1763
rect 10121 1729 10179 1763
rect 10213 1729 10271 1763
rect 10305 1729 10363 1763
rect 10397 1729 10455 1763
rect 10489 1729 10502 1763
rect 10581 1729 10639 1763
rect 10673 1729 10731 1763
rect 10765 1729 10823 1763
rect 10857 1729 10915 1763
rect 10949 1729 11007 1763
rect 11041 1729 11099 1763
rect 11133 1729 11191 1763
rect 11225 1729 11254 1763
rect 9782 1716 10502 1729
rect 10558 1716 11254 1729
rect 9782 1698 11254 1716
rect 11774 1774 13246 1794
rect 11774 1763 12494 1774
rect 12550 1763 13246 1774
rect 11774 1729 11803 1763
rect 11837 1729 11895 1763
rect 11929 1729 11987 1763
rect 12021 1729 12079 1763
rect 12113 1729 12171 1763
rect 12205 1729 12263 1763
rect 12297 1729 12355 1763
rect 12389 1729 12447 1763
rect 12481 1729 12494 1763
rect 12573 1729 12631 1763
rect 12665 1729 12723 1763
rect 12757 1729 12815 1763
rect 12849 1729 12907 1763
rect 12941 1729 12999 1763
rect 13033 1729 13091 1763
rect 13125 1729 13183 1763
rect 13217 1729 13246 1763
rect 11774 1716 12494 1729
rect 12550 1716 13246 1729
rect 11774 1698 13246 1716
rect 13726 1774 15198 1794
rect 13726 1763 14446 1774
rect 14502 1763 15198 1774
rect 13726 1729 13755 1763
rect 13789 1729 13847 1763
rect 13881 1729 13939 1763
rect 13973 1729 14031 1763
rect 14065 1729 14123 1763
rect 14157 1729 14215 1763
rect 14249 1729 14307 1763
rect 14341 1729 14399 1763
rect 14433 1729 14446 1763
rect 14525 1729 14583 1763
rect 14617 1729 14675 1763
rect 14709 1729 14767 1763
rect 14801 1729 14859 1763
rect 14893 1729 14951 1763
rect 14985 1729 15043 1763
rect 15077 1729 15135 1763
rect 15169 1729 15198 1763
rect 13726 1716 14446 1729
rect 14502 1716 15198 1729
rect 13726 1698 15198 1716
rect 15790 1774 17262 1794
rect 15790 1763 16510 1774
rect 16566 1763 17262 1774
rect 15790 1729 15819 1763
rect 15853 1729 15911 1763
rect 15945 1729 16003 1763
rect 16037 1729 16095 1763
rect 16129 1729 16187 1763
rect 16221 1729 16279 1763
rect 16313 1729 16371 1763
rect 16405 1729 16463 1763
rect 16497 1729 16510 1763
rect 16589 1729 16647 1763
rect 16681 1729 16739 1763
rect 16773 1729 16831 1763
rect 16865 1729 16923 1763
rect 16957 1729 17015 1763
rect 17049 1729 17107 1763
rect 17141 1729 17199 1763
rect 17233 1729 17262 1763
rect 15790 1716 16510 1729
rect 16566 1716 17262 1729
rect 15790 1698 17262 1716
rect 30368 862 30432 5710
rect 30230 820 30542 862
rect 30230 716 30332 820
rect 30436 716 30542 820
rect 30230 638 30542 716
<< via1 >>
rect 9540 17762 9600 17822
rect 6646 17504 6722 17576
rect 9536 17218 9594 17278
rect 11414 16986 11474 17042
rect 4590 16570 4642 16624
rect 4976 16020 5034 16074
rect 4746 15814 4808 15874
rect 6712 15706 6780 15768
rect 6608 15356 6660 15408
rect 4898 15270 4966 15332
rect 6130 15202 6198 15264
rect 7114 15156 7182 15218
rect 4582 14986 4648 15052
rect 5794 14654 5862 14716
rect 5012 14442 5078 14508
rect 4682 14244 4754 14314
rect 6350 14232 6418 14294
rect 7916 14222 7984 14284
rect 9456 16607 9508 16628
rect 9456 16574 9489 16607
rect 9489 16574 9508 16607
rect 10872 16344 10942 16410
rect 9842 16063 9900 16078
rect 9842 16029 9857 16063
rect 9857 16029 9900 16063
rect 9842 16024 9900 16029
rect 9612 15863 9674 15878
rect 9612 15829 9645 15863
rect 9645 15829 9674 15863
rect 9612 15818 9674 15829
rect 11578 15753 11646 15772
rect 11578 15719 11595 15753
rect 11595 15719 11629 15753
rect 11629 15719 11646 15753
rect 11578 15710 11646 15719
rect 9842 15494 9896 15506
rect 9842 15460 9872 15494
rect 9872 15460 9896 15494
rect 9842 15452 9896 15460
rect 9764 15319 9832 15336
rect 9764 15285 9771 15319
rect 9771 15285 9829 15319
rect 9829 15285 9832 15319
rect 9764 15274 9832 15285
rect 9448 15043 9514 15056
rect 9448 15009 9465 15043
rect 9465 15009 9499 15043
rect 9499 15009 9514 15043
rect 9448 14990 9514 15009
rect 11474 15404 11526 15412
rect 11474 15368 11498 15404
rect 11498 15368 11526 15404
rect 11474 15360 11526 15368
rect 10996 15253 11064 15268
rect 10996 15219 11013 15253
rect 11013 15219 11047 15253
rect 11047 15219 11064 15253
rect 10996 15206 11064 15219
rect 11980 15209 12048 15222
rect 11980 15175 11997 15209
rect 11997 15175 12048 15209
rect 11980 15160 12048 15175
rect 9878 14499 9944 14512
rect 9878 14465 9925 14499
rect 9925 14465 9944 14499
rect 9878 14446 9944 14465
rect 9548 14299 9620 14318
rect 9548 14265 9563 14299
rect 9563 14265 9597 14299
rect 9597 14265 9620 14299
rect 9548 14248 9620 14265
rect 6828 13856 6896 13918
rect 7652 13882 7704 13936
rect 9896 13842 9956 13904
rect 4884 13700 4956 13770
rect 9750 13755 9822 13774
rect 5862 13692 5930 13754
rect 7656 13676 7724 13738
rect 9750 13721 9781 13755
rect 9781 13721 9822 13755
rect 9750 13704 9822 13721
rect 5984 13390 6052 13450
rect 4576 13318 4648 13384
rect 7136 13316 7204 13378
rect 9442 13375 9514 13388
rect 9442 13341 9457 13375
rect 9457 13341 9491 13375
rect 9491 13341 9514 13375
rect 9442 13322 9514 13341
rect 10660 14709 10728 14720
rect 10660 14675 10679 14709
rect 10679 14675 10728 14709
rect 10660 14658 10728 14675
rect 11216 14287 11284 14298
rect 11216 14253 11271 14287
rect 11271 14253 11284 14287
rect 11216 14236 11284 14253
rect 16430 16660 16498 16722
rect 17188 16652 17256 16714
rect 18078 16654 18146 16716
rect 18686 16650 18754 16712
rect 19444 16642 19512 16704
rect 20334 16644 20402 16706
rect 21450 16644 21518 16706
rect 22208 16636 22276 16698
rect 23098 16638 23166 16700
rect 16410 16122 16478 16184
rect 17196 16112 17264 16174
rect 18076 16112 18144 16174
rect 18666 16112 18734 16174
rect 19452 16102 19520 16164
rect 20332 16102 20400 16164
rect 21430 16106 21498 16168
rect 22216 16096 22284 16158
rect 23096 16096 23164 16158
rect 24400 14810 24462 14870
rect 24144 14662 24196 14714
rect 12782 14271 12850 14288
rect 12782 14237 12801 14271
rect 12801 14237 12835 14271
rect 12835 14237 12850 14271
rect 12782 14226 12850 14237
rect 24452 14552 24504 14564
rect 24452 14518 24456 14552
rect 24456 14518 24492 14552
rect 24492 14518 24504 14552
rect 24452 14512 24504 14518
rect 24552 14554 24556 14578
rect 24556 14554 24592 14578
rect 24592 14554 24604 14578
rect 24552 14526 24604 14554
rect 24698 14528 24712 14536
rect 24712 14528 24746 14536
rect 24746 14528 24750 14536
rect 24698 14484 24750 14528
rect 23992 14258 24054 14318
rect 10164 13308 10226 13360
rect 10878 13884 10930 13894
rect 10878 13850 10886 13884
rect 10886 13850 10920 13884
rect 10920 13850 10930 13884
rect 10878 13842 10930 13850
rect 10976 13924 11028 13934
rect 10976 13890 10984 13924
rect 10984 13890 11018 13924
rect 11018 13890 11028 13924
rect 10976 13882 11028 13890
rect 11074 13834 11126 13890
rect 11694 13913 11762 13922
rect 11694 13879 11723 13913
rect 11723 13879 11762 13913
rect 11694 13860 11762 13879
rect 12518 13886 12570 13940
rect 12732 13964 12812 13984
rect 12732 13922 12746 13964
rect 12746 13922 12796 13964
rect 12796 13922 12812 13964
rect 12732 13908 12812 13922
rect 10728 13743 10796 13758
rect 10728 13709 10753 13743
rect 10753 13709 10796 13743
rect 10728 13696 10796 13709
rect 12522 13680 12590 13742
rect 10850 13445 10918 13454
rect 10850 13411 10877 13445
rect 10877 13411 10918 13445
rect 10850 13394 10918 13411
rect 11006 13338 11060 13342
rect 11006 13302 11012 13338
rect 11012 13302 11048 13338
rect 11048 13302 11060 13338
rect 11006 13290 11060 13302
rect 12002 13369 12070 13382
rect 12002 13335 12057 13369
rect 12057 13335 12070 13369
rect 12002 13320 12070 13335
rect 5996 12856 6064 12916
rect 11062 13070 11114 13086
rect 11062 13036 11098 13070
rect 11098 13036 11114 13070
rect 11062 13032 11114 13036
rect 4990 12778 5062 12844
rect 9856 12831 9928 12848
rect 9856 12797 9859 12831
rect 9859 12797 9917 12831
rect 9917 12797 9928 12831
rect 9856 12782 9928 12797
rect 4634 12576 4708 12642
rect 9500 12631 9574 12646
rect 9500 12597 9555 12631
rect 9555 12597 9574 12631
rect 9500 12580 9574 12597
rect 6280 12370 6348 12432
rect 9872 12326 9934 12394
rect 10862 12901 10930 12920
rect 10862 12867 10877 12901
rect 10877 12867 10930 12901
rect 10862 12860 10930 12867
rect 11146 12425 11214 12436
rect 11146 12391 11149 12425
rect 11149 12391 11207 12425
rect 11207 12391 11214 12425
rect 11146 12374 11214 12391
rect 11206 12200 11258 12212
rect 11206 12166 11212 12200
rect 11212 12166 11246 12200
rect 11246 12166 11258 12200
rect 11206 12160 11258 12166
rect 4906 12034 4980 12100
rect 9772 12087 9846 12104
rect 9772 12053 9773 12087
rect 9773 12053 9831 12087
rect 9831 12053 9846 12087
rect 9772 12038 9846 12053
rect 11016 12114 11068 12122
rect 11016 12080 11024 12114
rect 11024 12080 11060 12114
rect 11060 12080 11068 12114
rect 11016 12070 11068 12080
rect 6002 11830 6070 11892
rect 4560 11756 4640 11820
rect 9426 11811 9506 11824
rect 9426 11777 9467 11811
rect 9467 11777 9501 11811
rect 9501 11777 9506 11811
rect 9426 11760 9506 11777
rect 10868 11881 10936 11896
rect 10868 11847 10873 11881
rect 10873 11847 10931 11881
rect 10931 11847 10936 11881
rect 10868 11834 10936 11847
rect 4994 11214 5074 11278
rect 9860 11267 9940 11282
rect 9860 11233 9869 11267
rect 9869 11233 9927 11267
rect 9927 11233 9940 11267
rect 9860 11218 9940 11233
rect 4626 11010 4706 11074
rect 9492 11067 9572 11078
rect 9492 11033 9507 11067
rect 9507 11033 9565 11067
rect 9565 11033 9572 11067
rect 9492 11014 9572 11033
rect 5054 10676 5108 10732
rect 9920 10680 9974 10736
rect 4904 10476 4984 10540
rect 9770 10523 9850 10544
rect 9770 10489 9783 10523
rect 9783 10489 9841 10523
rect 9841 10489 9850 10523
rect 9770 10480 9850 10489
rect 6226 6617 6282 6638
rect 6226 6583 6233 6617
rect 6233 6583 6267 6617
rect 6267 6583 6282 6617
rect 6226 6580 6282 6583
rect 6168 6382 6220 6390
rect 6168 6348 6178 6382
rect 6178 6348 6212 6382
rect 6212 6348 6220 6382
rect 6168 6338 6220 6348
rect 6268 6384 6320 6396
rect 6268 6350 6274 6384
rect 6274 6350 6308 6384
rect 6308 6350 6320 6384
rect 6268 6344 6320 6350
rect 6170 6073 6226 6088
rect 6170 6039 6175 6073
rect 6175 6039 6226 6073
rect 6170 6030 6226 6039
rect 10406 5985 10464 6002
rect 10774 5985 10832 6000
rect 10406 5951 10415 5985
rect 10415 5951 10449 5985
rect 10449 5951 10464 5985
rect 10774 5951 10783 5985
rect 10783 5951 10817 5985
rect 10817 5951 10832 5985
rect 10406 5940 10464 5951
rect 10774 5936 10832 5951
rect 12796 5973 12852 5986
rect 12796 5939 12845 5973
rect 12845 5939 12852 5973
rect 12796 5928 12852 5939
rect 14754 5981 14810 5994
rect 14754 5947 14803 5981
rect 14803 5947 14810 5981
rect 14754 5936 14810 5947
rect 16748 5987 16804 6000
rect 16748 5953 16797 5987
rect 16797 5953 16804 5987
rect 16748 5942 16804 5953
rect 2564 5565 2620 5578
rect 2564 5531 2601 5565
rect 2601 5531 2620 5565
rect 2564 5520 2620 5531
rect 4686 5557 4742 5570
rect 4686 5523 4735 5557
rect 4735 5523 4742 5557
rect 4686 5512 4742 5523
rect 6638 5557 6694 5570
rect 6638 5523 6687 5557
rect 6687 5523 6694 5557
rect 6638 5512 6694 5523
rect 8640 5563 8696 5576
rect 8640 5529 8689 5563
rect 8689 5529 8696 5563
rect 10410 5614 10462 5618
rect 10410 5580 10418 5614
rect 10418 5580 10452 5614
rect 10452 5580 10462 5614
rect 10410 5566 10462 5580
rect 8640 5518 8696 5529
rect 11214 5441 11270 5452
rect 11214 5407 11243 5441
rect 11243 5407 11270 5441
rect 11214 5394 11270 5407
rect 12800 5429 12856 5440
rect 12800 5395 12845 5429
rect 12845 5395 12856 5429
rect 12800 5382 12856 5395
rect 14758 5437 14814 5448
rect 14758 5403 14803 5437
rect 14803 5403 14814 5437
rect 14758 5390 14814 5403
rect 16752 5443 16808 5454
rect 16752 5409 16797 5443
rect 16797 5409 16808 5443
rect 16752 5396 16808 5409
rect 18726 5364 18784 5428
rect 2228 5194 2280 5198
rect 2228 5160 2236 5194
rect 2236 5160 2270 5194
rect 2270 5160 2280 5194
rect 2228 5146 2280 5160
rect 10188 5111 10244 5120
rect 10188 5077 10201 5111
rect 10201 5077 10244 5111
rect 10188 5062 10244 5077
rect 2584 5021 2640 5040
rect 2584 4987 2601 5021
rect 2601 4987 2635 5021
rect 2635 4987 2640 5021
rect 2584 4982 2640 4987
rect 4690 5013 4746 5024
rect 4690 4979 4735 5013
rect 4735 4979 4746 5013
rect 4690 4966 4746 4979
rect 6642 5013 6698 5024
rect 6642 4979 6687 5013
rect 6687 4979 6698 5013
rect 6642 4966 6698 4979
rect 13032 5067 13088 5080
rect 8644 5019 8700 5030
rect 8644 4985 8689 5019
rect 8689 4985 8700 5019
rect 8644 4972 8700 4985
rect 13032 5033 13081 5067
rect 13081 5033 13088 5067
rect 13032 5022 13088 5033
rect 15034 5061 15090 5074
rect 15034 5027 15083 5061
rect 15083 5027 15090 5061
rect 15034 5016 15090 5027
rect 10438 4740 10490 4744
rect 10438 4706 10446 4740
rect 10446 4706 10480 4740
rect 10480 4706 10490 4740
rect 10438 4692 10490 4706
rect 17056 5043 17112 5056
rect 17056 5009 17105 5043
rect 17105 5009 17112 5043
rect 17056 4998 17112 5009
rect 19056 5042 19108 5050
rect 19056 5004 19064 5042
rect 19064 5004 19102 5042
rect 19102 5004 19108 5042
rect 19056 4998 19108 5004
rect 10788 4567 10844 4580
rect 10440 4533 10443 4566
rect 10443 4533 10477 4566
rect 10477 4533 10492 4566
rect 10788 4533 10811 4567
rect 10811 4533 10844 4567
rect 10440 4512 10492 4533
rect 10788 4522 10844 4533
rect 13036 4523 13092 4534
rect 13036 4489 13081 4523
rect 13081 4489 13092 4523
rect 13036 4476 13092 4489
rect 18720 4816 18778 4880
rect 15038 4517 15094 4528
rect 15038 4483 15083 4517
rect 15083 4483 15094 4517
rect 15038 4470 15094 4483
rect 17060 4499 17116 4510
rect 17060 4465 17105 4499
rect 17105 4465 17116 4499
rect 17060 4452 17116 4465
rect 6194 3320 6254 3382
rect 6138 3122 6190 3130
rect 6138 3088 6148 3122
rect 6148 3088 6182 3122
rect 6182 3088 6190 3122
rect 6138 3078 6190 3088
rect 6238 3124 6290 3136
rect 6238 3090 6244 3124
rect 6244 3090 6278 3124
rect 6278 3090 6290 3124
rect 6238 3084 6290 3090
rect 6176 2766 6236 2828
rect 2604 2305 2660 2318
rect 2604 2271 2605 2305
rect 2605 2271 2660 2305
rect 2604 2260 2660 2271
rect 4592 2301 4648 2314
rect 4592 2267 4641 2301
rect 4641 2267 4648 2301
rect 4592 2256 4648 2267
rect 6544 2301 6600 2314
rect 6544 2267 6593 2301
rect 6593 2267 6600 2301
rect 6544 2256 6600 2267
rect 8546 2307 8602 2320
rect 8546 2273 8595 2307
rect 8595 2273 8602 2307
rect 8546 2262 8602 2273
rect 10498 2307 10554 2320
rect 10498 2273 10547 2307
rect 10547 2273 10554 2307
rect 10498 2262 10554 2273
rect 12490 2307 12546 2320
rect 12490 2273 12539 2307
rect 12539 2273 12546 2307
rect 12490 2262 12546 2273
rect 14442 2307 14498 2320
rect 14442 2273 14491 2307
rect 14491 2273 14498 2307
rect 14442 2262 14498 2273
rect 16506 2307 16562 2320
rect 16506 2273 16555 2307
rect 16555 2273 16562 2307
rect 16506 2262 16562 2273
rect 2198 1934 2250 1938
rect 2198 1900 2206 1934
rect 2206 1900 2240 1934
rect 2240 1900 2250 1934
rect 2198 1886 2250 1900
rect 17402 1876 17454 1930
rect 2604 1761 2656 1778
rect 2604 1727 2605 1761
rect 2605 1727 2656 1761
rect 2604 1720 2656 1727
rect 4596 1757 4652 1768
rect 4596 1723 4641 1757
rect 4641 1723 4652 1757
rect 4596 1710 4652 1723
rect 6548 1757 6604 1768
rect 6548 1723 6593 1757
rect 6593 1723 6604 1757
rect 6548 1710 6604 1723
rect 8550 1763 8606 1774
rect 8550 1729 8595 1763
rect 8595 1729 8606 1763
rect 8550 1716 8606 1729
rect 10502 1763 10558 1774
rect 10502 1729 10547 1763
rect 10547 1729 10558 1763
rect 10502 1716 10558 1729
rect 12494 1763 12550 1774
rect 12494 1729 12539 1763
rect 12539 1729 12550 1763
rect 12494 1716 12550 1729
rect 14446 1763 14502 1774
rect 14446 1729 14491 1763
rect 14491 1729 14502 1763
rect 14446 1716 14502 1729
rect 16510 1763 16566 1774
rect 16510 1729 16555 1763
rect 16555 1729 16566 1763
rect 16510 1716 16566 1729
rect 30332 716 30436 820
<< metal2 >>
rect 9430 17822 9706 17844
rect 9430 17762 9540 17822
rect 9600 17762 9706 17822
rect 9430 17746 9706 17762
rect 6463 17587 6545 17588
rect 6463 17586 6759 17587
rect 6463 17576 6760 17586
rect 6463 17505 6646 17576
rect 4472 16624 4732 16636
rect 4472 16614 4590 16624
rect 4472 16558 4552 16614
rect 4642 16570 4732 16624
rect 4608 16558 4732 16570
rect 4472 16536 4732 16558
rect 4886 16076 5106 16090
rect 4886 16020 4976 16076
rect 5034 16020 5106 16076
rect 4886 15994 5106 16020
rect 4562 15874 4938 15880
rect 4562 15814 4746 15874
rect 4808 15814 4938 15874
rect 4562 15792 4938 15814
rect 6463 15424 6545 17505
rect 6604 17504 6646 17505
rect 6722 17504 6760 17576
rect 6604 17498 6760 17504
rect 9432 17278 9706 17302
rect 9432 17218 9536 17278
rect 9594 17218 9706 17278
rect 9432 17202 9706 17218
rect 11401 17054 11483 17055
rect 11400 17042 11506 17054
rect 11400 16986 11414 17042
rect 11474 17033 11506 17042
rect 11474 16986 11507 17033
rect 11400 16812 11507 16986
rect 11329 16730 11507 16812
rect 9338 16628 9598 16640
rect 9338 16618 9456 16628
rect 9338 16562 9418 16618
rect 9508 16574 9598 16628
rect 9474 16562 9598 16574
rect 9338 16540 9598 16562
rect 10812 16410 11014 16442
rect 10812 16344 10872 16410
rect 10942 16344 11014 16410
rect 10812 16316 11014 16344
rect 9752 16080 9972 16094
rect 9752 16024 9842 16080
rect 9900 16024 9972 16080
rect 9752 15998 9972 16024
rect 9428 15878 9804 15884
rect 9428 15818 9612 15878
rect 9674 15818 9804 15878
rect 9428 15796 9804 15818
rect 6608 15768 6894 15780
rect 6608 15706 6712 15768
rect 6780 15706 6894 15768
rect 6608 15684 6894 15706
rect 9824 15506 9932 15514
rect 9824 15452 9842 15506
rect 9896 15476 9932 15506
rect 9896 15452 10324 15476
rect 9824 15440 10324 15452
rect 6463 15408 6682 15424
rect 6463 15356 6608 15408
rect 6660 15356 6682 15408
rect 4836 15332 5028 15350
rect 6463 15342 6682 15356
rect 4836 15270 4898 15332
rect 4966 15270 5028 15332
rect 9702 15336 9894 15354
rect 4836 15254 5028 15270
rect 6108 15264 6254 15280
rect 6108 15202 6130 15264
rect 6198 15202 6254 15264
rect 9702 15274 9764 15336
rect 9832 15274 9894 15336
rect 9702 15258 9894 15274
rect 6108 15184 6254 15202
rect 7046 15218 7252 15238
rect 7046 15156 7114 15218
rect 7182 15156 7252 15218
rect 7046 15140 7252 15156
rect 4476 15052 4750 15070
rect 4476 14986 4582 15052
rect 4648 14986 4750 15052
rect 4476 14978 4750 14986
rect 9342 15056 9616 15074
rect 9342 14990 9448 15056
rect 9514 14990 9616 15056
rect 9342 14982 9616 14990
rect 5748 14716 5908 14736
rect 5748 14654 5794 14716
rect 5862 14654 5908 14716
rect 5748 14640 5908 14654
rect 4946 14508 5118 14524
rect 4946 14442 5012 14508
rect 5078 14442 5118 14508
rect 4946 14434 5118 14442
rect 7635 14487 8531 14581
rect 4576 14314 4870 14320
rect 4576 14244 4682 14314
rect 4754 14244 4870 14314
rect 4576 14232 4870 14244
rect 6322 14294 6470 14316
rect 6322 14232 6350 14294
rect 6418 14232 6470 14294
rect 6322 14218 6470 14232
rect 7635 13974 7729 14487
rect 7840 14284 8072 14296
rect 7840 14222 7916 14284
rect 7984 14222 8072 14284
rect 7840 14204 8072 14222
rect 6794 13918 6946 13938
rect 6794 13856 6828 13918
rect 6896 13856 6946 13918
rect 7635 13936 7806 13974
rect 7635 13882 7652 13936
rect 7704 13882 7806 13936
rect 7635 13857 7806 13882
rect 7724 13856 7806 13857
rect 6794 13842 6946 13856
rect 4820 13770 5040 13780
rect 4820 13700 4884 13770
rect 4956 13700 5040 13770
rect 4820 13684 5040 13700
rect 5824 13754 5974 13770
rect 5824 13692 5862 13754
rect 5930 13692 5974 13754
rect 5824 13672 5974 13692
rect 7642 13738 7744 13754
rect 7642 13676 7656 13738
rect 7724 13676 7744 13738
rect 7642 13658 7744 13676
rect 5950 13450 6084 13470
rect 4468 13384 4738 13396
rect 4468 13318 4576 13384
rect 4648 13318 4738 13384
rect 5950 13390 5984 13450
rect 6052 13390 6084 13450
rect 5950 13378 6084 13390
rect 7096 13378 7248 13396
rect 4468 13310 4738 13318
rect 7096 13316 7136 13378
rect 7204 13316 7248 13378
rect 7096 13300 7248 13316
rect 5948 12916 6100 12928
rect 5948 12856 5996 12916
rect 6064 12856 6100 12916
rect 4922 12844 5112 12854
rect 4922 12778 4990 12844
rect 5062 12778 5112 12844
rect 5948 12834 6100 12856
rect 4922 12766 5112 12778
rect 4574 12642 4780 12654
rect 4574 12576 4634 12642
rect 4708 12576 4780 12642
rect 4574 12560 4780 12576
rect 6230 12432 6402 12452
rect 6230 12370 6280 12432
rect 6348 12370 6402 12432
rect 6230 12356 6402 12370
rect 4858 12100 5024 12116
rect 4858 12034 4906 12100
rect 4980 12034 5024 12100
rect 4858 12022 5024 12034
rect 5944 11892 6100 11908
rect 4510 11820 4690 11834
rect 4510 11756 4560 11820
rect 4640 11756 4690 11820
rect 5944 11830 6002 11892
rect 6070 11830 6100 11892
rect 5944 11812 6100 11830
rect 4510 11746 4690 11756
rect 4938 11278 5118 11292
rect 4938 11214 4994 11278
rect 5074 11214 5118 11278
rect 4938 11204 5118 11214
rect 4580 11074 4776 11092
rect 4580 11010 4626 11074
rect 4706 11010 4776 11074
rect 4580 10996 4776 11010
rect 8437 10762 8531 14487
rect 9812 14512 9984 14528
rect 9812 14446 9878 14512
rect 9944 14446 9984 14512
rect 9812 14438 9984 14446
rect 9442 14318 9736 14324
rect 9442 14248 9548 14318
rect 9620 14248 9736 14318
rect 9442 14236 9736 14248
rect 10288 14102 10324 15440
rect 10614 14720 10774 14740
rect 10614 14658 10660 14720
rect 10728 14658 10774 14720
rect 10614 14644 10774 14658
rect 10876 14514 10944 16316
rect 11329 15428 11411 16730
rect 16346 16722 16558 16738
rect 16346 16660 16430 16722
rect 16498 16660 16558 16722
rect 16346 16646 16558 16660
rect 17116 16714 17328 16732
rect 17116 16652 17188 16714
rect 17256 16652 17328 16714
rect 17116 16640 17328 16652
rect 18008 16716 18220 16732
rect 18008 16654 18078 16716
rect 18146 16654 18220 16716
rect 18008 16640 18220 16654
rect 18602 16712 18814 16728
rect 18602 16650 18686 16712
rect 18754 16650 18814 16712
rect 18602 16636 18814 16650
rect 19372 16704 19584 16722
rect 19372 16642 19444 16704
rect 19512 16642 19584 16704
rect 19372 16630 19584 16642
rect 20264 16706 20476 16722
rect 20264 16644 20334 16706
rect 20402 16644 20476 16706
rect 20264 16630 20476 16644
rect 21366 16706 21578 16722
rect 21366 16644 21450 16706
rect 21518 16644 21578 16706
rect 21366 16630 21578 16644
rect 22136 16698 22348 16716
rect 22136 16636 22208 16698
rect 22276 16636 22348 16698
rect 22136 16624 22348 16636
rect 23028 16700 23240 16716
rect 23028 16638 23098 16700
rect 23166 16638 23240 16700
rect 23028 16624 23240 16638
rect 16336 16184 16548 16194
rect 16336 16122 16410 16184
rect 16478 16122 16548 16184
rect 16336 16102 16548 16122
rect 17126 16174 17338 16186
rect 17126 16112 17196 16174
rect 17264 16112 17338 16174
rect 17126 16094 17338 16112
rect 17996 16174 18208 16186
rect 17996 16112 18076 16174
rect 18144 16112 18208 16174
rect 17996 16094 18208 16112
rect 18592 16174 18804 16184
rect 18592 16112 18666 16174
rect 18734 16112 18804 16174
rect 18592 16092 18804 16112
rect 19382 16164 19594 16176
rect 19382 16102 19452 16164
rect 19520 16102 19594 16164
rect 19382 16084 19594 16102
rect 20252 16164 20464 16176
rect 20252 16102 20332 16164
rect 20400 16102 20464 16164
rect 20252 16084 20464 16102
rect 21356 16168 21568 16178
rect 21356 16106 21430 16168
rect 21498 16106 21568 16168
rect 21356 16086 21568 16106
rect 22146 16158 22358 16170
rect 22146 16096 22216 16158
rect 22284 16096 22358 16158
rect 22146 16078 22358 16096
rect 23016 16158 23228 16170
rect 23016 16096 23096 16158
rect 23164 16096 23228 16158
rect 23016 16078 23228 16096
rect 11474 15772 11760 15784
rect 11474 15710 11578 15772
rect 11646 15710 11760 15772
rect 11474 15688 11760 15710
rect 11329 15412 11548 15428
rect 11329 15360 11474 15412
rect 11526 15360 11548 15412
rect 11329 15346 11548 15360
rect 10974 15268 11120 15284
rect 10974 15206 10996 15268
rect 11064 15206 11120 15268
rect 10974 15188 11120 15206
rect 11912 15222 12118 15242
rect 11912 15160 11980 15222
rect 12048 15160 12118 15222
rect 11912 15144 12118 15160
rect 24312 14870 24542 14880
rect 24312 14810 24400 14870
rect 24462 14810 24542 14870
rect 24312 14788 24542 14810
rect 26389 14843 27464 14921
rect 26389 14740 26467 14843
rect 26948 14766 27172 14794
rect 26389 14726 26466 14740
rect 24138 14714 26466 14726
rect 24138 14662 24144 14714
rect 24196 14662 26466 14714
rect 24138 14658 26466 14662
rect 10876 14446 11034 14514
rect 10288 14066 10898 14102
rect 10862 13940 10898 14066
rect 9834 13904 10004 13916
rect 9834 13842 9896 13904
rect 9956 13884 10004 13904
rect 10862 13894 10938 13940
rect 10862 13884 10878 13894
rect 9956 13842 10580 13884
rect 9834 13836 10580 13842
rect 10860 13842 10878 13884
rect 10930 13842 10938 13894
rect 10860 13836 10938 13842
rect 9834 13822 10004 13836
rect 9686 13774 9906 13784
rect 9686 13704 9750 13774
rect 9822 13704 9906 13774
rect 9686 13688 9906 13704
rect 10530 13596 10578 13836
rect 10868 13798 10938 13836
rect 10966 13934 11034 14446
rect 12501 14491 13397 14585
rect 11188 14298 11336 14320
rect 11188 14236 11216 14298
rect 11284 14236 11336 14298
rect 11188 14222 11336 14236
rect 10966 13882 10976 13934
rect 11028 13882 11034 13934
rect 10966 13796 11034 13882
rect 11067 13890 11141 13989
rect 12501 13978 12595 14491
rect 12706 14288 12938 14300
rect 12706 14226 12782 14288
rect 12850 14226 12938 14288
rect 12706 14208 12938 14226
rect 12704 13984 12842 13996
rect 11067 13834 11074 13890
rect 11126 13834 11141 13890
rect 11660 13922 11812 13942
rect 11660 13860 11694 13922
rect 11762 13860 11812 13922
rect 12501 13940 12672 13978
rect 12501 13886 12518 13940
rect 12570 13886 12672 13940
rect 12704 13908 12732 13984
rect 12812 13908 12842 13984
rect 12704 13894 12842 13908
rect 12501 13861 12672 13886
rect 12590 13860 12672 13861
rect 11660 13846 11812 13860
rect 11067 13805 11141 13834
rect 10690 13758 10840 13774
rect 10690 13696 10728 13758
rect 10796 13696 10840 13758
rect 11067 13731 11209 13805
rect 10690 13676 10840 13696
rect 10530 13548 11040 13596
rect 10816 13454 10950 13474
rect 9334 13388 9604 13400
rect 9334 13322 9442 13388
rect 9514 13322 9604 13388
rect 10816 13394 10850 13454
rect 10918 13394 10950 13454
rect 10816 13382 10950 13394
rect 10992 13376 11040 13548
rect 10226 13370 10632 13372
rect 9334 13314 9604 13322
rect 10156 13360 10632 13370
rect 10156 13308 10164 13360
rect 10226 13308 10632 13360
rect 10156 13300 10632 13308
rect 10560 13174 10632 13300
rect 10986 13342 11084 13376
rect 10986 13290 11006 13342
rect 11060 13290 11084 13342
rect 10986 13272 11084 13290
rect 11135 13176 11209 13731
rect 12508 13742 12610 13758
rect 12508 13680 12522 13742
rect 12590 13680 12610 13742
rect 12508 13662 12610 13680
rect 12724 13660 12792 13894
rect 12704 13658 12792 13660
rect 12644 13590 12792 13658
rect 11962 13382 12114 13400
rect 11962 13320 12002 13382
rect 12070 13320 12114 13382
rect 11962 13304 12114 13320
rect 11006 13174 11209 13176
rect 10560 13102 11209 13174
rect 11052 13086 11124 13102
rect 11052 13032 11062 13086
rect 11114 13032 11124 13086
rect 11052 12948 11124 13032
rect 10814 12920 10966 12932
rect 10814 12860 10862 12920
rect 10930 12860 10966 12920
rect 9788 12848 9978 12858
rect 9788 12782 9856 12848
rect 9928 12782 9978 12848
rect 10814 12838 10966 12860
rect 9788 12770 9978 12782
rect 9440 12646 9646 12658
rect 9440 12580 9500 12646
rect 9574 12580 9646 12646
rect 9440 12564 9646 12580
rect 11096 12436 11268 12456
rect 9826 12394 9976 12408
rect 9826 12326 9872 12394
rect 9934 12342 9976 12394
rect 11096 12374 11146 12436
rect 11214 12374 11268 12436
rect 11096 12360 11268 12374
rect 9934 12326 11056 12342
rect 9826 12310 11056 12326
rect 11024 12130 11056 12310
rect 12644 12222 12712 13590
rect 11200 12212 12712 12222
rect 11200 12160 11206 12212
rect 11258 12160 12712 12212
rect 11200 12154 12712 12160
rect 11008 12122 11078 12130
rect 9724 12104 9890 12120
rect 9724 12038 9772 12104
rect 9846 12038 9890 12104
rect 11008 12070 11016 12122
rect 11068 12070 11078 12122
rect 11008 12064 11078 12070
rect 9724 12026 9890 12038
rect 10810 11896 10966 11912
rect 9376 11824 9556 11838
rect 9376 11760 9426 11824
rect 9506 11760 9556 11824
rect 10810 11834 10868 11896
rect 10936 11834 10966 11896
rect 10810 11816 10966 11834
rect 9376 11750 9556 11760
rect 9804 11282 9984 11296
rect 9804 11218 9860 11282
rect 9940 11218 9984 11282
rect 9804 11208 9984 11218
rect 9446 11078 9642 11096
rect 9446 11014 9492 11078
rect 9572 11014 9642 11078
rect 9446 11000 9642 11014
rect 13303 10766 13397 14491
rect 24138 14488 24198 14658
rect 26389 14657 26466 14658
rect 26948 14646 27000 14766
rect 27122 14726 27172 14766
rect 27122 14658 27176 14726
rect 27122 14646 27172 14658
rect 24448 14564 24504 14620
rect 24448 14512 24452 14564
rect 23850 14318 24212 14334
rect 23850 14258 23992 14318
rect 24054 14258 24212 14318
rect 23850 14240 24212 14258
rect 24448 14112 24504 14512
rect 24546 14578 24606 14622
rect 24546 14526 24552 14578
rect 24604 14526 24606 14578
rect 24448 14056 24502 14112
rect 4970 10732 8531 10762
rect 4970 10676 5054 10732
rect 5108 10676 8531 10732
rect 4970 10668 8531 10676
rect 9836 10736 13397 10766
rect 9836 10680 9920 10736
rect 9974 10680 13397 10736
rect 9836 10672 13397 10680
rect 23258 14000 24502 14056
rect 4970 10652 5202 10668
rect 9836 10656 10068 10672
rect 4856 10540 5036 10546
rect 4856 10476 4904 10540
rect 4984 10476 5036 10540
rect 4856 10458 5036 10476
rect 9722 10544 9902 10550
rect 9722 10480 9770 10544
rect 9850 10480 9902 10544
rect 9722 10462 9902 10480
rect 6112 6638 6388 6648
rect 6112 6580 6226 6638
rect 6282 6580 6388 6638
rect 6112 6558 6388 6580
rect 5585 6398 5651 6404
rect 2222 6390 6228 6398
rect 2222 6338 6168 6390
rect 6220 6338 6228 6390
rect 6262 6396 13156 6398
rect 6262 6344 6268 6396
rect 6320 6394 13156 6396
rect 23258 6394 23314 14000
rect 24546 13290 24606 14526
rect 24684 14536 24776 14624
rect 26948 14604 27172 14646
rect 24684 14484 24698 14536
rect 24750 14514 24776 14536
rect 26993 14514 27071 14604
rect 24750 14484 27071 14514
rect 24684 14436 27071 14484
rect 27386 14514 27464 14843
rect 27386 14510 27604 14514
rect 27386 14492 27730 14510
rect 27386 14436 27550 14492
rect 27512 14372 27550 14436
rect 27682 14372 27730 14492
rect 27512 14336 27730 14372
rect 6320 6344 23314 6394
rect 6262 6340 23314 6344
rect 6262 6338 16050 6340
rect 17150 6338 23314 6340
rect 24252 13230 24608 13290
rect 2222 6332 6228 6338
rect 18793 6336 18848 6338
rect 2222 5198 2290 6332
rect 6110 6088 6274 6104
rect 6110 6030 6170 6088
rect 6226 6030 6274 6088
rect 6110 6018 6274 6030
rect 10404 6002 10472 6018
rect 10404 5940 10406 6002
rect 10464 5940 10472 6002
rect 10404 5618 10472 5940
rect 10708 6000 10888 6016
rect 10708 5936 10774 6000
rect 10832 5936 10888 6000
rect 10708 5922 10888 5936
rect 12738 5986 12918 6002
rect 12738 5928 12796 5986
rect 12852 5928 12918 5986
rect 12738 5908 12918 5928
rect 14696 5994 14876 6010
rect 14696 5936 14754 5994
rect 14810 5936 14876 5994
rect 14696 5916 14876 5936
rect 16690 6000 16870 6016
rect 16690 5942 16748 6000
rect 16804 5942 16870 6000
rect 16690 5922 16870 5942
rect 2510 5578 2690 5596
rect 2510 5520 2564 5578
rect 2620 5520 2690 5578
rect 2510 5502 2690 5520
rect 4628 5570 4808 5586
rect 4628 5512 4686 5570
rect 4742 5512 4808 5570
rect 4628 5492 4808 5512
rect 6580 5570 6760 5586
rect 6580 5512 6638 5570
rect 6694 5512 6760 5570
rect 6580 5492 6760 5512
rect 8582 5576 8762 5592
rect 8582 5518 8640 5576
rect 8696 5518 8762 5576
rect 10404 5566 10410 5618
rect 10462 5566 10472 5618
rect 10404 5562 10472 5566
rect 8582 5498 8762 5518
rect 11142 5452 11324 5474
rect 11142 5394 11214 5452
rect 11270 5394 11324 5452
rect 11142 5378 11324 5394
rect 12738 5440 12918 5458
rect 12738 5382 12800 5440
rect 12856 5382 12918 5440
rect 12738 5364 12918 5382
rect 14696 5448 14876 5466
rect 14696 5390 14758 5448
rect 14814 5390 14876 5448
rect 14696 5372 14876 5390
rect 16690 5454 16870 5472
rect 16690 5396 16752 5454
rect 16808 5396 16870 5454
rect 16690 5378 16870 5396
rect 18658 5428 18838 5444
rect 18658 5364 18726 5428
rect 18784 5364 18838 5428
rect 18658 5348 18838 5364
rect 2222 5146 2228 5198
rect 2280 5146 2290 5198
rect 19193 5175 19248 6338
rect 2222 5142 2290 5146
rect 10128 5120 10308 5142
rect 10128 5062 10188 5120
rect 10244 5062 10308 5120
rect 19196 5098 19244 5175
rect 2520 5040 2700 5050
rect 2520 4982 2584 5040
rect 2640 4982 2700 5040
rect 2520 4956 2700 4982
rect 4628 5024 4808 5042
rect 4628 4966 4690 5024
rect 4746 4966 4808 5024
rect 4628 4948 4808 4966
rect 6580 5024 6760 5042
rect 6580 4966 6642 5024
rect 6698 4966 6760 5024
rect 6580 4948 6760 4966
rect 8582 5030 8762 5048
rect 10128 5046 10308 5062
rect 12974 5080 13154 5096
rect 8582 4972 8644 5030
rect 8700 4972 8762 5030
rect 12974 5022 13032 5080
rect 13088 5022 13154 5080
rect 12974 5002 13154 5022
rect 14976 5074 15156 5090
rect 14976 5016 15034 5074
rect 15090 5016 15156 5074
rect 14976 4996 15156 5016
rect 16998 5056 17178 5072
rect 16998 4998 17056 5056
rect 17112 4998 17178 5056
rect 16998 4978 17178 4998
rect 19048 5050 19244 5098
rect 19048 4998 19056 5050
rect 19108 4998 19112 5050
rect 8582 4954 8762 4972
rect 19048 4942 19112 4998
rect 18662 4880 18842 4894
rect 18662 4816 18720 4880
rect 18778 4816 18842 4880
rect 10432 4744 10500 4802
rect 18662 4798 18842 4816
rect 10432 4692 10438 4744
rect 10490 4692 10500 4744
rect 10432 4566 10500 4692
rect 10432 4512 10440 4566
rect 10492 4512 10500 4566
rect 10432 4502 10500 4512
rect 10734 4580 10914 4594
rect 10734 4522 10788 4580
rect 10844 4522 10914 4580
rect 10734 4498 10914 4522
rect 12974 4534 13154 4552
rect 12974 4476 13036 4534
rect 13092 4476 13154 4534
rect 12974 4458 13154 4476
rect 14976 4528 15156 4546
rect 14976 4470 15038 4528
rect 15094 4470 15156 4528
rect 14976 4452 15156 4470
rect 16998 4510 17178 4528
rect 16998 4452 17060 4510
rect 17116 4452 17178 4510
rect 16998 4434 17178 4452
rect 6082 3382 6354 3386
rect 6082 3320 6194 3382
rect 6254 3320 6354 3382
rect 6082 3292 6354 3320
rect 24252 3138 24312 13230
rect 2192 3130 6198 3138
rect 2192 3078 6138 3130
rect 6190 3078 6198 3130
rect 6232 3136 24312 3138
rect 6232 3084 6238 3136
rect 6290 3084 24312 3136
rect 6232 3078 24312 3084
rect 2192 3072 6198 3078
rect 2192 1938 2260 3072
rect 6080 2828 6300 2842
rect 6080 2766 6176 2828
rect 6236 2766 6300 2828
rect 6080 2752 6300 2766
rect 2540 2318 2720 2336
rect 2540 2260 2604 2318
rect 2660 2260 2720 2318
rect 2540 2242 2720 2260
rect 4534 2314 4714 2330
rect 4534 2256 4592 2314
rect 4648 2256 4714 2314
rect 4534 2236 4714 2256
rect 6486 2314 6666 2330
rect 6486 2256 6544 2314
rect 6600 2256 6666 2314
rect 6486 2236 6666 2256
rect 8488 2320 8668 2336
rect 8488 2262 8546 2320
rect 8602 2262 8668 2320
rect 8488 2242 8668 2262
rect 10440 2320 10620 2336
rect 10440 2262 10498 2320
rect 10554 2262 10620 2320
rect 10440 2242 10620 2262
rect 12432 2320 12612 2336
rect 12432 2262 12490 2320
rect 12546 2262 12612 2320
rect 12432 2242 12612 2262
rect 14384 2320 14564 2336
rect 14384 2262 14442 2320
rect 14498 2262 14564 2320
rect 14384 2242 14564 2262
rect 16448 2320 16628 2336
rect 16448 2262 16506 2320
rect 16562 2262 16628 2320
rect 16448 2242 16628 2262
rect 17390 1982 17450 3078
rect 2192 1886 2198 1938
rect 2250 1886 2260 1938
rect 2192 1882 2260 1886
rect 17362 1930 17488 1982
rect 17362 1876 17402 1930
rect 17454 1876 17488 1930
rect 17362 1828 17488 1876
rect 2538 1778 2718 1794
rect 2538 1720 2604 1778
rect 2660 1720 2718 1778
rect 2538 1700 2718 1720
rect 4534 1768 4714 1786
rect 4534 1710 4596 1768
rect 4652 1710 4714 1768
rect 4534 1692 4714 1710
rect 6486 1768 6666 1786
rect 6486 1710 6548 1768
rect 6604 1710 6666 1768
rect 6486 1692 6666 1710
rect 8488 1774 8668 1792
rect 8488 1716 8550 1774
rect 8606 1716 8668 1774
rect 8488 1698 8668 1716
rect 10440 1774 10620 1792
rect 10440 1716 10502 1774
rect 10558 1716 10620 1774
rect 10440 1698 10620 1716
rect 12432 1774 12612 1792
rect 12432 1716 12494 1774
rect 12550 1716 12612 1774
rect 12432 1698 12612 1716
rect 14384 1774 14564 1792
rect 14384 1716 14446 1774
rect 14502 1716 14564 1774
rect 14384 1698 14564 1716
rect 16448 1774 16628 1792
rect 16448 1716 16510 1774
rect 16566 1716 16628 1774
rect 16448 1698 16628 1716
rect 30230 820 30542 862
rect 30230 716 30332 820
rect 30436 716 30542 820
rect 30230 638 30542 716
<< via2 >>
rect 9540 17762 9600 17822
rect 4552 16570 4590 16614
rect 4590 16570 4608 16614
rect 4552 16558 4608 16570
rect 4976 16074 5034 16076
rect 4976 16020 5034 16074
rect 4746 15814 4808 15874
rect 9536 17218 9594 17278
rect 9418 16574 9456 16618
rect 9456 16574 9474 16618
rect 9418 16562 9474 16574
rect 9842 16078 9900 16080
rect 9842 16024 9900 16078
rect 9612 15818 9674 15878
rect 6712 15706 6780 15768
rect 4898 15270 4966 15332
rect 6130 15202 6198 15264
rect 9764 15274 9832 15336
rect 7114 15156 7182 15218
rect 4582 14986 4648 15052
rect 9448 14990 9514 15056
rect 5794 14654 5862 14716
rect 5012 14442 5078 14508
rect 4682 14244 4754 14314
rect 6350 14232 6418 14294
rect 7916 14222 7984 14284
rect 6828 13856 6896 13918
rect 4884 13700 4956 13770
rect 5862 13692 5930 13754
rect 7656 13676 7724 13738
rect 4576 13318 4648 13384
rect 5984 13390 6052 13450
rect 7136 13316 7204 13378
rect 5996 12856 6064 12916
rect 4990 12778 5062 12844
rect 4634 12576 4708 12642
rect 6280 12370 6348 12432
rect 4906 12034 4980 12100
rect 4560 11756 4640 11820
rect 6002 11830 6070 11892
rect 4994 11214 5074 11278
rect 4626 11010 4706 11074
rect 9878 14446 9944 14512
rect 9548 14248 9620 14318
rect 10660 14658 10728 14720
rect 16430 16660 16498 16722
rect 17188 16652 17256 16714
rect 18078 16654 18146 16716
rect 18686 16650 18754 16712
rect 19444 16642 19512 16704
rect 20334 16644 20402 16706
rect 21450 16644 21518 16706
rect 22208 16636 22276 16698
rect 23098 16638 23166 16700
rect 16410 16122 16478 16184
rect 17196 16112 17264 16174
rect 18076 16112 18144 16174
rect 18666 16112 18734 16174
rect 19452 16102 19520 16164
rect 20332 16102 20400 16164
rect 21430 16106 21498 16168
rect 22216 16096 22284 16158
rect 23096 16096 23164 16158
rect 11578 15710 11646 15772
rect 10996 15206 11064 15268
rect 11980 15160 12048 15222
rect 24400 14810 24462 14870
rect 9750 13704 9822 13774
rect 11216 14236 11284 14298
rect 12782 14226 12850 14288
rect 11694 13860 11762 13922
rect 10728 13696 10796 13758
rect 9442 13322 9514 13388
rect 10850 13394 10918 13454
rect 12522 13680 12590 13742
rect 12002 13320 12070 13382
rect 10862 12860 10930 12920
rect 9856 12782 9928 12848
rect 9500 12580 9574 12646
rect 11146 12374 11214 12436
rect 9772 12038 9846 12104
rect 9426 11760 9506 11824
rect 10868 11834 10936 11896
rect 9860 11218 9940 11282
rect 9492 11014 9572 11078
rect 27000 14646 27122 14766
rect 23992 14258 24054 14318
rect 4904 10476 4984 10540
rect 9770 10480 9850 10544
rect 6226 6580 6282 6638
rect 27550 14372 27682 14492
rect 6170 6030 6226 6088
rect 10774 5936 10832 6000
rect 12796 5928 12852 5986
rect 14754 5936 14810 5994
rect 16748 5942 16804 6000
rect 2564 5520 2620 5578
rect 4686 5512 4742 5570
rect 6638 5512 6694 5570
rect 8640 5518 8696 5576
rect 11214 5394 11270 5452
rect 12800 5382 12856 5440
rect 14758 5390 14814 5448
rect 16752 5396 16808 5454
rect 18726 5364 18784 5428
rect 10188 5062 10244 5120
rect 2584 4982 2640 5040
rect 4690 4966 4746 5024
rect 6642 4966 6698 5024
rect 8644 4972 8700 5030
rect 13032 5022 13088 5080
rect 15034 5016 15090 5074
rect 17056 4998 17112 5056
rect 18720 4816 18778 4880
rect 10788 4522 10844 4580
rect 13036 4476 13092 4534
rect 15038 4470 15094 4528
rect 17060 4452 17116 4510
rect 6194 3320 6254 3382
rect 6176 2766 6236 2828
rect 2604 2260 2660 2318
rect 4592 2256 4648 2314
rect 6544 2256 6600 2314
rect 8546 2262 8602 2320
rect 10498 2262 10554 2320
rect 12490 2262 12546 2320
rect 14442 2262 14498 2320
rect 16506 2262 16562 2320
rect 2604 1720 2656 1778
rect 2656 1720 2660 1778
rect 4596 1710 4652 1768
rect 6548 1710 6604 1768
rect 8550 1716 8606 1774
rect 10502 1716 10558 1774
rect 12494 1716 12550 1774
rect 14446 1716 14502 1774
rect 16510 1716 16566 1774
rect 30332 716 30436 820
<< metal3 >>
rect 814 17848 23871 17936
rect 814 17780 996 17848
rect 1066 17822 23871 17848
rect 1066 17780 9540 17822
rect 814 17762 9540 17780
rect 9600 17762 23871 17822
rect 814 17722 23871 17762
rect 18799 17720 19013 17722
rect 200 17278 13306 17330
rect 200 17218 9536 17278
rect 9594 17218 13306 17278
rect 200 17104 13306 17218
rect 200 16942 322 17104
rect 474 17038 13306 17104
rect 474 17022 21152 17038
rect 474 16942 23276 17022
rect 200 16810 23276 16942
rect 200 16808 13306 16810
rect 4036 16628 4280 16808
rect 4036 16614 4844 16628
rect 4036 16558 4552 16614
rect 4608 16558 4844 16614
rect 4036 16536 4844 16558
rect 4036 15884 4280 16536
rect 4880 16076 5584 16082
rect 4880 16020 4976 16076
rect 5034 16020 5584 16076
rect 4880 15994 5584 16020
rect 5342 15912 5584 15994
rect 4036 15874 4938 15884
rect 4036 15814 4746 15874
rect 4808 15814 4938 15874
rect 4036 15792 4938 15814
rect 4036 15066 4280 15792
rect 5340 15344 5584 15912
rect 4834 15332 5584 15344
rect 4834 15270 4898 15332
rect 4966 15270 5584 15332
rect 6320 15780 6502 16808
rect 6320 15768 6896 15780
rect 6320 15706 6712 15768
rect 6780 15706 6896 15768
rect 6320 15684 6896 15706
rect 6320 15278 6502 15684
rect 4834 15256 5584 15270
rect 4036 15052 4900 15066
rect 4036 14986 4582 15052
rect 4648 14986 4900 15052
rect 4036 14974 4900 14986
rect 4036 14324 4280 14974
rect 5340 14738 5584 15256
rect 6088 15264 6502 15278
rect 6088 15202 6130 15264
rect 6198 15202 6502 15264
rect 6088 15180 6502 15202
rect 5340 14716 6026 14738
rect 5340 14654 5794 14716
rect 5862 14654 6026 14716
rect 5340 14642 6026 14654
rect 5340 14522 5584 14642
rect 4942 14508 5584 14522
rect 4942 14442 5012 14508
rect 5078 14442 5584 14508
rect 4942 14434 5584 14442
rect 4036 14314 4880 14324
rect 4036 14244 4682 14314
rect 4754 14244 4880 14314
rect 4036 14232 4880 14244
rect 4036 13404 4280 14232
rect 5340 13776 5584 14434
rect 6320 14433 6502 15180
rect 7050 15218 7552 15236
rect 7050 15156 7114 15218
rect 7182 15156 7552 15218
rect 7050 15140 7552 15156
rect 6321 14430 6502 14433
rect 6321 14334 6684 14430
rect 6321 14328 6502 14334
rect 6320 14294 6502 14328
rect 6320 14232 6350 14294
rect 6418 14232 6502 14294
rect 6320 14213 6502 14232
rect 6589 13938 6684 14334
rect 6584 13918 6948 13938
rect 6584 13856 6828 13918
rect 6896 13856 6948 13918
rect 6584 13846 6948 13856
rect 4822 13772 5584 13776
rect 4822 13770 6086 13772
rect 4822 13700 4884 13770
rect 4956 13754 6086 13770
rect 4956 13700 5862 13754
rect 4822 13692 5862 13700
rect 5930 13692 6086 13754
rect 4822 13688 6086 13692
rect 5340 13676 6086 13688
rect 4036 13384 4884 13404
rect 4036 13318 4576 13384
rect 4648 13318 4884 13384
rect 4036 13312 4884 13318
rect 4036 12658 4280 13312
rect 5340 12928 5584 13676
rect 6589 13470 6684 13846
rect 5948 13450 6684 13470
rect 5948 13390 5984 13450
rect 6052 13390 6684 13450
rect 7348 13752 7552 15140
rect 7838 14284 8072 16808
rect 7838 14222 7916 14284
rect 7984 14222 8072 14284
rect 7838 14188 8072 14222
rect 8902 16792 9242 16808
rect 11186 16792 11464 16808
rect 12704 16792 13034 16808
rect 8902 16632 9146 16792
rect 8902 16618 9710 16632
rect 8902 16562 9418 16618
rect 9474 16562 9710 16618
rect 8902 16540 9710 16562
rect 8902 15888 9146 16540
rect 9746 16080 10450 16086
rect 9746 16024 9842 16080
rect 9900 16024 10450 16080
rect 9746 15998 10450 16024
rect 10208 15916 10450 15998
rect 8902 15878 9804 15888
rect 8902 15818 9612 15878
rect 9674 15818 9804 15878
rect 8902 15796 9804 15818
rect 8902 15070 9146 15796
rect 10206 15348 10450 15916
rect 9700 15336 10450 15348
rect 9700 15274 9764 15336
rect 9832 15274 10450 15336
rect 11186 15784 11368 16792
rect 11186 15772 11762 15784
rect 11186 15710 11578 15772
rect 11646 15710 11762 15772
rect 11186 15688 11762 15710
rect 11186 15282 11368 15688
rect 9700 15260 10450 15274
rect 8902 15056 9766 15070
rect 8902 14990 9448 15056
rect 9514 14990 9766 15056
rect 8902 14978 9766 14990
rect 8902 14328 9146 14978
rect 10206 14742 10450 15260
rect 10954 15268 11368 15282
rect 10954 15206 10996 15268
rect 11064 15206 11368 15268
rect 10954 15184 11368 15206
rect 10206 14720 10892 14742
rect 10206 14658 10660 14720
rect 10728 14658 10892 14720
rect 10206 14646 10892 14658
rect 10206 14526 10450 14646
rect 9808 14512 10450 14526
rect 9808 14446 9878 14512
rect 9944 14446 10450 14512
rect 9808 14438 10450 14446
rect 8902 14318 9746 14328
rect 8902 14248 9548 14318
rect 9620 14248 9746 14318
rect 8902 14236 9746 14248
rect 7348 13738 7746 13752
rect 7348 13676 7656 13738
rect 7724 13676 7746 13738
rect 7348 13656 7746 13676
rect 7348 13394 7552 13656
rect 5948 13378 6684 13390
rect 5340 12916 6098 12928
rect 5340 12856 5996 12916
rect 6064 12856 6098 12916
rect 5340 12854 6098 12856
rect 4926 12844 6098 12854
rect 4926 12778 4990 12844
rect 5062 12832 6098 12844
rect 5062 12778 5584 12832
rect 4926 12766 5584 12778
rect 4036 12642 4952 12658
rect 4036 12576 4634 12642
rect 4708 12576 4952 12642
rect 4036 12566 4952 12576
rect 4036 11840 4280 12566
rect 5340 12110 5584 12766
rect 6589 12454 6684 13378
rect 7092 13378 7552 13394
rect 7092 13316 7136 13378
rect 7204 13316 7552 13378
rect 7092 13298 7552 13316
rect 6193 12432 6684 12454
rect 6193 12370 6280 12432
rect 6348 12370 6684 12432
rect 6193 12359 6684 12370
rect 4850 12100 5584 12110
rect 4850 12034 4906 12100
rect 4980 12034 5584 12100
rect 4850 12022 5584 12034
rect 5340 11906 5584 12022
rect 5340 11892 6100 11906
rect 4036 11820 4838 11840
rect 4036 11756 4560 11820
rect 4640 11756 4838 11820
rect 4036 11748 4838 11756
rect 5340 11830 6002 11892
rect 6070 11830 6100 11892
rect 5340 11810 6100 11830
rect 4036 11090 4280 11748
rect 5340 11294 5584 11810
rect 4936 11278 5584 11294
rect 4936 11214 4994 11278
rect 5074 11214 5584 11278
rect 4936 11200 5584 11214
rect 4036 11074 4904 11090
rect 4036 11010 4626 11074
rect 4706 11010 4904 11074
rect 4036 10998 4904 11010
rect 4036 10996 4280 10998
rect 5340 10554 5584 11200
rect 4852 10540 5584 10554
rect 4852 10476 4904 10540
rect 4984 10476 5584 10540
rect 4852 10448 5584 10476
rect 5340 9882 5584 10448
rect 7348 9882 7552 13298
rect 8902 13408 9146 14236
rect 10206 13780 10450 14438
rect 11186 14437 11368 15184
rect 11916 15222 12418 15240
rect 11916 15160 11980 15222
rect 12048 15160 12418 15222
rect 11916 15144 12418 15160
rect 11187 14434 11368 14437
rect 11187 14338 11550 14434
rect 11187 14332 11368 14338
rect 11186 14298 11368 14332
rect 11186 14236 11216 14298
rect 11284 14236 11368 14298
rect 11186 14217 11368 14236
rect 11455 13942 11550 14338
rect 11450 13922 11814 13942
rect 11450 13860 11694 13922
rect 11762 13860 11814 13922
rect 11450 13850 11814 13860
rect 9688 13776 10450 13780
rect 9688 13774 10952 13776
rect 9688 13704 9750 13774
rect 9822 13758 10952 13774
rect 9822 13704 10728 13758
rect 9688 13696 10728 13704
rect 10796 13696 10952 13758
rect 9688 13692 10952 13696
rect 10206 13680 10952 13692
rect 8902 13388 9750 13408
rect 8902 13322 9442 13388
rect 9514 13322 9750 13388
rect 8902 13316 9750 13322
rect 8902 12662 9146 13316
rect 10206 12932 10450 13680
rect 11455 13474 11550 13850
rect 10814 13454 11550 13474
rect 10814 13394 10850 13454
rect 10918 13394 11550 13454
rect 12214 13756 12418 15144
rect 12704 14288 12938 16792
rect 15198 15406 15426 16810
rect 16340 16722 16568 16810
rect 16340 16660 16430 16722
rect 16498 16660 16568 16722
rect 16340 16652 16568 16660
rect 17108 16714 17336 16810
rect 17108 16652 17188 16714
rect 17256 16652 17336 16714
rect 17108 16642 17336 16652
rect 17998 16716 18226 16810
rect 18452 16800 20542 16810
rect 17998 16654 18078 16716
rect 18146 16654 18226 16716
rect 17998 16638 18226 16654
rect 18596 16712 18824 16800
rect 18596 16650 18686 16712
rect 18754 16650 18824 16712
rect 18596 16642 18824 16650
rect 19364 16704 19592 16800
rect 19364 16642 19444 16704
rect 19512 16642 19592 16704
rect 19364 16632 19592 16642
rect 20254 16706 20482 16800
rect 20990 16794 23276 16810
rect 20254 16644 20334 16706
rect 20402 16644 20482 16706
rect 20254 16628 20482 16644
rect 21360 16706 21588 16794
rect 21360 16644 21450 16706
rect 21518 16644 21588 16706
rect 21360 16636 21588 16644
rect 22128 16698 22356 16794
rect 22128 16636 22208 16698
rect 22276 16636 22356 16698
rect 22128 16626 22356 16636
rect 23018 16700 23246 16794
rect 23018 16638 23098 16700
rect 23166 16638 23246 16700
rect 23018 16622 23246 16638
rect 16333 16184 16547 16199
rect 16333 16122 16410 16184
rect 16478 16122 16547 16184
rect 16333 16027 16547 16122
rect 17127 16174 17341 16185
rect 17127 16112 17196 16174
rect 17264 16112 17341 16174
rect 17127 16027 17341 16112
rect 17993 16174 18207 16191
rect 17993 16112 18076 16174
rect 18144 16112 18207 16174
rect 17993 16027 18207 16112
rect 18589 16174 18803 16189
rect 18589 16112 18666 16174
rect 18734 16112 18803 16174
rect 16197 16018 18300 16027
rect 16197 16017 18510 16018
rect 18589 16017 18803 16112
rect 19383 16164 19597 16175
rect 19383 16102 19452 16164
rect 19520 16102 19597 16164
rect 19383 16017 19597 16102
rect 20249 16164 20463 16181
rect 20249 16102 20332 16164
rect 20400 16102 20463 16164
rect 20249 16017 20463 16102
rect 21353 16168 21567 16183
rect 21353 16106 21430 16168
rect 21498 16106 21567 16168
rect 21353 16017 21567 16106
rect 16197 16011 21567 16017
rect 22147 16158 22361 16169
rect 22147 16096 22216 16158
rect 22284 16096 22361 16158
rect 22147 16011 22361 16096
rect 23013 16158 23227 16175
rect 23013 16096 23096 16158
rect 23164 16096 23227 16158
rect 23013 16027 23227 16096
rect 23657 16027 23871 17722
rect 22627 16011 23871 16027
rect 16197 16010 21710 16011
rect 21790 16010 21966 16011
rect 16197 16006 21966 16010
rect 22094 16006 23871 16011
rect 16197 15896 23871 16006
rect 16197 15813 23874 15896
rect 18292 15803 23874 15813
rect 20597 15797 23874 15803
rect 23270 15794 23874 15797
rect 15198 15178 24536 15406
rect 24310 15150 24536 15178
rect 24310 14870 24538 15150
rect 24310 14810 24400 14870
rect 24462 14810 24538 14870
rect 24310 14790 24538 14810
rect 26956 14766 27174 14788
rect 26956 14646 27000 14766
rect 27122 14646 27174 14766
rect 26956 14604 27174 14646
rect 27512 14492 27730 14510
rect 27512 14372 27550 14492
rect 27682 14372 27730 14492
rect 27512 14336 27730 14372
rect 12704 14226 12782 14288
rect 12850 14226 12938 14288
rect 12704 14192 12938 14226
rect 23852 14318 24212 14334
rect 23852 14258 23992 14318
rect 24054 14258 24212 14318
rect 23852 14128 24212 14258
rect 23852 13946 24204 14128
rect 12214 13742 12612 13756
rect 12214 13680 12522 13742
rect 12590 13680 12612 13742
rect 12214 13660 12612 13680
rect 15110 13726 24204 13946
rect 12214 13398 12418 13660
rect 10814 13382 11550 13394
rect 10206 12920 10964 12932
rect 10206 12860 10862 12920
rect 10930 12860 10964 12920
rect 10206 12858 10964 12860
rect 9792 12848 10964 12858
rect 9792 12782 9856 12848
rect 9928 12836 10964 12848
rect 9928 12782 10450 12836
rect 9792 12770 10450 12782
rect 8902 12646 9818 12662
rect 8902 12580 9500 12646
rect 9574 12580 9818 12646
rect 8902 12570 9818 12580
rect 8902 11844 9146 12570
rect 10206 12114 10450 12770
rect 11455 12458 11550 13382
rect 11958 13382 12418 13398
rect 11958 13320 12002 13382
rect 12070 13320 12418 13382
rect 11958 13302 12418 13320
rect 11059 12436 11550 12458
rect 11059 12374 11146 12436
rect 11214 12374 11550 12436
rect 11059 12363 11550 12374
rect 9716 12104 10450 12114
rect 9716 12038 9772 12104
rect 9846 12038 10450 12104
rect 9716 12026 10450 12038
rect 10206 11910 10450 12026
rect 10206 11896 10966 11910
rect 8902 11824 9704 11844
rect 8902 11760 9426 11824
rect 9506 11760 9704 11824
rect 8902 11752 9704 11760
rect 10206 11834 10868 11896
rect 10936 11834 10966 11896
rect 10206 11814 10966 11834
rect 8902 11094 9146 11752
rect 10206 11298 10450 11814
rect 9802 11282 10450 11298
rect 9802 11218 9860 11282
rect 9940 11218 10450 11282
rect 9802 11204 10450 11218
rect 8902 11078 9770 11094
rect 8902 11014 9492 11078
rect 9572 11014 9770 11078
rect 8902 11002 9770 11014
rect 8902 11000 9146 11002
rect 10206 10558 10450 11204
rect 9718 10544 10450 10558
rect 9718 10480 9770 10544
rect 9850 10480 10450 10544
rect 9718 10452 10450 10480
rect 10206 9944 10450 10452
rect 12214 9944 12418 13302
rect 15110 13586 24208 13726
rect 10206 9922 10540 9944
rect 12214 9922 12508 9944
rect 13258 9922 13626 9926
rect 8392 9890 14696 9922
rect 15110 9890 15470 13586
rect 8392 9886 15470 9890
rect 8312 9882 15470 9886
rect 800 9724 15470 9882
rect 800 9562 994 9724
rect 1146 9562 15470 9724
rect 800 9530 15470 9562
rect 800 9376 13253 9530
rect 6108 6638 6646 6736
rect 6108 6580 6226 6638
rect 6282 6580 6646 6638
rect 6108 6556 6646 6580
rect 372 6088 6274 6108
rect 372 6074 6170 6088
rect 372 5986 392 6074
rect 498 6030 6170 6074
rect 6226 6030 6274 6088
rect 498 5986 6274 6030
rect 372 5954 6274 5986
rect 6466 5814 6646 6556
rect 9652 6050 18838 6222
rect 9652 6042 11818 6050
rect 9652 5814 9832 6042
rect 802 5774 9844 5814
rect 802 5670 936 5774
rect 1052 5670 9844 5774
rect 802 5634 9844 5670
rect 2512 5578 2692 5634
rect 4378 5620 4558 5634
rect 2512 5520 2564 5578
rect 2620 5520 2692 5578
rect 2512 5506 2692 5520
rect 4628 5574 4808 5634
rect 6104 5620 6284 5634
rect 6572 5602 6766 5634
rect 8010 5620 8190 5634
rect 6572 5574 6762 5602
rect 4628 5570 4810 5574
rect 4628 5512 4686 5570
rect 4742 5512 4810 5570
rect 4628 5492 4810 5512
rect 6570 5570 6762 5574
rect 6570 5512 6638 5570
rect 6694 5512 6762 5570
rect 6570 5492 6762 5512
rect 8584 5576 8762 5634
rect 8584 5518 8640 5576
rect 8696 5574 8762 5576
rect 8696 5518 8764 5574
rect 8584 5498 8764 5518
rect 4628 5478 4808 5492
rect 6570 5488 6750 5492
rect 10128 5120 10308 6042
rect 10708 6000 10888 6042
rect 10708 5936 10774 6000
rect 10832 5936 10888 6000
rect 10708 5924 10888 5936
rect 12736 5986 12922 6050
rect 12736 5928 12796 5986
rect 12852 5928 12922 5986
rect 12736 5922 12922 5928
rect 12740 5908 12920 5922
rect 10972 5452 12936 5480
rect 10972 5394 11214 5452
rect 11270 5440 12936 5452
rect 11270 5394 12800 5440
rect 10972 5382 12800 5394
rect 12856 5382 12936 5440
rect 10972 5300 12936 5382
rect 10128 5062 10188 5120
rect 10244 5062 10308 5120
rect 2520 5040 2700 5048
rect 2520 4982 2584 5040
rect 2640 4982 2700 5040
rect 2520 4850 2700 4982
rect 4628 5024 4808 5048
rect 4628 4966 4690 5024
rect 4746 4966 4808 5024
rect 4380 4850 4560 4858
rect 4628 4850 4808 4966
rect 6580 5024 6760 5048
rect 6580 4966 6642 5024
rect 6698 4966 6760 5024
rect 6580 4948 6760 4966
rect 6092 4850 6272 4858
rect 6574 4850 6760 4948
rect 8582 5030 8762 5054
rect 10128 5046 10308 5062
rect 8582 4972 8644 5030
rect 8700 4972 8762 5030
rect 8002 4852 8182 4858
rect 8582 4852 8762 4972
rect 7674 4850 9835 4852
rect 198 4814 9835 4850
rect 198 4710 330 4814
rect 446 4710 9835 4814
rect 198 4670 9835 4710
rect 9652 4496 9832 4670
rect 10732 4580 10912 4598
rect 10732 4522 10788 4580
rect 10844 4522 10912 4580
rect 9652 4376 9834 4496
rect 10732 4376 10912 4522
rect 11576 4376 11756 5300
rect 13626 5174 13798 6050
rect 14696 5994 14882 6050
rect 14696 5952 14754 5994
rect 14698 5936 14754 5952
rect 14810 5952 14882 5994
rect 16690 6000 16876 6050
rect 17510 6042 18838 6050
rect 16690 5958 16748 6000
rect 14810 5936 14878 5952
rect 14698 5916 14878 5936
rect 16692 5942 16748 5958
rect 16804 5958 16876 6000
rect 16804 5942 16872 5958
rect 16692 5922 16872 5942
rect 14688 5454 16890 5480
rect 14688 5448 16752 5454
rect 14688 5390 14758 5448
rect 14814 5396 16752 5448
rect 16808 5396 16890 5454
rect 14814 5390 16890 5396
rect 14688 5308 16890 5390
rect 12976 5124 15154 5174
rect 12976 5080 15156 5124
rect 12976 5022 13032 5080
rect 13088 5074 15156 5080
rect 13088 5022 15034 5074
rect 12976 5016 15034 5022
rect 15090 5072 15156 5074
rect 15090 5016 15158 5072
rect 12976 5002 15158 5016
rect 14978 4996 15158 5002
rect 12974 4534 13154 4558
rect 12974 4476 13036 4534
rect 13092 4476 13154 4534
rect 9652 4368 11818 4376
rect 12974 4368 13154 4476
rect 14976 4528 15156 4552
rect 14976 4470 15038 4528
rect 15094 4470 15156 4528
rect 14976 4368 15156 4470
rect 15878 4368 16050 5308
rect 17648 5168 17828 6042
rect 18658 5428 18838 6042
rect 18658 5364 18726 5428
rect 18784 5364 18838 5428
rect 18658 5354 18838 5364
rect 17002 5106 17828 5168
rect 17000 5056 17828 5106
rect 17000 4998 17056 5056
rect 17112 4998 17828 5056
rect 17000 4988 17828 4998
rect 17000 4978 17180 4988
rect 18662 4880 18842 4888
rect 18662 4816 18720 4880
rect 18778 4816 18842 4880
rect 9652 4352 16050 4368
rect 16998 4510 17178 4534
rect 16998 4452 17060 4510
rect 17116 4452 17178 4510
rect 16998 4368 17178 4452
rect 18662 4376 18842 4816
rect 17510 4368 18840 4376
rect 16998 4352 18840 4368
rect 9652 4328 18840 4352
rect 9656 4196 18840 4328
rect 6082 3382 6656 3408
rect 6082 3320 6194 3382
rect 6254 3320 6656 3382
rect 6082 3228 6656 3320
rect 294 2828 6298 2858
rect 294 2808 6176 2828
rect 294 2714 384 2808
rect 484 2766 6176 2808
rect 6236 2766 6298 2828
rect 484 2714 6298 2766
rect 294 2664 6298 2714
rect 6476 2554 6656 3228
rect 794 2518 16633 2554
rect 794 2410 936 2518
rect 1068 2410 16633 2518
rect 794 2380 16633 2410
rect 794 2374 3426 2380
rect 3626 2374 5476 2380
rect 5676 2376 16633 2380
rect 2540 2318 2720 2374
rect 2540 2260 2604 2318
rect 2660 2260 2720 2318
rect 2540 2244 2720 2260
rect 4536 2314 4716 2374
rect 4536 2256 4592 2314
rect 4648 2256 4716 2314
rect 4536 2236 4716 2256
rect 6476 2314 6668 2376
rect 6476 2256 6544 2314
rect 6600 2256 6668 2314
rect 6476 2236 6668 2256
rect 8490 2320 8670 2376
rect 8490 2262 8546 2320
rect 8602 2262 8670 2320
rect 8490 2242 8670 2262
rect 10430 2320 10622 2376
rect 10430 2262 10498 2320
rect 10554 2262 10622 2320
rect 10430 2242 10622 2262
rect 12434 2320 12614 2376
rect 12434 2262 12490 2320
rect 12546 2262 12614 2320
rect 12434 2242 12614 2262
rect 14374 2320 14566 2376
rect 14374 2262 14442 2320
rect 14498 2262 14566 2320
rect 14374 2242 14566 2262
rect 16438 2320 16630 2376
rect 16438 2262 16506 2320
rect 16562 2262 16630 2320
rect 16438 2242 16630 2262
rect 10430 2238 10610 2242
rect 14374 2238 14554 2242
rect 16438 2238 16618 2242
rect 6476 2232 6656 2236
rect 2542 1778 2722 1790
rect 2542 1720 2604 1778
rect 2660 1720 2722 1778
rect 2542 1590 2722 1720
rect 4534 1768 4714 1792
rect 4534 1710 4596 1768
rect 4652 1710 4714 1768
rect 4534 1590 4714 1710
rect 6486 1768 6666 1792
rect 6486 1710 6548 1768
rect 6604 1710 6666 1768
rect 6486 1692 6666 1710
rect 6480 1590 6666 1692
rect 8488 1774 8668 1798
rect 8488 1716 8550 1774
rect 8606 1716 8668 1774
rect 8488 1596 8668 1716
rect 10440 1774 10620 1798
rect 10440 1716 10502 1774
rect 10558 1716 10620 1774
rect 10440 1698 10620 1716
rect 10434 1596 10620 1698
rect 12432 1774 12612 1798
rect 12432 1716 12494 1774
rect 12550 1716 12612 1774
rect 12432 1596 12612 1716
rect 14384 1774 14564 1798
rect 14384 1716 14446 1774
rect 14502 1716 14564 1774
rect 16448 1774 16628 1798
rect 16448 1716 16510 1774
rect 16566 1716 16628 1774
rect 14384 1698 14564 1716
rect 14378 1596 14564 1698
rect 16442 1686 16628 1716
rect 16442 1656 16626 1686
rect 7580 1592 9430 1596
rect 9630 1592 11402 1596
rect 11524 1592 13374 1596
rect 13574 1592 15346 1596
rect 7456 1590 15346 1592
rect 210 1586 3426 1590
rect 3626 1586 5476 1590
rect 5676 1588 15630 1590
rect 16446 1588 16626 1656
rect 5676 1586 16626 1588
rect 210 1548 16626 1586
rect 210 1438 336 1548
rect 456 1438 16626 1548
rect 210 1410 16626 1438
rect 30230 820 30542 862
rect 30230 716 30332 820
rect 30436 716 30542 820
rect 30230 638 30542 716
<< via3 >>
rect 996 17780 1066 17848
rect 322 16942 474 17104
rect 27000 14646 27122 14766
rect 27550 14372 27682 14492
rect 994 9562 1146 9724
rect 392 5986 498 6074
rect 936 5670 1052 5774
rect 330 4710 446 4814
rect 384 2714 484 2808
rect 936 2410 1068 2518
rect 336 1438 456 1548
rect 30332 716 30436 820
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44952 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 200 17104 600 44152
rect 200 16942 322 17104
rect 474 16942 600 17104
rect 200 6074 600 16942
rect 200 5986 392 6074
rect 498 5986 600 6074
rect 200 4814 600 5986
rect 200 4710 330 4814
rect 446 4710 600 4814
rect 200 2808 600 4710
rect 200 2714 384 2808
rect 484 2714 600 2808
rect 200 1548 600 2714
rect 200 1438 336 1548
rect 456 1438 600 1548
rect 200 1000 600 1438
rect 800 17848 1200 44152
rect 800 17780 996 17848
rect 1066 17780 1200 17848
rect 800 9724 1200 17780
rect 27110 14788 27170 45152
rect 26956 14766 27174 14788
rect 26956 14646 27000 14766
rect 27122 14646 27174 14766
rect 26956 14604 27174 14646
rect 27662 14510 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 27512 14492 27730 14510
rect 27512 14372 27550 14492
rect 27682 14372 27730 14492
rect 27512 14336 27730 14372
rect 800 9562 994 9724
rect 1146 9562 1200 9724
rect 800 5774 1200 9562
rect 800 5670 936 5774
rect 1052 5670 1200 5774
rect 800 2518 1200 5670
rect 800 2410 936 2518
rect 1068 2410 1200 2518
rect 800 1000 1200 2410
rect 30230 820 30542 862
rect 30230 716 30332 820
rect 30436 716 30542 820
rect 30230 638 30542 716
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 0 30542 638
use CLA  CLA_0
timestamp 1754940301
transform 1 0 4568 0 1 15292
box -138 -4838 3744 1342
use CLA  CLA_1
timestamp 1754940301
transform 1 0 9434 0 1 15296
box -138 -4838 3744 1342
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1754938408
transform -1 0 3278 0 -1 2288
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_1
timestamp 1754938408
transform -1 0 5348 0 -1 2284
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_2
timestamp 1754938408
transform -1 0 7300 0 -1 2284
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_3
timestamp 1754938408
transform -1 0 9302 0 -1 2290
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_4
timestamp 1754938408
transform -1 0 11254 0 -1 2290
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_5
timestamp 1754938408
transform -1 0 13246 0 -1 2290
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_6
timestamp 1754938408
transform -1 0 15198 0 -1 2290
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_7
timestamp 1754938408
transform -1 0 17262 0 -1 2290
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_8
timestamp 1754938408
transform -1 0 5442 0 -1 5540
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_9
timestamp 1754938408
transform -1 0 7394 0 -1 5540
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_10
timestamp 1754938408
transform -1 0 3308 0 -1 5548
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_11
timestamp 1754938408
transform -1 0 9396 0 -1 5546
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_12
timestamp 1754938408
transform -1 0 13552 0 -1 5956
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_13
timestamp 1754938408
transform -1 0 11490 0 -1 5968
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_14
timestamp 1754938408
transform -1 0 15510 0 -1 5964
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_15
timestamp 1754938408
transform -1 0 17504 0 -1 5970
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_16
timestamp 1754938408
transform -1 0 13788 0 -1 5050
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_17
timestamp 1754938408
transform -1 0 11518 0 -1 5094
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_18
timestamp 1754938408
transform -1 0 15790 0 -1 5044
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_19
timestamp 1754938408
transform -1 0 17812 0 -1 5026
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1754938408
transform -1 0 6358 0 -1 3340
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1754938408
transform -1 0 6388 0 -1 6600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1754938408
transform -1 0 9706 0 -1 17794
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1754938408
transform 1 0 16336 0 1 16150
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_4
timestamp 1754938408
transform 1 0 17104 0 1 16140
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_5
timestamp 1754938408
transform 1 0 17978 0 1 16142
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_6
timestamp 1754938408
transform 1 0 18592 0 1 16140
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_7
timestamp 1754938408
transform 1 0 19360 0 1 16130
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_8
timestamp 1754938408
transform 1 0 20234 0 1 16132
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_9
timestamp 1754938408
transform 1 0 21356 0 1 16134
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_10
timestamp 1754938408
transform 1 0 22124 0 1 16124
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_11
timestamp 1754938408
transform 1 0 22998 0 1 16126
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sky130_fd_sc_hd__mux2_1_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1754938408
transform -1 0 19130 0 -1 5396
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1754938408
transform 1 0 23484 0 1 14288
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 1760 0 -1 2284
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1723858470
transform -1 0 3826 0 -1 2286
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1723858470
transform -1 0 5778 0 -1 2286
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1723858470
transform -1 0 7780 0 -1 2292
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1723858470
transform -1 0 9732 0 -1 2292
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1723858470
transform -1 0 11724 0 -1 2292
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1723858470
transform -1 0 13676 0 -1 2292
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1723858470
transform -1 0 19290 0 -1 5412
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1723858470
transform -1 0 6086 0 -1 3340
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1723858470
transform 1 0 25454 0 1 14290
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_10
timestamp 1723858470
transform 1 0 23312 0 1 16130
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_11
timestamp 1723858470
transform 1 0 22454 0 1 16118
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_12
timestamp 1723858470
transform 1 0 21670 0 1 16140
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_13
timestamp 1723858470
transform 1 0 20554 0 1 16138
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_14
timestamp 1723858470
transform 1 0 19674 0 1 16134
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_15
timestamp 1723858470
transform 1 0 18910 0 1 16146
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_16
timestamp 1723858470
transform 1 0 17846 0 1 16146
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_17
timestamp 1723858470
transform 1 0 17418 0 1 16146
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_18
timestamp 1723858470
transform 1 0 16196 0 1 16150
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_19
timestamp 1723858470
transform -1 0 6544 0 -1 6598
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_20
timestamp 1723858470
transform -1 0 9848 0 -1 17790
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_21
timestamp 1723858470
transform 1 0 4300 0 1 16040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_22
timestamp 1723858470
transform 1 0 4434 0 1 15294
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_23
timestamp 1723858470
transform 1 0 4340 0 1 14478
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_24
timestamp 1723858470
transform 1 0 4432 0 1 13728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_25
timestamp 1723858470
transform 1 0 4336 0 1 12802
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_26
timestamp 1723858470
transform 1 0 4420 0 1 12062
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_27
timestamp 1723858470
transform 1 0 4336 0 1 11242
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_28
timestamp 1723858470
transform 1 0 4434 0 1 10504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_29
timestamp 1723858470
transform 1 0 5786 0 1 11852
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_30
timestamp 1723858470
transform 1 0 5800 0 1 12880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_31
timestamp 1723858470
transform 1 0 5682 0 1 13718
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_32
timestamp 1723858470
transform 1 0 5614 0 1 14694
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_33
timestamp 1723858470
transform 1 0 6480 0 1 15184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_34
timestamp 1723858470
transform 1 0 7288 0 1 13348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_35
timestamp 1723858470
transform 1 0 8314 0 1 13710
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_36
timestamp 1723858470
transform 1 0 12154 0 1 13352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_37
timestamp 1723858470
transform 1 0 13180 0 1 13714
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_38
timestamp 1723858470
transform 1 0 11346 0 1 15188
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_39
timestamp 1723858470
transform 1 0 10480 0 1 14698
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_40
timestamp 1723858470
transform 1 0 9206 0 1 14482
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_41
timestamp 1723858470
transform 1 0 9300 0 1 15298
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_42
timestamp 1723858470
transform 1 0 9166 0 1 16044
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_43
timestamp 1723858470
transform 1 0 10548 0 1 13722
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_44
timestamp 1723858470
transform 1 0 9298 0 1 13732
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_45
timestamp 1723858470
transform 1 0 10666 0 1 12884
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_46
timestamp 1723858470
transform 1 0 10652 0 1 11856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_47
timestamp 1723858470
transform 1 0 9300 0 1 10508
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_48
timestamp 1723858470
transform 1 0 9202 0 1 11246
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_49
timestamp 1723858470
transform 1 0 9286 0 1 12066
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_50
timestamp 1723858470
transform 1 0 9202 0 1 12806
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_51
timestamp 1723858470
transform -1 0 1780 0 -1 5546
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_52
timestamp 1723858470
transform -1 0 15750 0 -1 2292
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_53
timestamp 1723858470
transform -1 0 9976 0 -1 5964
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_54
timestamp 1723858470
transform -1 0 11672 0 -1 5106
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_55
timestamp 1723858470
transform -1 0 3920 0 -1 5542
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_56
timestamp 1723858470
transform -1 0 5872 0 -1 5542
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_57
timestamp 1723858470
transform -1 0 7874 0 -1 5548
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_58
timestamp 1723858470
transform -1 0 12030 0 -1 5958
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_59
timestamp 1723858470
transform -1 0 13988 0 -1 5966
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_60
timestamp 1723858470
transform -1 0 15982 0 -1 5972
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_61
timestamp 1723858470
transform -1 0 12266 0 -1 5052
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_62
timestamp 1723858470
transform -1 0 14268 0 -1 5046
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_63
timestamp 1723858470
transform -1 0 16290 0 -1 5028
box -38 -48 130 592
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
