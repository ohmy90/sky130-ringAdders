VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_ohmy90_adders
  CLASS BLOCK ;
  FOREIGN tt_um_ohmy90_adders ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564000 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 92.790 209.550 94.395 217.740 ;
      LAYER pwell ;
        RECT 94.725 217.105 95.510 217.535 ;
        RECT 94.685 210.055 95.595 217.040 ;
        RECT 94.685 209.885 95.785 210.055 ;
        RECT 94.685 209.810 95.595 209.885 ;
      LAYER nwell ;
        RECT 92.710 200.990 94.315 207.810 ;
      LAYER pwell ;
        RECT 94.645 207.175 95.430 207.605 ;
        RECT 94.605 201.495 95.515 207.155 ;
        RECT 94.605 201.350 95.705 201.495 ;
        RECT 95.535 201.325 95.705 201.350 ;
      LAYER nwell ;
        RECT 92.750 193.850 94.355 198.830 ;
      LAYER pwell ;
        RECT 94.685 198.195 95.470 198.625 ;
        RECT 94.645 194.355 95.555 198.080 ;
        RECT 94.645 194.210 95.745 194.355 ;
        RECT 95.575 194.185 95.745 194.210 ;
      LAYER nwell ;
        RECT 92.820 188.460 94.425 192.520 ;
      LAYER pwell ;
        RECT 94.755 191.885 95.540 192.315 ;
        RECT 94.715 188.965 95.625 191.865 ;
        RECT 94.715 188.795 95.815 188.965 ;
        RECT 94.715 188.705 95.625 188.795 ;
      LAYER nwell ;
        RECT 92.880 183.630 94.485 186.750 ;
      LAYER pwell ;
        RECT 94.815 186.115 95.600 186.545 ;
        RECT 94.775 184.135 95.685 186.065 ;
        RECT 94.775 183.965 95.875 184.135 ;
        RECT 94.775 183.875 95.685 183.965 ;
      LAYER nwell ;
        RECT 92.920 180.110 94.525 182.330 ;
      LAYER pwell ;
        RECT 94.855 181.695 95.640 182.125 ;
        RECT 94.815 180.615 95.725 181.665 ;
        RECT 94.815 180.445 95.915 180.615 ;
        RECT 94.815 180.315 95.725 180.445 ;
      LAYER nwell ;
        RECT 92.140 166.740 93.745 176.320 ;
      LAYER pwell ;
        RECT 94.075 175.685 94.860 176.115 ;
        RECT 94.035 172.900 94.945 175.665 ;
        RECT 94.265 171.360 94.945 172.900 ;
        RECT 94.045 170.450 94.945 171.360 ;
        RECT 94.265 167.245 94.945 170.450 ;
        RECT 94.265 167.075 95.135 167.245 ;
        RECT 94.265 166.935 94.945 167.075 ;
      LAYER nwell ;
        RECT 92.180 155.210 93.785 164.790 ;
      LAYER pwell ;
        RECT 94.115 164.155 94.900 164.585 ;
        RECT 94.075 161.370 94.985 164.135 ;
        RECT 94.305 159.830 94.985 161.370 ;
        RECT 94.085 158.920 94.985 159.830 ;
        RECT 94.305 155.715 94.985 158.920 ;
        RECT 94.305 155.545 95.175 155.715 ;
        RECT 94.305 155.405 94.985 155.545 ;
      LAYER nwell ;
        RECT 92.220 144.140 93.825 153.720 ;
      LAYER pwell ;
        RECT 94.155 153.085 94.940 153.515 ;
        RECT 94.115 150.300 95.025 153.065 ;
        RECT 94.345 148.760 95.025 150.300 ;
        RECT 94.125 147.850 95.025 148.760 ;
        RECT 94.345 144.645 95.025 147.850 ;
        RECT 94.345 144.475 95.215 144.645 ;
        RECT 94.345 144.335 95.025 144.475 ;
      LAYER nwell ;
        RECT 92.130 133.140 93.735 142.720 ;
      LAYER pwell ;
        RECT 94.065 142.085 94.850 142.515 ;
        RECT 94.025 139.300 94.935 142.065 ;
        RECT 94.255 137.760 94.935 139.300 ;
        RECT 94.035 136.850 94.935 137.760 ;
        RECT 94.255 133.645 94.935 136.850 ;
        RECT 94.255 133.475 95.125 133.645 ;
        RECT 94.255 133.335 94.935 133.475 ;
      LAYER nwell ;
        RECT 92.170 122.070 93.775 131.650 ;
      LAYER pwell ;
        RECT 94.105 131.015 94.890 131.445 ;
        RECT 94.065 128.230 94.975 130.995 ;
        RECT 94.295 126.690 94.975 128.230 ;
        RECT 94.075 125.780 94.975 126.690 ;
        RECT 94.295 122.575 94.975 125.780 ;
        RECT 94.295 122.405 95.165 122.575 ;
        RECT 94.295 122.265 94.975 122.405 ;
      LAYER nwell ;
        RECT 37.540 115.525 47.120 117.130 ;
        RECT 48.610 115.565 58.190 117.170 ;
        RECT 59.610 115.475 69.190 117.080 ;
        RECT 70.680 115.515 80.260 117.120 ;
        RECT 82.210 115.555 91.790 117.160 ;
      LAYER pwell ;
        RECT 41.250 115.005 42.160 115.225 ;
        RECT 43.700 115.005 46.465 115.235 ;
        RECT 37.735 114.325 46.465 115.005 ;
        RECT 46.485 114.410 46.915 115.195 ;
        RECT 52.320 115.045 53.230 115.265 ;
        RECT 54.770 115.045 57.535 115.275 ;
        RECT 48.805 114.365 57.535 115.045 ;
        RECT 57.555 114.450 57.985 115.235 ;
        RECT 63.320 114.955 64.230 115.175 ;
        RECT 65.770 114.955 68.535 115.185 ;
        RECT 37.875 114.135 38.045 114.325 ;
        RECT 48.945 114.175 49.115 114.365 ;
        RECT 59.805 114.275 68.535 114.955 ;
        RECT 68.555 114.360 68.985 115.145 ;
        RECT 74.390 114.995 75.300 115.215 ;
        RECT 76.840 114.995 79.605 115.225 ;
        RECT 70.875 114.315 79.605 114.995 ;
        RECT 79.625 114.400 80.055 115.185 ;
        RECT 85.920 115.035 86.830 115.255 ;
        RECT 88.370 115.035 91.135 115.265 ;
        RECT 82.405 114.355 91.135 115.035 ;
        RECT 91.155 114.440 91.585 115.225 ;
        RECT 59.945 114.085 60.115 114.275 ;
        RECT 71.015 114.125 71.185 114.315 ;
        RECT 82.545 114.165 82.715 114.355 ;
        RECT 48.215 88.885 48.385 89.055 ;
        RECT 48.215 88.865 48.320 88.885 ;
        RECT 47.390 87.955 48.320 88.865 ;
        RECT 48.465 87.995 48.895 88.780 ;
        RECT 82.790 88.335 82.960 88.505 ;
        RECT 87.160 88.345 87.330 88.515 ;
        RECT 82.790 88.315 82.895 88.335 ;
        RECT 87.160 88.325 87.265 88.345 ;
        RECT 78.900 88.145 79.070 88.315 ;
        RECT 78.900 88.125 79.005 88.145 ;
      LAYER nwell ;
        RECT 46.960 86.060 49.100 87.665 ;
      LAYER pwell ;
        RECT 77.420 87.255 77.850 88.040 ;
        RECT 78.075 87.215 79.005 88.125 ;
        RECT 81.350 87.445 81.780 88.230 ;
        RECT 81.965 87.405 82.895 88.315 ;
        RECT 85.680 87.455 86.110 88.240 ;
        RECT 86.335 87.415 87.265 88.325 ;
        RECT 91.000 88.295 91.170 88.465 ;
        RECT 96.610 88.305 96.780 88.475 ;
        RECT 100.980 88.315 101.150 88.485 ;
        RECT 91.000 88.275 91.105 88.295 ;
        RECT 96.610 88.285 96.715 88.305 ;
        RECT 100.980 88.295 101.085 88.315 ;
        RECT 89.570 87.405 90.000 88.190 ;
        RECT 90.175 87.365 91.105 88.275 ;
        RECT 95.150 87.415 95.580 88.200 ;
        RECT 95.785 87.375 96.715 88.285 ;
        RECT 99.480 87.425 99.910 88.210 ;
        RECT 100.155 87.385 101.085 88.295 ;
        RECT 104.820 88.265 104.990 88.435 ;
        RECT 104.820 88.245 104.925 88.265 ;
        RECT 103.330 87.375 103.760 88.160 ;
        RECT 103.995 87.335 104.925 88.245 ;
        RECT 107.890 88.255 108.060 88.425 ;
        RECT 112.260 88.265 112.430 88.435 ;
        RECT 107.890 88.235 107.995 88.255 ;
        RECT 112.260 88.245 112.365 88.265 ;
        RECT 107.065 87.325 107.995 88.235 ;
        RECT 108.220 87.365 108.650 88.150 ;
        RECT 110.760 87.375 111.190 88.160 ;
        RECT 111.435 87.335 112.365 88.245 ;
        RECT 116.100 88.215 116.270 88.385 ;
        RECT 116.100 88.195 116.205 88.215 ;
        RECT 115.275 87.285 116.205 88.195 ;
        RECT 116.420 87.325 116.850 88.110 ;
      LAYER nwell ;
        RECT 77.215 85.320 79.405 86.925 ;
        RECT 81.145 85.510 83.295 87.115 ;
        RECT 85.475 85.520 87.665 87.125 ;
        RECT 89.365 85.470 91.505 87.075 ;
        RECT 94.945 85.480 97.115 87.085 ;
        RECT 99.275 85.490 101.485 87.095 ;
        RECT 103.125 85.440 105.325 87.045 ;
        RECT 106.635 85.430 108.855 87.035 ;
        RECT 110.555 85.440 112.765 87.045 ;
        RECT 114.845 85.390 117.055 86.995 ;
        RECT 21.690 81.515 25.750 83.120 ;
        RECT 46.020 81.535 50.080 83.140 ;
        RECT 81.040 82.055 83.250 83.660 ;
        RECT 85.330 82.005 87.540 83.610 ;
        RECT 89.240 82.015 91.460 83.620 ;
        RECT 92.770 82.005 94.970 83.610 ;
        RECT 96.610 81.955 98.820 83.560 ;
        RECT 100.980 81.965 103.150 83.570 ;
        RECT 106.590 81.975 108.730 83.580 ;
        RECT 110.430 81.925 112.620 83.530 ;
        RECT 114.800 81.935 116.950 83.540 ;
      LAYER pwell ;
        RECT 21.895 80.400 22.325 81.185 ;
        RECT 22.385 80.315 25.555 81.225 ;
        RECT 46.225 80.420 46.655 81.205 ;
        RECT 46.715 80.335 49.885 81.245 ;
        RECT 81.245 80.940 81.675 81.725 ;
        RECT 81.890 80.855 82.820 81.765 ;
        RECT 81.890 80.835 81.995 80.855 ;
        RECT 81.825 80.665 81.995 80.835 ;
        RECT 85.730 80.805 86.660 81.715 ;
        RECT 86.905 80.890 87.335 81.675 ;
        RECT 89.445 80.900 89.875 81.685 ;
        RECT 90.100 80.815 91.030 81.725 ;
        RECT 85.730 80.785 85.835 80.805 ;
        RECT 90.100 80.795 90.205 80.815 ;
        RECT 85.665 80.615 85.835 80.785 ;
        RECT 90.035 80.625 90.205 80.795 ;
        RECT 93.170 80.805 94.100 81.715 ;
        RECT 94.335 80.890 94.765 81.675 ;
        RECT 93.170 80.785 93.275 80.805 ;
        RECT 93.105 80.615 93.275 80.785 ;
        RECT 97.010 80.755 97.940 81.665 ;
        RECT 98.185 80.840 98.615 81.625 ;
        RECT 101.380 80.765 102.310 81.675 ;
        RECT 102.515 80.850 102.945 81.635 ;
        RECT 106.990 80.775 107.920 81.685 ;
        RECT 108.095 80.860 108.525 81.645 ;
        RECT 97.010 80.735 97.115 80.755 ;
        RECT 101.380 80.745 101.485 80.765 ;
        RECT 106.990 80.755 107.095 80.775 ;
        RECT 96.945 80.565 97.115 80.735 ;
        RECT 101.315 80.575 101.485 80.745 ;
        RECT 106.925 80.585 107.095 80.755 ;
        RECT 110.830 80.725 111.760 81.635 ;
        RECT 111.985 80.810 112.415 81.595 ;
        RECT 115.200 80.735 116.130 81.645 ;
        RECT 116.315 80.820 116.745 81.605 ;
        RECT 110.830 80.705 110.935 80.725 ;
        RECT 115.200 80.715 115.305 80.735 ;
        RECT 110.765 80.535 110.935 80.705 ;
        RECT 115.135 80.545 115.305 80.715 ;
        RECT 22.485 80.125 22.655 80.315 ;
        RECT 46.815 80.145 46.985 80.335 ;
      LAYER nwell ;
        RECT 22.190 77.795 25.320 79.400 ;
      LAYER pwell ;
        RECT 22.395 76.680 22.825 77.465 ;
        RECT 23.975 77.415 24.925 77.505 ;
        RECT 22.995 76.595 24.925 77.415 ;
      LAYER nwell ;
        RECT 32.850 77.245 36.910 78.850 ;
        RECT 46.520 77.815 49.650 79.420 ;
      LAYER pwell ;
        RECT 35.120 76.725 36.255 76.955 ;
        RECT 22.995 76.575 23.145 76.595 ;
        RECT 22.975 76.405 23.145 76.575 ;
      LAYER nwell ;
        RECT 21.740 73.695 25.800 75.300 ;
        RECT 28.560 74.745 31.700 76.350 ;
      LAYER pwell ;
        RECT 33.045 76.045 36.255 76.725 ;
        RECT 36.275 76.130 36.705 76.915 ;
        RECT 46.725 76.700 47.155 77.485 ;
        RECT 48.305 77.435 49.255 77.525 ;
        RECT 47.325 76.615 49.255 77.435 ;
      LAYER nwell ;
        RECT 57.180 77.265 61.240 78.870 ;
      LAYER pwell ;
        RECT 59.450 76.745 60.585 76.975 ;
        RECT 47.325 76.595 47.475 76.615 ;
        RECT 47.305 76.425 47.475 76.595 ;
        RECT 33.185 75.855 33.355 76.045 ;
        RECT 29.895 74.365 30.845 74.455 ;
        RECT 28.915 73.545 30.845 74.365 ;
        RECT 31.065 73.630 31.495 74.415 ;
      LAYER nwell ;
        RECT 46.070 73.715 50.130 75.320 ;
        RECT 52.890 74.765 56.030 76.370 ;
      LAYER pwell ;
        RECT 57.375 76.065 60.585 76.745 ;
        RECT 60.605 76.150 61.035 76.935 ;
        RECT 57.515 75.875 57.685 76.065 ;
        RECT 54.225 74.385 55.175 74.475 ;
        RECT 53.245 73.565 55.175 74.385 ;
        RECT 55.395 73.650 55.825 74.435 ;
        RECT 53.245 73.545 53.395 73.565 ;
        RECT 28.915 73.525 29.065 73.545 ;
        RECT 21.945 72.580 22.375 73.365 ;
        RECT 22.435 72.495 25.605 73.405 ;
        RECT 28.895 73.355 29.065 73.525 ;
        RECT 46.275 72.600 46.705 73.385 ;
        RECT 46.765 72.515 49.935 73.425 ;
        RECT 53.225 73.375 53.395 73.545 ;
      LAYER nwell ;
        RECT 117.230 72.745 127.730 74.350 ;
      LAYER pwell ;
        RECT 22.535 72.305 22.705 72.495 ;
        RECT 46.865 72.325 47.035 72.515 ;
        RECT 120.630 72.440 121.980 72.475 ;
        RECT 119.690 72.395 121.980 72.440 ;
        RECT 118.750 72.225 121.980 72.395 ;
        RECT 125.055 72.455 125.975 72.475 ;
        RECT 125.055 72.225 127.075 72.455 ;
        RECT 117.425 71.795 127.075 72.225 ;
        RECT 117.425 71.760 120.620 71.795 ;
        RECT 117.425 71.715 119.680 71.760 ;
      LAYER nwell ;
        RECT 22.240 69.975 25.370 71.580 ;
        RECT 28.470 69.915 32.530 71.520 ;
        RECT 38.420 69.835 42.020 71.440 ;
        RECT 46.560 69.995 49.700 71.600 ;
      LAYER pwell ;
        RECT 117.425 71.545 119.185 71.715 ;
        RECT 121.980 71.545 127.075 71.795 ;
        RECT 127.095 71.630 127.525 72.415 ;
      LAYER nwell ;
        RECT 52.800 69.935 56.860 71.540 ;
        RECT 62.750 69.855 66.350 71.460 ;
      LAYER pwell ;
        RECT 117.565 71.355 117.735 71.545 ;
        RECT 22.445 68.860 22.875 69.645 ;
        RECT 24.025 69.595 24.975 69.685 ;
        RECT 23.045 68.775 24.975 69.595 ;
        RECT 28.675 68.800 29.105 69.585 ;
        RECT 31.200 69.395 32.335 69.625 ;
        RECT 23.045 68.755 23.195 68.775 ;
        RECT 23.025 68.585 23.195 68.755 ;
        RECT 29.125 68.715 32.335 69.395 ;
        RECT 29.265 68.525 29.435 68.715 ;
      LAYER nwell ;
        RECT 33.780 68.045 36.900 69.650 ;
      LAYER pwell ;
        RECT 40.420 69.345 41.365 69.545 ;
        RECT 38.615 68.665 41.365 69.345 ;
        RECT 41.385 68.720 41.815 69.505 ;
        RECT 46.765 68.880 47.195 69.665 ;
        RECT 48.355 69.615 49.305 69.705 ;
        RECT 47.375 68.795 49.305 69.615 ;
        RECT 53.005 68.820 53.435 69.605 ;
        RECT 55.530 69.415 56.665 69.645 ;
        RECT 47.375 68.775 47.525 68.795 ;
        RECT 38.760 68.445 38.930 68.665 ;
        RECT 40.420 68.635 41.365 68.665 ;
        RECT 47.355 68.605 47.525 68.775 ;
        RECT 53.455 68.735 56.665 69.415 ;
        RECT 53.595 68.545 53.765 68.735 ;
      LAYER nwell ;
        RECT 58.110 68.065 61.240 69.670 ;
      LAYER pwell ;
        RECT 64.750 69.365 65.695 69.565 ;
        RECT 62.945 68.685 65.695 69.365 ;
        RECT 65.715 68.740 66.145 69.525 ;
        RECT 63.090 68.465 63.260 68.685 ;
        RECT 64.750 68.655 65.695 68.685 ;
        RECT 35.025 67.525 35.955 67.755 ;
      LAYER nwell ;
        RECT 21.700 65.355 25.760 66.960 ;
        RECT 29.090 65.705 32.230 67.310 ;
      LAYER pwell ;
        RECT 34.120 66.845 35.955 67.525 ;
        RECT 36.265 66.930 36.695 67.715 ;
        RECT 59.355 67.545 60.285 67.775 ;
        RECT 34.120 66.825 34.285 66.845 ;
        RECT 34.115 66.655 34.285 66.825 ;
        RECT 21.905 64.240 22.335 65.025 ;
        RECT 22.395 64.155 25.565 65.065 ;
        RECT 29.295 64.590 29.725 65.375 ;
        RECT 31.115 65.185 32.035 65.415 ;
      LAYER nwell ;
        RECT 46.030 65.375 50.090 66.980 ;
        RECT 53.420 65.725 56.560 67.330 ;
      LAYER pwell ;
        RECT 58.450 66.865 60.285 67.545 ;
        RECT 60.605 66.950 61.035 67.735 ;
        RECT 58.450 66.845 58.615 66.865 ;
        RECT 58.445 66.675 58.615 66.845 ;
        RECT 29.745 64.505 32.035 65.185 ;
        RECT 29.885 64.315 30.055 64.505 ;
        RECT 46.235 64.260 46.665 65.045 ;
        RECT 46.725 64.175 49.895 65.085 ;
        RECT 53.625 64.610 54.055 65.395 ;
        RECT 55.445 65.205 56.365 65.435 ;
        RECT 54.075 64.525 56.365 65.205 ;
        RECT 54.215 64.335 54.385 64.525 ;
        RECT 22.495 63.965 22.665 64.155 ;
        RECT 46.825 63.985 46.995 64.175 ;
      LAYER nwell ;
        RECT 22.200 61.635 25.330 63.240 ;
      LAYER pwell ;
        RECT 22.405 60.520 22.835 61.305 ;
        RECT 23.985 61.255 24.935 61.345 ;
        RECT 23.005 60.435 24.935 61.255 ;
      LAYER nwell ;
        RECT 29.070 60.605 32.210 62.210 ;
        RECT 46.520 61.655 49.660 63.260 ;
      LAYER pwell ;
        RECT 46.725 60.540 47.155 61.325 ;
        RECT 48.315 61.275 49.265 61.365 ;
        RECT 47.335 60.455 49.265 61.275 ;
      LAYER nwell ;
        RECT 53.400 60.625 56.540 62.230 ;
      LAYER pwell ;
        RECT 47.335 60.435 47.485 60.455 ;
        RECT 23.005 60.415 23.155 60.435 ;
        RECT 22.985 60.245 23.155 60.415 ;
        RECT 29.275 59.490 29.705 60.275 ;
        RECT 30.865 60.225 31.815 60.315 ;
        RECT 47.315 60.265 47.485 60.435 ;
        RECT 29.885 59.405 31.815 60.225 ;
        RECT 53.605 59.510 54.035 60.295 ;
        RECT 55.195 60.245 56.145 60.335 ;
        RECT 54.215 59.425 56.145 60.245 ;
        RECT 54.215 59.405 54.365 59.425 ;
        RECT 29.885 59.385 30.035 59.405 ;
        RECT 29.865 59.215 30.035 59.385 ;
        RECT 54.195 59.235 54.365 59.405 ;
      LAYER nwell ;
        RECT 21.750 57.535 25.810 59.140 ;
        RECT 46.080 57.555 50.140 59.160 ;
      LAYER pwell ;
        RECT 21.955 56.420 22.385 57.205 ;
        RECT 22.445 56.335 25.615 57.245 ;
        RECT 46.285 56.440 46.715 57.225 ;
        RECT 46.775 56.355 49.945 57.265 ;
        RECT 22.545 56.145 22.715 56.335 ;
        RECT 46.875 56.165 47.045 56.355 ;
      LAYER nwell ;
        RECT 22.240 53.815 25.380 55.420 ;
        RECT 46.570 53.835 49.710 55.440 ;
      LAYER pwell ;
        RECT 22.445 52.700 22.875 53.485 ;
        RECT 24.035 53.435 24.985 53.525 ;
        RECT 23.055 52.615 24.985 53.435 ;
        RECT 46.775 52.720 47.205 53.505 ;
        RECT 48.365 53.455 49.315 53.545 ;
        RECT 47.385 52.635 49.315 53.455 ;
        RECT 47.385 52.615 47.535 52.635 ;
        RECT 23.055 52.595 23.205 52.615 ;
        RECT 23.035 52.425 23.205 52.595 ;
        RECT 47.365 52.445 47.535 52.615 ;
        RECT 31.625 32.915 31.795 33.085 ;
        RECT 31.625 32.895 31.730 32.915 ;
        RECT 30.800 31.985 31.730 32.895 ;
        RECT 31.905 32.025 32.335 32.810 ;
      LAYER nwell ;
        RECT 30.370 30.090 32.540 31.695 ;
      LAYER pwell ;
        RECT 57.130 29.735 57.300 29.925 ;
        RECT 49.655 28.865 50.085 29.650 ;
        RECT 50.270 29.055 57.445 29.735 ;
        RECT 67.440 29.675 67.610 29.865 ;
        RECT 77.230 29.715 77.400 29.905 ;
        RECT 87.200 29.745 87.370 29.935 ;
        RECT 50.270 28.825 51.200 29.055 ;
        RECT 56.515 28.825 57.445 29.055 ;
        RECT 59.955 28.805 60.385 29.590 ;
        RECT 60.580 28.995 67.755 29.675 ;
        RECT 60.580 28.765 61.510 28.995 ;
        RECT 66.825 28.765 67.755 28.995 ;
        RECT 69.745 28.845 70.175 29.630 ;
        RECT 70.370 29.035 77.545 29.715 ;
        RECT 70.370 28.805 71.300 29.035 ;
        RECT 76.615 28.805 77.545 29.035 ;
        RECT 79.725 28.875 80.155 29.660 ;
        RECT 80.340 29.065 87.515 29.745 ;
        RECT 80.340 28.835 81.270 29.065 ;
        RECT 86.585 28.835 87.515 29.065 ;
        RECT 16.220 27.635 16.390 27.825 ;
        RECT 8.745 26.765 9.175 27.550 ;
        RECT 9.360 26.955 16.535 27.635 ;
        RECT 26.890 27.595 27.060 27.785 ;
        RECT 36.650 27.595 36.820 27.785 ;
        RECT 46.660 27.625 46.830 27.815 ;
        RECT 9.360 26.725 10.290 26.955 ;
        RECT 15.605 26.725 16.535 26.955 ;
        RECT 19.415 26.725 19.845 27.510 ;
        RECT 20.030 26.915 27.205 27.595 ;
        RECT 20.030 26.685 20.960 26.915 ;
        RECT 26.275 26.685 27.205 26.915 ;
        RECT 29.165 26.725 29.595 27.510 ;
        RECT 29.790 26.915 36.965 27.595 ;
        RECT 29.790 26.685 30.720 26.915 ;
        RECT 36.035 26.685 36.965 26.915 ;
        RECT 39.175 26.755 39.605 27.540 ;
        RECT 39.800 26.945 46.975 27.625 ;
        RECT 39.800 26.715 40.730 26.945 ;
        RECT 46.045 26.715 46.975 26.945 ;
      LAYER nwell ;
        RECT 49.450 26.930 57.640 28.535 ;
        RECT 59.750 26.870 67.950 28.475 ;
        RECT 69.540 26.910 77.740 28.515 ;
        RECT 79.520 26.940 87.710 28.545 ;
      LAYER pwell ;
        RECT 95.060 26.875 95.230 27.065 ;
      LAYER nwell ;
        RECT 8.540 24.830 16.730 26.435 ;
        RECT 19.210 24.790 27.400 26.395 ;
        RECT 28.960 24.790 37.160 26.395 ;
        RECT 38.970 24.820 47.170 26.425 ;
      LAYER pwell ;
        RECT 91.745 26.195 95.645 26.875 ;
        RECT 94.715 25.965 95.645 26.195 ;
        RECT 95.665 26.005 96.095 26.790 ;
        RECT 57.270 25.365 57.440 25.555 ;
        RECT 50.410 24.685 57.585 25.365 ;
        RECT 50.410 24.455 51.340 24.685 ;
        RECT 56.655 24.455 57.585 24.685 ;
        RECT 57.605 24.495 58.035 25.280 ;
        RECT 68.620 25.145 68.790 25.335 ;
        RECT 61.155 24.275 61.585 25.060 ;
        RECT 61.760 24.465 68.935 25.145 ;
        RECT 78.630 25.115 78.800 25.305 ;
        RECT 61.760 24.235 62.690 24.465 ;
        RECT 68.005 24.235 68.935 24.465 ;
        RECT 71.155 24.245 71.585 25.030 ;
        RECT 71.770 24.435 78.945 25.115 ;
        RECT 88.740 25.025 88.910 25.215 ;
        RECT 71.770 24.205 72.700 24.435 ;
        RECT 78.015 24.205 78.945 24.435 ;
      LAYER nwell ;
        RECT 50.040 22.560 58.240 24.165 ;
      LAYER pwell ;
        RECT 81.275 24.155 81.705 24.940 ;
        RECT 81.880 24.345 89.055 25.025 ;
        RECT 81.880 24.115 82.810 24.345 ;
        RECT 88.125 24.115 89.055 24.345 ;
      LAYER nwell ;
        RECT 91.320 24.070 96.300 25.675 ;
        RECT 60.950 22.340 69.130 23.945 ;
        RECT 70.950 22.310 79.140 23.915 ;
        RECT 81.070 22.220 89.250 23.825 ;
      LAYER pwell ;
        RECT 31.475 16.615 31.645 16.785 ;
        RECT 31.475 16.595 31.580 16.615 ;
        RECT 29.985 15.725 30.415 16.510 ;
        RECT 30.650 15.685 31.580 16.595 ;
      LAYER nwell ;
        RECT 29.780 13.790 31.980 15.395 ;
      LAYER pwell ;
        RECT 16.070 11.335 16.240 11.525 ;
        RECT 8.595 10.465 9.025 11.250 ;
        RECT 9.210 10.655 16.385 11.335 ;
        RECT 26.420 11.315 26.590 11.505 ;
        RECT 36.180 11.315 36.350 11.505 ;
        RECT 46.190 11.345 46.360 11.535 ;
        RECT 55.950 11.345 56.120 11.535 ;
        RECT 65.910 11.345 66.080 11.535 ;
        RECT 75.670 11.345 75.840 11.535 ;
        RECT 85.990 11.345 86.160 11.535 ;
        RECT 9.210 10.425 10.140 10.655 ;
        RECT 15.455 10.425 16.385 10.655 ;
        RECT 18.945 10.445 19.375 11.230 ;
        RECT 19.560 10.635 26.735 11.315 ;
        RECT 19.560 10.405 20.490 10.635 ;
        RECT 25.805 10.405 26.735 10.635 ;
        RECT 28.725 10.445 29.155 11.230 ;
        RECT 29.320 10.635 36.495 11.315 ;
        RECT 29.320 10.405 30.250 10.635 ;
        RECT 35.565 10.405 36.495 10.635 ;
        RECT 38.715 10.475 39.145 11.260 ;
        RECT 39.330 10.665 46.505 11.345 ;
        RECT 39.330 10.435 40.260 10.665 ;
        RECT 45.575 10.435 46.505 10.665 ;
        RECT 48.495 10.475 48.925 11.260 ;
        RECT 49.090 10.665 56.265 11.345 ;
        RECT 49.090 10.435 50.020 10.665 ;
        RECT 55.335 10.435 56.265 10.665 ;
        RECT 58.435 10.475 58.865 11.260 ;
        RECT 59.050 10.665 66.225 11.345 ;
        RECT 59.050 10.435 59.980 10.665 ;
        RECT 65.295 10.435 66.225 10.665 ;
        RECT 68.205 10.475 68.635 11.260 ;
        RECT 68.810 10.665 75.985 11.345 ;
        RECT 68.810 10.435 69.740 10.665 ;
        RECT 75.055 10.435 75.985 10.665 ;
        RECT 78.515 10.475 78.945 11.260 ;
        RECT 79.130 10.665 86.305 11.345 ;
        RECT 79.130 10.435 80.060 10.665 ;
        RECT 85.375 10.435 86.305 10.665 ;
      LAYER nwell ;
        RECT 8.390 8.530 16.580 10.135 ;
        RECT 18.740 8.510 26.930 10.115 ;
        RECT 28.520 8.510 36.690 10.115 ;
        RECT 38.510 8.540 46.700 10.145 ;
        RECT 48.290 8.540 56.460 10.145 ;
        RECT 58.230 8.540 66.420 10.145 ;
        RECT 68.000 8.540 76.180 10.145 ;
        RECT 78.310 8.540 86.500 10.145 ;
      LAYER li1 ;
        RECT 92.895 217.465 93.065 217.550 ;
        RECT 95.615 217.465 95.785 217.550 ;
        RECT 92.895 217.175 94.230 217.465 ;
        RECT 94.890 217.175 95.785 217.465 ;
        RECT 92.895 216.910 93.065 217.175 ;
        RECT 95.615 216.910 95.785 217.175 ;
        RECT 92.895 216.700 93.865 216.910 ;
        RECT 94.815 216.700 95.785 216.910 ;
        RECT 92.895 216.030 93.065 216.700 ;
        RECT 93.235 216.200 95.445 216.530 ;
        RECT 92.895 215.860 93.865 216.030 ;
        RECT 92.895 215.190 93.065 215.860 ;
        RECT 94.035 215.690 94.205 216.200 ;
        RECT 93.235 215.360 94.205 215.690 ;
        RECT 92.895 215.020 93.865 215.190 ;
        RECT 92.895 214.350 93.065 215.020 ;
        RECT 94.035 214.850 94.205 215.360 ;
        RECT 94.795 215.690 94.985 216.200 ;
        RECT 95.615 216.030 95.785 216.700 ;
        RECT 95.155 215.860 95.785 216.030 ;
        RECT 94.795 215.360 95.445 215.690 ;
        RECT 93.235 214.520 94.205 214.850 ;
        RECT 92.895 214.180 93.865 214.350 ;
        RECT 92.895 213.510 93.065 214.180 ;
        RECT 94.035 214.010 94.205 214.520 ;
        RECT 93.235 213.680 94.205 214.010 ;
        RECT 92.895 213.340 93.865 213.510 ;
        RECT 92.895 212.670 93.065 213.340 ;
        RECT 94.035 213.170 94.205 213.680 ;
        RECT 93.235 212.840 94.205 213.170 ;
        RECT 92.895 212.500 93.865 212.670 ;
        RECT 92.895 211.830 93.065 212.500 ;
        RECT 94.035 212.330 94.205 212.840 ;
        RECT 93.235 212.000 94.205 212.330 ;
        RECT 92.895 211.660 93.865 211.830 ;
        RECT 92.895 210.990 93.065 211.660 ;
        RECT 94.035 211.490 94.205 212.000 ;
        RECT 93.235 211.160 94.205 211.490 ;
        RECT 92.895 210.820 93.865 210.990 ;
        RECT 92.895 210.150 93.065 210.820 ;
        RECT 94.035 210.650 94.205 211.160 ;
        RECT 93.235 210.320 94.205 210.650 ;
        RECT 92.895 209.940 94.215 210.150 ;
        RECT 92.895 209.740 93.065 209.940 ;
        RECT 94.385 209.825 94.625 215.265 ;
        RECT 94.795 214.850 94.985 215.360 ;
        RECT 95.615 215.190 95.785 215.860 ;
        RECT 95.155 215.020 95.785 215.190 ;
        RECT 94.795 214.520 95.445 214.850 ;
        RECT 94.795 214.010 94.985 214.520 ;
        RECT 95.615 214.350 95.785 215.020 ;
        RECT 95.155 214.180 95.785 214.350 ;
        RECT 94.795 213.680 95.445 214.010 ;
        RECT 94.795 213.170 94.985 213.680 ;
        RECT 95.615 213.510 95.785 214.180 ;
        RECT 95.155 213.340 95.785 213.510 ;
        RECT 94.795 212.840 95.445 213.170 ;
        RECT 94.795 212.330 94.985 212.840 ;
        RECT 95.615 212.670 95.785 213.340 ;
        RECT 95.155 212.500 95.785 212.670 ;
        RECT 94.795 212.000 95.445 212.330 ;
        RECT 94.795 211.490 94.985 212.000 ;
        RECT 95.615 211.830 95.785 212.500 ;
        RECT 95.155 211.660 95.785 211.830 ;
        RECT 94.795 211.160 95.445 211.490 ;
        RECT 94.795 210.650 94.985 211.160 ;
        RECT 95.615 210.990 95.785 211.660 ;
        RECT 95.155 210.820 95.785 210.990 ;
        RECT 94.795 210.320 95.445 210.650 ;
        RECT 95.615 210.150 95.785 210.820 ;
        RECT 94.815 209.920 95.785 210.150 ;
        RECT 95.615 209.740 95.785 209.920 ;
        RECT 92.815 207.535 92.985 207.620 ;
        RECT 95.535 207.535 95.705 207.620 ;
        RECT 92.815 207.245 94.150 207.535 ;
        RECT 94.810 207.245 95.705 207.535 ;
        RECT 92.815 207.075 92.985 207.245 ;
        RECT 95.535 207.075 95.705 207.245 ;
        RECT 92.815 206.735 93.785 207.075 ;
        RECT 92.815 205.890 92.985 206.735 ;
        RECT 93.955 206.725 94.905 207.075 ;
        RECT 95.075 206.735 95.705 207.075 ;
        RECT 93.955 206.390 94.125 206.725 ;
        RECT 93.155 206.060 94.125 206.390 ;
        RECT 92.815 205.720 93.785 205.890 ;
        RECT 92.815 205.050 92.985 205.720 ;
        RECT 93.955 205.550 94.125 206.060 ;
        RECT 93.155 205.220 94.125 205.550 ;
        RECT 92.815 204.880 93.785 205.050 ;
        RECT 92.815 204.210 92.985 204.880 ;
        RECT 93.955 204.710 94.125 205.220 ;
        RECT 93.155 204.380 94.125 204.710 ;
        RECT 92.815 204.040 93.785 204.210 ;
        RECT 92.815 203.370 92.985 204.040 ;
        RECT 93.955 203.870 94.125 204.380 ;
        RECT 93.155 203.540 94.125 203.870 ;
        RECT 92.815 203.200 93.785 203.370 ;
        RECT 92.815 202.530 92.985 203.200 ;
        RECT 93.955 203.030 94.125 203.540 ;
        RECT 93.155 202.700 94.125 203.030 ;
        RECT 92.815 202.360 93.785 202.530 ;
        RECT 92.815 201.690 92.985 202.360 ;
        RECT 93.955 202.190 94.125 202.700 ;
        RECT 93.155 201.860 94.125 202.190 ;
        RECT 94.295 201.860 94.545 206.450 ;
        RECT 94.715 206.390 94.905 206.725 ;
        RECT 94.715 206.060 95.365 206.390 ;
        RECT 94.715 205.550 94.905 206.060 ;
        RECT 95.535 205.890 95.705 206.735 ;
        RECT 95.075 205.720 95.705 205.890 ;
        RECT 94.715 205.220 95.365 205.550 ;
        RECT 94.715 204.710 94.905 205.220 ;
        RECT 95.535 205.050 95.705 205.720 ;
        RECT 95.075 204.880 95.705 205.050 ;
        RECT 94.715 204.380 95.365 204.710 ;
        RECT 94.715 203.870 94.905 204.380 ;
        RECT 95.535 204.210 95.705 204.880 ;
        RECT 95.075 204.040 95.705 204.210 ;
        RECT 94.715 203.540 95.365 203.870 ;
        RECT 94.715 203.030 94.905 203.540 ;
        RECT 95.535 203.370 95.705 204.040 ;
        RECT 95.075 203.200 95.705 203.370 ;
        RECT 94.715 202.700 95.365 203.030 ;
        RECT 94.715 202.190 94.905 202.700 ;
        RECT 95.535 202.530 95.705 203.200 ;
        RECT 95.075 202.360 95.705 202.530 ;
        RECT 94.715 201.860 95.365 202.190 ;
        RECT 93.955 201.690 94.125 201.860 ;
        RECT 94.715 201.690 94.905 201.860 ;
        RECT 95.535 201.690 95.705 202.360 ;
        RECT 92.815 201.435 93.785 201.690 ;
        RECT 92.815 201.180 92.985 201.435 ;
        RECT 93.955 201.265 94.905 201.690 ;
        RECT 95.075 201.435 95.705 201.690 ;
        RECT 95.535 201.180 95.705 201.435 ;
        RECT 92.855 198.555 93.025 198.640 ;
        RECT 95.575 198.555 95.745 198.640 ;
        RECT 92.855 198.265 94.190 198.555 ;
        RECT 94.850 198.265 95.745 198.555 ;
        RECT 92.855 198.040 93.025 198.265 ;
        RECT 92.855 197.740 93.825 198.040 ;
        RECT 93.995 197.775 94.945 198.095 ;
        RECT 95.575 198.045 95.745 198.265 ;
        RECT 92.855 197.070 93.025 197.740 ;
        RECT 93.995 197.570 94.165 197.775 ;
        RECT 93.195 197.240 94.165 197.570 ;
        RECT 92.855 196.900 93.825 197.070 ;
        RECT 92.855 196.230 93.025 196.900 ;
        RECT 93.995 196.730 94.165 197.240 ;
        RECT 93.195 196.400 94.165 196.730 ;
        RECT 92.855 196.060 93.825 196.230 ;
        RECT 92.855 195.390 93.025 196.060 ;
        RECT 93.995 195.890 94.165 196.400 ;
        RECT 93.195 195.560 94.165 195.890 ;
        RECT 92.855 195.220 93.825 195.390 ;
        RECT 92.855 194.550 93.025 195.220 ;
        RECT 93.995 195.050 94.165 195.560 ;
        RECT 93.195 194.720 94.165 195.050 ;
        RECT 94.335 194.720 94.585 197.575 ;
        RECT 94.755 197.570 94.945 197.775 ;
        RECT 95.115 197.740 95.745 198.045 ;
        RECT 94.755 197.240 95.405 197.570 ;
        RECT 94.755 196.730 94.945 197.240 ;
        RECT 95.575 197.070 95.745 197.740 ;
        RECT 95.115 196.900 95.745 197.070 ;
        RECT 94.755 196.400 95.405 196.730 ;
        RECT 94.755 195.890 94.945 196.400 ;
        RECT 95.575 196.230 95.745 196.900 ;
        RECT 95.115 196.060 95.745 196.230 ;
        RECT 94.755 195.560 95.405 195.890 ;
        RECT 94.755 195.050 94.945 195.560 ;
        RECT 95.575 195.390 95.745 196.060 ;
        RECT 95.115 195.220 95.745 195.390 ;
        RECT 94.755 194.720 95.405 195.050 ;
        RECT 92.855 194.295 93.825 194.550 ;
        RECT 93.995 194.470 94.165 194.720 ;
        RECT 94.755 194.470 94.945 194.720 ;
        RECT 95.575 194.550 95.745 195.220 ;
        RECT 92.855 194.040 93.025 194.295 ;
        RECT 93.995 194.125 94.945 194.470 ;
        RECT 95.115 194.295 95.745 194.550 ;
        RECT 95.575 194.040 95.745 194.295 ;
        RECT 92.925 192.245 93.095 192.330 ;
        RECT 95.645 192.245 95.815 192.330 ;
        RECT 92.925 191.955 94.260 192.245 ;
        RECT 94.920 191.955 95.815 192.245 ;
        RECT 92.925 191.685 93.095 191.955 ;
        RECT 92.925 191.515 93.555 191.685 ;
        RECT 92.925 190.845 93.095 191.515 ;
        RECT 94.045 191.435 95.005 191.785 ;
        RECT 95.645 191.685 95.815 191.955 ;
        RECT 95.180 191.435 95.815 191.685 ;
        RECT 94.045 191.345 94.235 191.435 ;
        RECT 93.265 191.015 94.235 191.345 ;
        RECT 94.825 191.265 95.005 191.435 ;
        RECT 92.925 190.675 93.895 190.845 ;
        RECT 92.925 190.005 93.095 190.675 ;
        RECT 94.065 190.505 94.235 191.015 ;
        RECT 93.265 190.175 94.235 190.505 ;
        RECT 92.925 189.835 93.895 190.005 ;
        RECT 92.925 189.075 93.095 189.835 ;
        RECT 94.065 189.665 94.235 190.175 ;
        RECT 93.265 189.335 94.235 189.665 ;
        RECT 92.925 188.780 94.235 189.075 ;
        RECT 92.925 188.650 93.095 188.780 ;
        RECT 94.405 188.755 94.655 191.265 ;
        RECT 94.825 191.095 95.475 191.265 ;
        RECT 94.825 190.425 95.005 191.095 ;
        RECT 95.645 190.845 95.815 191.435 ;
        RECT 95.185 190.675 95.815 190.845 ;
        RECT 94.825 190.255 95.475 190.425 ;
        RECT 94.825 189.585 95.005 190.255 ;
        RECT 95.645 190.005 95.815 190.675 ;
        RECT 95.185 189.835 95.815 190.005 ;
        RECT 94.825 189.415 95.475 189.585 ;
        RECT 95.645 189.045 95.815 189.835 ;
        RECT 95.185 188.780 95.815 189.045 ;
        RECT 95.645 188.650 95.815 188.780 ;
        RECT 92.985 186.475 93.155 186.560 ;
        RECT 95.705 186.475 95.875 186.560 ;
        RECT 92.985 186.185 94.320 186.475 ;
        RECT 94.980 186.185 95.875 186.475 ;
        RECT 92.985 185.935 93.155 186.185 ;
        RECT 92.985 185.725 93.615 185.935 ;
        RECT 94.105 185.725 95.065 185.990 ;
        RECT 95.705 185.975 95.875 186.185 ;
        RECT 95.240 185.725 95.875 185.975 ;
        RECT 92.985 185.055 93.155 185.725 ;
        RECT 94.105 185.555 94.295 185.725 ;
        RECT 94.885 185.555 95.065 185.725 ;
        RECT 93.325 185.225 94.295 185.555 ;
        RECT 92.985 184.885 93.955 185.055 ;
        RECT 92.985 184.215 93.155 184.885 ;
        RECT 94.125 184.715 94.295 185.225 ;
        RECT 93.325 184.385 94.295 184.715 ;
        RECT 92.985 183.950 94.295 184.215 ;
        RECT 92.985 183.820 93.155 183.950 ;
        RECT 94.465 183.925 94.715 185.555 ;
        RECT 94.885 185.225 95.535 185.555 ;
        RECT 94.885 184.715 95.065 185.225 ;
        RECT 95.705 185.055 95.875 185.725 ;
        RECT 95.245 184.885 95.875 185.055 ;
        RECT 94.885 184.385 95.535 184.715 ;
        RECT 95.705 184.215 95.875 184.885 ;
        RECT 95.245 183.950 95.875 184.215 ;
        RECT 95.705 183.820 95.875 183.950 ;
        RECT 93.025 182.055 93.195 182.140 ;
        RECT 95.745 182.055 95.915 182.140 ;
        RECT 93.025 181.765 94.360 182.055 ;
        RECT 95.020 181.765 95.915 182.055 ;
        RECT 93.025 181.535 93.195 181.765 ;
        RECT 95.745 181.535 95.915 181.765 ;
        RECT 93.025 181.325 94.335 181.535 ;
        RECT 94.925 181.325 95.915 181.535 ;
        RECT 93.025 180.655 93.195 181.325 ;
        RECT 93.365 180.905 95.575 181.155 ;
        RECT 93.365 180.825 94.345 180.905 ;
        RECT 94.945 180.825 95.575 180.905 ;
        RECT 93.025 180.425 94.335 180.655 ;
        RECT 93.025 180.300 93.195 180.425 ;
        RECT 94.505 180.405 94.755 180.735 ;
        RECT 95.745 180.655 95.915 181.325 ;
        RECT 94.925 180.425 95.915 180.655 ;
        RECT 95.745 180.300 95.915 180.425 ;
        RECT 92.245 176.045 92.415 176.130 ;
        RECT 94.965 176.045 95.135 176.130 ;
        RECT 92.245 175.755 93.580 176.045 ;
        RECT 94.240 175.755 95.135 176.045 ;
        RECT 92.245 175.075 92.415 175.755 ;
        RECT 92.585 175.345 94.795 175.580 ;
        RECT 92.585 175.245 93.570 175.345 ;
        RECT 94.140 175.325 94.795 175.345 ;
        RECT 92.245 174.860 93.555 175.075 ;
        RECT 92.245 173.650 92.415 174.860 ;
        RECT 93.725 174.670 94.055 175.175 ;
        RECT 94.965 175.155 95.135 175.755 ;
        RECT 94.505 174.835 95.135 175.155 ;
        RECT 92.605 174.600 94.055 174.670 ;
        RECT 92.605 174.400 94.705 174.600 ;
        RECT 92.605 174.340 93.335 174.400 ;
        RECT 94.435 174.350 94.705 174.400 ;
        RECT 93.475 174.160 94.310 174.230 ;
        RECT 93.475 174.150 94.745 174.160 ;
        RECT 92.630 174.040 94.745 174.150 ;
        RECT 92.630 173.995 93.605 174.040 ;
        RECT 92.630 173.820 93.555 173.995 ;
        RECT 94.185 173.985 94.745 174.040 ;
        RECT 92.245 173.480 93.425 173.650 ;
        RECT 92.245 172.735 92.415 173.480 ;
        RECT 93.725 173.320 94.055 173.870 ;
        RECT 94.225 173.830 94.745 173.985 ;
        RECT 94.965 173.660 95.135 174.835 ;
        RECT 94.355 173.490 95.135 173.660 ;
        RECT 93.725 173.310 94.750 173.320 ;
        RECT 92.585 173.120 94.750 173.310 ;
        RECT 92.585 172.970 93.520 173.120 ;
        RECT 94.225 172.990 94.750 173.120 ;
        RECT 92.245 172.420 92.915 172.735 ;
        RECT 92.245 170.710 92.415 172.420 ;
        RECT 93.145 172.410 93.520 172.970 ;
        RECT 93.725 172.240 94.055 172.950 ;
        RECT 94.965 172.725 95.135 173.490 ;
        RECT 94.435 172.515 95.135 172.725 ;
        RECT 92.715 172.070 94.685 172.240 ;
        RECT 92.715 171.355 92.885 172.070 ;
        RECT 93.055 171.580 94.345 171.900 ;
        RECT 94.015 171.435 94.345 171.580 ;
        RECT 94.515 171.455 94.685 172.070 ;
        RECT 93.085 171.220 93.805 171.410 ;
        RECT 92.585 171.050 92.915 171.130 ;
        RECT 94.515 171.050 94.685 171.285 ;
        RECT 92.585 170.880 94.685 171.050 ;
        RECT 92.245 170.540 93.215 170.710 ;
        RECT 93.475 170.540 93.805 170.710 ;
        RECT 92.245 168.635 92.415 170.540 ;
        RECT 93.475 170.370 93.735 170.540 ;
        RECT 93.985 170.420 94.285 170.880 ;
        RECT 94.965 170.700 95.135 172.515 ;
        RECT 92.690 170.200 93.735 170.370 ;
        RECT 93.955 170.220 94.285 170.420 ;
        RECT 94.465 170.330 95.135 170.700 ;
        RECT 92.690 169.265 92.860 170.200 ;
        RECT 93.030 169.670 93.395 170.030 ;
        RECT 93.565 170.010 93.735 170.200 ;
        RECT 93.565 169.840 94.685 170.010 ;
        RECT 93.030 169.500 94.315 169.670 ;
        RECT 93.330 169.090 93.925 169.330 ;
        RECT 94.095 169.145 94.315 169.500 ;
        RECT 94.515 169.335 94.685 169.840 ;
        RECT 92.585 168.920 93.140 169.055 ;
        RECT 94.515 168.975 94.685 169.140 ;
        RECT 94.245 168.920 94.685 168.975 ;
        RECT 92.585 168.805 94.685 168.920 ;
        RECT 93.010 168.750 94.375 168.805 ;
        RECT 94.965 168.635 95.135 170.330 ;
        RECT 92.245 168.370 92.875 168.635 ;
        RECT 92.245 167.775 92.415 168.370 ;
        RECT 93.385 168.300 94.335 168.580 ;
        RECT 94.505 168.385 95.135 168.635 ;
        RECT 92.585 167.945 94.705 168.130 ;
        RECT 94.965 167.775 95.135 168.385 ;
        RECT 92.245 167.445 92.915 167.775 ;
        RECT 93.085 167.540 94.415 167.770 ;
        RECT 92.245 166.930 92.415 167.445 ;
        RECT 93.085 167.275 93.255 167.540 ;
        RECT 92.585 167.105 93.255 167.275 ;
        RECT 93.425 167.020 94.075 167.370 ;
        RECT 94.245 167.275 94.415 167.540 ;
        RECT 94.585 167.445 95.135 167.775 ;
        RECT 94.245 167.105 94.705 167.275 ;
        RECT 94.965 166.930 95.135 167.445 ;
        RECT 92.285 164.515 92.455 164.600 ;
        RECT 95.005 164.515 95.175 164.600 ;
        RECT 92.285 164.225 93.620 164.515 ;
        RECT 94.280 164.225 95.175 164.515 ;
        RECT 92.285 163.545 92.455 164.225 ;
        RECT 92.625 163.815 94.835 164.050 ;
        RECT 92.625 163.715 93.610 163.815 ;
        RECT 94.180 163.795 94.835 163.815 ;
        RECT 92.285 163.330 93.595 163.545 ;
        RECT 92.285 162.120 92.455 163.330 ;
        RECT 93.765 163.140 94.095 163.645 ;
        RECT 95.005 163.625 95.175 164.225 ;
        RECT 94.545 163.305 95.175 163.625 ;
        RECT 92.645 163.070 94.095 163.140 ;
        RECT 92.645 162.870 94.745 163.070 ;
        RECT 92.645 162.810 93.375 162.870 ;
        RECT 94.475 162.820 94.745 162.870 ;
        RECT 93.515 162.630 94.350 162.700 ;
        RECT 93.515 162.620 94.785 162.630 ;
        RECT 92.670 162.510 94.785 162.620 ;
        RECT 92.670 162.465 93.645 162.510 ;
        RECT 92.670 162.290 93.595 162.465 ;
        RECT 94.225 162.455 94.785 162.510 ;
        RECT 92.285 161.950 93.465 162.120 ;
        RECT 92.285 161.205 92.455 161.950 ;
        RECT 93.765 161.790 94.095 162.340 ;
        RECT 94.265 162.300 94.785 162.455 ;
        RECT 95.005 162.130 95.175 163.305 ;
        RECT 94.395 161.960 95.175 162.130 ;
        RECT 93.765 161.780 94.790 161.790 ;
        RECT 92.625 161.590 94.790 161.780 ;
        RECT 92.625 161.440 93.560 161.590 ;
        RECT 94.265 161.460 94.790 161.590 ;
        RECT 92.285 160.890 92.955 161.205 ;
        RECT 92.285 159.180 92.455 160.890 ;
        RECT 93.185 160.880 93.560 161.440 ;
        RECT 93.765 160.710 94.095 161.420 ;
        RECT 95.005 161.195 95.175 161.960 ;
        RECT 94.475 160.985 95.175 161.195 ;
        RECT 92.755 160.540 94.725 160.710 ;
        RECT 92.755 159.825 92.925 160.540 ;
        RECT 93.095 160.050 94.385 160.370 ;
        RECT 94.055 159.905 94.385 160.050 ;
        RECT 94.555 159.925 94.725 160.540 ;
        RECT 93.125 159.690 93.845 159.880 ;
        RECT 92.625 159.520 92.955 159.600 ;
        RECT 94.555 159.520 94.725 159.755 ;
        RECT 92.625 159.350 94.725 159.520 ;
        RECT 92.285 159.010 93.255 159.180 ;
        RECT 93.515 159.010 93.845 159.180 ;
        RECT 92.285 157.105 92.455 159.010 ;
        RECT 93.515 158.840 93.775 159.010 ;
        RECT 94.025 158.890 94.325 159.350 ;
        RECT 95.005 159.170 95.175 160.985 ;
        RECT 92.730 158.670 93.775 158.840 ;
        RECT 93.995 158.690 94.325 158.890 ;
        RECT 94.505 158.800 95.175 159.170 ;
        RECT 92.730 157.735 92.900 158.670 ;
        RECT 93.070 158.140 93.435 158.500 ;
        RECT 93.605 158.480 93.775 158.670 ;
        RECT 93.605 158.310 94.725 158.480 ;
        RECT 93.070 157.970 94.355 158.140 ;
        RECT 93.370 157.560 93.965 157.800 ;
        RECT 94.135 157.615 94.355 157.970 ;
        RECT 94.555 157.805 94.725 158.310 ;
        RECT 92.625 157.390 93.180 157.525 ;
        RECT 94.555 157.445 94.725 157.610 ;
        RECT 94.285 157.390 94.725 157.445 ;
        RECT 92.625 157.275 94.725 157.390 ;
        RECT 93.050 157.220 94.415 157.275 ;
        RECT 95.005 157.105 95.175 158.800 ;
        RECT 92.285 156.840 92.915 157.105 ;
        RECT 92.285 156.245 92.455 156.840 ;
        RECT 93.425 156.770 94.375 157.050 ;
        RECT 94.545 156.855 95.175 157.105 ;
        RECT 92.625 156.415 94.745 156.600 ;
        RECT 95.005 156.245 95.175 156.855 ;
        RECT 92.285 155.915 92.955 156.245 ;
        RECT 93.125 156.010 94.455 156.240 ;
        RECT 92.285 155.400 92.455 155.915 ;
        RECT 93.125 155.745 93.295 156.010 ;
        RECT 92.625 155.575 93.295 155.745 ;
        RECT 93.465 155.490 94.115 155.840 ;
        RECT 94.285 155.745 94.455 156.010 ;
        RECT 94.625 155.915 95.175 156.245 ;
        RECT 94.285 155.575 94.745 155.745 ;
        RECT 95.005 155.400 95.175 155.915 ;
        RECT 92.325 153.445 92.495 153.530 ;
        RECT 95.045 153.445 95.215 153.530 ;
        RECT 92.325 153.155 93.660 153.445 ;
        RECT 94.320 153.155 95.215 153.445 ;
        RECT 92.325 152.475 92.495 153.155 ;
        RECT 92.665 152.745 94.875 152.980 ;
        RECT 92.665 152.645 93.650 152.745 ;
        RECT 94.220 152.725 94.875 152.745 ;
        RECT 92.325 152.260 93.635 152.475 ;
        RECT 92.325 151.050 92.495 152.260 ;
        RECT 93.805 152.070 94.135 152.575 ;
        RECT 95.045 152.555 95.215 153.155 ;
        RECT 94.585 152.235 95.215 152.555 ;
        RECT 92.685 152.000 94.135 152.070 ;
        RECT 92.685 151.800 94.785 152.000 ;
        RECT 92.685 151.740 93.415 151.800 ;
        RECT 94.515 151.750 94.785 151.800 ;
        RECT 93.555 151.560 94.390 151.630 ;
        RECT 93.555 151.550 94.825 151.560 ;
        RECT 92.710 151.440 94.825 151.550 ;
        RECT 92.710 151.395 93.685 151.440 ;
        RECT 92.710 151.220 93.635 151.395 ;
        RECT 94.265 151.385 94.825 151.440 ;
        RECT 92.325 150.880 93.505 151.050 ;
        RECT 92.325 150.135 92.495 150.880 ;
        RECT 93.805 150.720 94.135 151.270 ;
        RECT 94.305 151.230 94.825 151.385 ;
        RECT 95.045 151.060 95.215 152.235 ;
        RECT 94.435 150.890 95.215 151.060 ;
        RECT 93.805 150.710 94.830 150.720 ;
        RECT 92.665 150.520 94.830 150.710 ;
        RECT 92.665 150.370 93.600 150.520 ;
        RECT 94.305 150.390 94.830 150.520 ;
        RECT 92.325 149.820 92.995 150.135 ;
        RECT 92.325 148.110 92.495 149.820 ;
        RECT 93.225 149.810 93.600 150.370 ;
        RECT 93.805 149.640 94.135 150.350 ;
        RECT 95.045 150.125 95.215 150.890 ;
        RECT 94.515 149.915 95.215 150.125 ;
        RECT 92.795 149.470 94.765 149.640 ;
        RECT 92.795 148.755 92.965 149.470 ;
        RECT 93.135 148.980 94.425 149.300 ;
        RECT 94.095 148.835 94.425 148.980 ;
        RECT 94.595 148.855 94.765 149.470 ;
        RECT 93.165 148.620 93.885 148.810 ;
        RECT 92.665 148.450 92.995 148.530 ;
        RECT 94.595 148.450 94.765 148.685 ;
        RECT 92.665 148.280 94.765 148.450 ;
        RECT 92.325 147.940 93.295 148.110 ;
        RECT 93.555 147.940 93.885 148.110 ;
        RECT 92.325 146.035 92.495 147.940 ;
        RECT 93.555 147.770 93.815 147.940 ;
        RECT 94.065 147.820 94.365 148.280 ;
        RECT 95.045 148.100 95.215 149.915 ;
        RECT 92.770 147.600 93.815 147.770 ;
        RECT 94.035 147.620 94.365 147.820 ;
        RECT 94.545 147.730 95.215 148.100 ;
        RECT 92.770 146.665 92.940 147.600 ;
        RECT 93.110 147.070 93.475 147.430 ;
        RECT 93.645 147.410 93.815 147.600 ;
        RECT 93.645 147.240 94.765 147.410 ;
        RECT 93.110 146.900 94.395 147.070 ;
        RECT 93.410 146.490 94.005 146.730 ;
        RECT 94.175 146.545 94.395 146.900 ;
        RECT 94.595 146.735 94.765 147.240 ;
        RECT 92.665 146.320 93.220 146.455 ;
        RECT 94.595 146.375 94.765 146.540 ;
        RECT 94.325 146.320 94.765 146.375 ;
        RECT 92.665 146.205 94.765 146.320 ;
        RECT 93.090 146.150 94.455 146.205 ;
        RECT 95.045 146.035 95.215 147.730 ;
        RECT 92.325 145.770 92.955 146.035 ;
        RECT 92.325 145.175 92.495 145.770 ;
        RECT 93.465 145.700 94.415 145.980 ;
        RECT 94.585 145.785 95.215 146.035 ;
        RECT 92.665 145.345 94.785 145.530 ;
        RECT 95.045 145.175 95.215 145.785 ;
        RECT 92.325 144.845 92.995 145.175 ;
        RECT 93.165 144.940 94.495 145.170 ;
        RECT 92.325 144.330 92.495 144.845 ;
        RECT 93.165 144.675 93.335 144.940 ;
        RECT 92.665 144.505 93.335 144.675 ;
        RECT 93.505 144.420 94.155 144.770 ;
        RECT 94.325 144.675 94.495 144.940 ;
        RECT 94.665 144.845 95.215 145.175 ;
        RECT 94.325 144.505 94.785 144.675 ;
        RECT 95.045 144.330 95.215 144.845 ;
        RECT 92.235 142.445 92.405 142.530 ;
        RECT 94.955 142.445 95.125 142.530 ;
        RECT 92.235 142.155 93.570 142.445 ;
        RECT 94.230 142.155 95.125 142.445 ;
        RECT 92.235 141.475 92.405 142.155 ;
        RECT 92.575 141.745 94.785 141.980 ;
        RECT 92.575 141.645 93.560 141.745 ;
        RECT 94.130 141.725 94.785 141.745 ;
        RECT 92.235 141.260 93.545 141.475 ;
        RECT 92.235 140.050 92.405 141.260 ;
        RECT 93.715 141.070 94.045 141.575 ;
        RECT 94.955 141.555 95.125 142.155 ;
        RECT 94.495 141.235 95.125 141.555 ;
        RECT 92.595 141.000 94.045 141.070 ;
        RECT 92.595 140.800 94.695 141.000 ;
        RECT 92.595 140.740 93.325 140.800 ;
        RECT 94.425 140.750 94.695 140.800 ;
        RECT 93.465 140.560 94.300 140.630 ;
        RECT 93.465 140.550 94.735 140.560 ;
        RECT 92.620 140.440 94.735 140.550 ;
        RECT 92.620 140.395 93.595 140.440 ;
        RECT 92.620 140.220 93.545 140.395 ;
        RECT 94.175 140.385 94.735 140.440 ;
        RECT 92.235 139.880 93.415 140.050 ;
        RECT 92.235 139.135 92.405 139.880 ;
        RECT 93.715 139.720 94.045 140.270 ;
        RECT 94.215 140.230 94.735 140.385 ;
        RECT 94.955 140.060 95.125 141.235 ;
        RECT 94.345 139.890 95.125 140.060 ;
        RECT 93.715 139.710 94.740 139.720 ;
        RECT 92.575 139.520 94.740 139.710 ;
        RECT 92.575 139.370 93.510 139.520 ;
        RECT 94.215 139.390 94.740 139.520 ;
        RECT 92.235 138.820 92.905 139.135 ;
        RECT 92.235 137.110 92.405 138.820 ;
        RECT 93.135 138.810 93.510 139.370 ;
        RECT 93.715 138.640 94.045 139.350 ;
        RECT 94.955 139.125 95.125 139.890 ;
        RECT 94.425 138.915 95.125 139.125 ;
        RECT 92.705 138.470 94.675 138.640 ;
        RECT 92.705 137.755 92.875 138.470 ;
        RECT 93.045 137.980 94.335 138.300 ;
        RECT 94.005 137.835 94.335 137.980 ;
        RECT 94.505 137.855 94.675 138.470 ;
        RECT 93.075 137.620 93.795 137.810 ;
        RECT 92.575 137.450 92.905 137.530 ;
        RECT 94.505 137.450 94.675 137.685 ;
        RECT 92.575 137.280 94.675 137.450 ;
        RECT 92.235 136.940 93.205 137.110 ;
        RECT 93.465 136.940 93.795 137.110 ;
        RECT 92.235 135.035 92.405 136.940 ;
        RECT 93.465 136.770 93.725 136.940 ;
        RECT 93.975 136.820 94.275 137.280 ;
        RECT 94.955 137.100 95.125 138.915 ;
        RECT 92.680 136.600 93.725 136.770 ;
        RECT 93.945 136.620 94.275 136.820 ;
        RECT 94.455 136.730 95.125 137.100 ;
        RECT 92.680 135.665 92.850 136.600 ;
        RECT 93.020 136.070 93.385 136.430 ;
        RECT 93.555 136.410 93.725 136.600 ;
        RECT 93.555 136.240 94.675 136.410 ;
        RECT 93.020 135.900 94.305 136.070 ;
        RECT 93.320 135.490 93.915 135.730 ;
        RECT 94.085 135.545 94.305 135.900 ;
        RECT 94.505 135.735 94.675 136.240 ;
        RECT 92.575 135.320 93.130 135.455 ;
        RECT 94.505 135.375 94.675 135.540 ;
        RECT 94.235 135.320 94.675 135.375 ;
        RECT 92.575 135.205 94.675 135.320 ;
        RECT 93.000 135.150 94.365 135.205 ;
        RECT 94.955 135.035 95.125 136.730 ;
        RECT 92.235 134.770 92.865 135.035 ;
        RECT 92.235 134.175 92.405 134.770 ;
        RECT 93.375 134.700 94.325 134.980 ;
        RECT 94.495 134.785 95.125 135.035 ;
        RECT 92.575 134.345 94.695 134.530 ;
        RECT 94.955 134.175 95.125 134.785 ;
        RECT 92.235 133.845 92.905 134.175 ;
        RECT 93.075 133.940 94.405 134.170 ;
        RECT 92.235 133.330 92.405 133.845 ;
        RECT 93.075 133.675 93.245 133.940 ;
        RECT 92.575 133.505 93.245 133.675 ;
        RECT 93.415 133.420 94.065 133.770 ;
        RECT 94.235 133.675 94.405 133.940 ;
        RECT 94.575 133.845 95.125 134.175 ;
        RECT 94.235 133.505 94.695 133.675 ;
        RECT 94.955 133.330 95.125 133.845 ;
        RECT 92.275 131.375 92.445 131.460 ;
        RECT 94.995 131.375 95.165 131.460 ;
        RECT 92.275 131.085 93.610 131.375 ;
        RECT 94.270 131.085 95.165 131.375 ;
        RECT 92.275 130.405 92.445 131.085 ;
        RECT 92.615 130.675 94.825 130.910 ;
        RECT 92.615 130.575 93.600 130.675 ;
        RECT 94.170 130.655 94.825 130.675 ;
        RECT 92.275 130.190 93.585 130.405 ;
        RECT 92.275 128.980 92.445 130.190 ;
        RECT 93.755 130.000 94.085 130.505 ;
        RECT 94.995 130.485 95.165 131.085 ;
        RECT 94.535 130.165 95.165 130.485 ;
        RECT 92.635 129.930 94.085 130.000 ;
        RECT 92.635 129.730 94.735 129.930 ;
        RECT 92.635 129.670 93.365 129.730 ;
        RECT 94.465 129.680 94.735 129.730 ;
        RECT 93.505 129.490 94.340 129.560 ;
        RECT 93.505 129.480 94.775 129.490 ;
        RECT 92.660 129.370 94.775 129.480 ;
        RECT 92.660 129.325 93.635 129.370 ;
        RECT 92.660 129.150 93.585 129.325 ;
        RECT 94.215 129.315 94.775 129.370 ;
        RECT 92.275 128.810 93.455 128.980 ;
        RECT 92.275 128.065 92.445 128.810 ;
        RECT 93.755 128.650 94.085 129.200 ;
        RECT 94.255 129.160 94.775 129.315 ;
        RECT 94.995 128.990 95.165 130.165 ;
        RECT 94.385 128.820 95.165 128.990 ;
        RECT 93.755 128.640 94.780 128.650 ;
        RECT 92.615 128.450 94.780 128.640 ;
        RECT 92.615 128.300 93.550 128.450 ;
        RECT 94.255 128.320 94.780 128.450 ;
        RECT 92.275 127.750 92.945 128.065 ;
        RECT 92.275 126.040 92.445 127.750 ;
        RECT 93.175 127.740 93.550 128.300 ;
        RECT 93.755 127.570 94.085 128.280 ;
        RECT 94.995 128.055 95.165 128.820 ;
        RECT 94.465 127.845 95.165 128.055 ;
        RECT 92.745 127.400 94.715 127.570 ;
        RECT 92.745 126.685 92.915 127.400 ;
        RECT 93.085 126.910 94.375 127.230 ;
        RECT 94.045 126.765 94.375 126.910 ;
        RECT 94.545 126.785 94.715 127.400 ;
        RECT 93.115 126.550 93.835 126.740 ;
        RECT 92.615 126.380 92.945 126.460 ;
        RECT 94.545 126.380 94.715 126.615 ;
        RECT 92.615 126.210 94.715 126.380 ;
        RECT 92.275 125.870 93.245 126.040 ;
        RECT 93.505 125.870 93.835 126.040 ;
        RECT 92.275 123.965 92.445 125.870 ;
        RECT 93.505 125.700 93.765 125.870 ;
        RECT 94.015 125.750 94.315 126.210 ;
        RECT 94.995 126.030 95.165 127.845 ;
        RECT 92.720 125.530 93.765 125.700 ;
        RECT 93.985 125.550 94.315 125.750 ;
        RECT 94.495 125.660 95.165 126.030 ;
        RECT 92.720 124.595 92.890 125.530 ;
        RECT 93.060 125.000 93.425 125.360 ;
        RECT 93.595 125.340 93.765 125.530 ;
        RECT 93.595 125.170 94.715 125.340 ;
        RECT 93.060 124.830 94.345 125.000 ;
        RECT 93.360 124.420 93.955 124.660 ;
        RECT 94.125 124.475 94.345 124.830 ;
        RECT 94.545 124.665 94.715 125.170 ;
        RECT 92.615 124.250 93.170 124.385 ;
        RECT 94.545 124.305 94.715 124.470 ;
        RECT 94.275 124.250 94.715 124.305 ;
        RECT 92.615 124.135 94.715 124.250 ;
        RECT 93.040 124.080 94.405 124.135 ;
        RECT 94.995 123.965 95.165 125.660 ;
        RECT 92.275 123.700 92.905 123.965 ;
        RECT 92.275 123.105 92.445 123.700 ;
        RECT 93.415 123.630 94.365 123.910 ;
        RECT 94.535 123.715 95.165 123.965 ;
        RECT 92.615 123.275 94.735 123.460 ;
        RECT 94.995 123.105 95.165 123.715 ;
        RECT 92.275 122.775 92.945 123.105 ;
        RECT 93.115 122.870 94.445 123.100 ;
        RECT 92.275 122.260 92.445 122.775 ;
        RECT 93.115 122.605 93.285 122.870 ;
        RECT 92.615 122.435 93.285 122.605 ;
        RECT 93.455 122.350 94.105 122.700 ;
        RECT 94.275 122.605 94.445 122.870 ;
        RECT 94.615 122.775 95.165 123.105 ;
        RECT 94.275 122.435 94.735 122.605 ;
        RECT 94.995 122.260 95.165 122.775 ;
        RECT 37.730 116.855 46.930 117.025 ;
        RECT 48.800 116.895 58.000 117.065 ;
        RECT 37.905 116.185 38.075 116.685 ;
        RECT 38.245 116.355 38.575 116.855 ;
        RECT 37.905 116.015 38.570 116.185 ;
        RECT 37.820 115.195 38.170 115.845 ;
        RECT 38.340 115.025 38.570 116.015 ;
        RECT 37.905 114.855 38.570 115.025 ;
        RECT 37.905 114.565 38.075 114.855 ;
        RECT 38.245 114.305 38.575 114.685 ;
        RECT 38.745 114.565 38.930 116.685 ;
        RECT 39.170 116.395 39.435 116.855 ;
        RECT 39.605 116.260 39.855 116.685 ;
        RECT 40.065 116.410 41.170 116.580 ;
        RECT 39.550 116.130 39.855 116.260 ;
        RECT 39.100 114.935 39.380 115.885 ;
        RECT 39.550 115.025 39.720 116.130 ;
        RECT 39.890 115.345 40.130 115.940 ;
        RECT 40.300 115.875 40.830 116.240 ;
        RECT 40.300 115.175 40.470 115.875 ;
        RECT 41.000 115.795 41.170 116.410 ;
        RECT 41.340 116.055 41.510 116.855 ;
        RECT 41.680 116.355 41.930 116.685 ;
        RECT 42.155 116.385 43.040 116.555 ;
        RECT 41.000 115.705 41.510 115.795 ;
        RECT 39.550 114.895 39.775 115.025 ;
        RECT 39.945 114.955 40.470 115.175 ;
        RECT 40.640 115.535 41.510 115.705 ;
        RECT 39.185 114.305 39.435 114.765 ;
        RECT 39.605 114.755 39.775 114.895 ;
        RECT 40.640 114.755 40.810 115.535 ;
        RECT 41.340 115.465 41.510 115.535 ;
        RECT 41.020 115.285 41.220 115.315 ;
        RECT 41.680 115.285 41.850 116.355 ;
        RECT 42.020 115.465 42.210 116.185 ;
        RECT 41.020 114.985 41.850 115.285 ;
        RECT 42.380 115.255 42.700 116.215 ;
        RECT 39.605 114.585 39.940 114.755 ;
        RECT 40.135 114.585 40.810 114.755 ;
        RECT 41.130 114.305 41.500 114.805 ;
        RECT 41.680 114.755 41.850 114.985 ;
        RECT 42.235 114.925 42.700 115.255 ;
        RECT 42.870 115.545 43.040 116.385 ;
        RECT 43.220 116.355 43.535 116.855 ;
        RECT 43.770 116.125 44.110 116.685 ;
        RECT 43.210 115.750 44.110 116.125 ;
        RECT 44.280 115.845 44.450 116.855 ;
        RECT 43.920 115.545 44.110 115.750 ;
        RECT 44.620 115.795 44.950 116.640 ;
        RECT 45.140 115.935 45.470 116.665 ;
        RECT 44.620 115.715 45.030 115.795 ;
        RECT 44.795 115.665 45.030 115.715 ;
        RECT 42.870 115.215 43.750 115.545 ;
        RECT 43.920 115.215 44.670 115.545 ;
        RECT 42.870 114.755 43.040 115.215 ;
        RECT 43.920 115.045 44.120 115.215 ;
        RECT 44.840 115.085 45.030 115.665 ;
        RECT 44.785 115.045 45.030 115.085 ;
        RECT 41.680 114.585 42.085 114.755 ;
        RECT 42.255 114.585 43.040 114.755 ;
        RECT 43.315 114.305 43.525 114.835 ;
        RECT 43.790 114.520 44.120 115.045 ;
        RECT 44.630 114.960 45.030 115.045 ;
        RECT 45.200 115.545 45.470 115.935 ;
        RECT 45.660 115.715 45.875 116.855 ;
        RECT 46.045 115.700 46.380 116.685 ;
        RECT 45.200 115.215 45.975 115.545 ;
        RECT 44.290 114.305 44.460 114.915 ;
        RECT 44.630 114.525 44.960 114.960 ;
        RECT 45.200 114.835 45.400 115.215 ;
        RECT 46.145 115.130 46.380 115.700 ;
        RECT 46.555 115.690 46.845 116.855 ;
        RECT 48.975 116.225 49.145 116.725 ;
        RECT 49.315 116.395 49.645 116.895 ;
        RECT 48.975 116.055 49.640 116.225 ;
        RECT 48.890 115.235 49.240 115.885 ;
        RECT 45.150 114.565 45.400 114.835 ;
        RECT 45.635 114.305 45.955 114.765 ;
        RECT 46.125 114.475 46.380 115.130 ;
        RECT 49.410 115.065 49.640 116.055 ;
        RECT 46.555 114.305 46.845 115.030 ;
        RECT 48.975 114.895 49.640 115.065 ;
        RECT 48.975 114.605 49.145 114.895 ;
        RECT 49.315 114.345 49.645 114.725 ;
        RECT 49.815 114.605 50.000 116.725 ;
        RECT 50.240 116.435 50.505 116.895 ;
        RECT 50.675 116.300 50.925 116.725 ;
        RECT 51.135 116.450 52.240 116.620 ;
        RECT 50.620 116.170 50.925 116.300 ;
        RECT 50.170 114.975 50.450 115.925 ;
        RECT 50.620 115.065 50.790 116.170 ;
        RECT 50.960 115.385 51.200 115.980 ;
        RECT 51.370 115.915 51.900 116.280 ;
        RECT 51.370 115.215 51.540 115.915 ;
        RECT 52.070 115.835 52.240 116.450 ;
        RECT 52.410 116.095 52.580 116.895 ;
        RECT 52.750 116.395 53.000 116.725 ;
        RECT 53.225 116.425 54.110 116.595 ;
        RECT 52.070 115.745 52.580 115.835 ;
        RECT 50.620 114.935 50.845 115.065 ;
        RECT 51.015 114.995 51.540 115.215 ;
        RECT 51.710 115.575 52.580 115.745 ;
        RECT 50.255 114.345 50.505 114.805 ;
        RECT 50.675 114.795 50.845 114.935 ;
        RECT 51.710 114.795 51.880 115.575 ;
        RECT 52.410 115.505 52.580 115.575 ;
        RECT 52.090 115.325 52.290 115.355 ;
        RECT 52.750 115.325 52.920 116.395 ;
        RECT 53.090 115.505 53.280 116.225 ;
        RECT 52.090 115.025 52.920 115.325 ;
        RECT 53.450 115.295 53.770 116.255 ;
        RECT 50.675 114.625 51.010 114.795 ;
        RECT 51.205 114.625 51.880 114.795 ;
        RECT 52.200 114.345 52.570 114.845 ;
        RECT 52.750 114.795 52.920 115.025 ;
        RECT 53.305 114.965 53.770 115.295 ;
        RECT 53.940 115.585 54.110 116.425 ;
        RECT 54.290 116.395 54.605 116.895 ;
        RECT 54.840 116.165 55.180 116.725 ;
        RECT 54.280 115.790 55.180 116.165 ;
        RECT 55.350 115.885 55.520 116.895 ;
        RECT 54.990 115.585 55.180 115.790 ;
        RECT 55.690 115.835 56.020 116.680 ;
        RECT 56.210 115.975 56.540 116.705 ;
        RECT 55.690 115.755 56.100 115.835 ;
        RECT 55.865 115.705 56.100 115.755 ;
        RECT 53.940 115.255 54.820 115.585 ;
        RECT 54.990 115.255 55.740 115.585 ;
        RECT 53.940 114.795 54.110 115.255 ;
        RECT 54.990 115.085 55.190 115.255 ;
        RECT 55.910 115.125 56.100 115.705 ;
        RECT 55.855 115.085 56.100 115.125 ;
        RECT 52.750 114.625 53.155 114.795 ;
        RECT 53.325 114.625 54.110 114.795 ;
        RECT 54.385 114.345 54.595 114.875 ;
        RECT 54.860 114.560 55.190 115.085 ;
        RECT 55.700 115.000 56.100 115.085 ;
        RECT 56.270 115.585 56.540 115.975 ;
        RECT 56.730 115.755 56.945 116.895 ;
        RECT 57.115 115.740 57.450 116.725 ;
        RECT 56.270 115.255 57.045 115.585 ;
        RECT 55.360 114.345 55.530 114.955 ;
        RECT 55.700 114.565 56.030 115.000 ;
        RECT 56.270 114.875 56.470 115.255 ;
        RECT 57.215 115.170 57.450 115.740 ;
        RECT 57.625 115.730 57.915 116.895 ;
        RECT 59.800 116.805 69.000 116.975 ;
        RECT 70.870 116.845 80.070 117.015 ;
        RECT 82.400 116.885 91.600 117.055 ;
        RECT 59.975 116.135 60.145 116.635 ;
        RECT 60.315 116.305 60.645 116.805 ;
        RECT 59.975 115.965 60.640 116.135 ;
        RECT 56.220 114.605 56.470 114.875 ;
        RECT 56.705 114.345 57.025 114.805 ;
        RECT 57.195 114.515 57.450 115.170 ;
        RECT 59.890 115.145 60.240 115.795 ;
        RECT 57.625 114.345 57.915 115.070 ;
        RECT 60.410 114.975 60.640 115.965 ;
        RECT 59.975 114.805 60.640 114.975 ;
        RECT 59.975 114.515 60.145 114.805 ;
        RECT 37.730 114.135 46.930 114.305 ;
        RECT 48.800 114.175 58.000 114.345 ;
        RECT 60.315 114.255 60.645 114.635 ;
        RECT 60.815 114.515 61.000 116.635 ;
        RECT 61.240 116.345 61.505 116.805 ;
        RECT 61.675 116.210 61.925 116.635 ;
        RECT 62.135 116.360 63.240 116.530 ;
        RECT 61.620 116.080 61.925 116.210 ;
        RECT 61.170 114.885 61.450 115.835 ;
        RECT 61.620 114.975 61.790 116.080 ;
        RECT 61.960 115.295 62.200 115.890 ;
        RECT 62.370 115.825 62.900 116.190 ;
        RECT 62.370 115.125 62.540 115.825 ;
        RECT 63.070 115.745 63.240 116.360 ;
        RECT 63.410 116.005 63.580 116.805 ;
        RECT 63.750 116.305 64.000 116.635 ;
        RECT 64.225 116.335 65.110 116.505 ;
        RECT 63.070 115.655 63.580 115.745 ;
        RECT 61.620 114.845 61.845 114.975 ;
        RECT 62.015 114.905 62.540 115.125 ;
        RECT 62.710 115.485 63.580 115.655 ;
        RECT 61.255 114.255 61.505 114.715 ;
        RECT 61.675 114.705 61.845 114.845 ;
        RECT 62.710 114.705 62.880 115.485 ;
        RECT 63.410 115.415 63.580 115.485 ;
        RECT 63.090 115.235 63.290 115.265 ;
        RECT 63.750 115.235 63.920 116.305 ;
        RECT 64.090 115.415 64.280 116.135 ;
        RECT 63.090 114.935 63.920 115.235 ;
        RECT 64.450 115.205 64.770 116.165 ;
        RECT 61.675 114.535 62.010 114.705 ;
        RECT 62.205 114.535 62.880 114.705 ;
        RECT 63.200 114.255 63.570 114.755 ;
        RECT 63.750 114.705 63.920 114.935 ;
        RECT 64.305 114.875 64.770 115.205 ;
        RECT 64.940 115.495 65.110 116.335 ;
        RECT 65.290 116.305 65.605 116.805 ;
        RECT 65.840 116.075 66.180 116.635 ;
        RECT 65.280 115.700 66.180 116.075 ;
        RECT 66.350 115.795 66.520 116.805 ;
        RECT 65.990 115.495 66.180 115.700 ;
        RECT 66.690 115.745 67.020 116.590 ;
        RECT 67.210 115.885 67.540 116.615 ;
        RECT 66.690 115.665 67.100 115.745 ;
        RECT 66.865 115.615 67.100 115.665 ;
        RECT 64.940 115.165 65.820 115.495 ;
        RECT 65.990 115.165 66.740 115.495 ;
        RECT 64.940 114.705 65.110 115.165 ;
        RECT 65.990 114.995 66.190 115.165 ;
        RECT 66.910 115.035 67.100 115.615 ;
        RECT 66.855 114.995 67.100 115.035 ;
        RECT 63.750 114.535 64.155 114.705 ;
        RECT 64.325 114.535 65.110 114.705 ;
        RECT 65.385 114.255 65.595 114.785 ;
        RECT 65.860 114.470 66.190 114.995 ;
        RECT 66.700 114.910 67.100 114.995 ;
        RECT 67.270 115.495 67.540 115.885 ;
        RECT 67.730 115.665 67.945 116.805 ;
        RECT 68.115 115.650 68.450 116.635 ;
        RECT 67.270 115.165 68.045 115.495 ;
        RECT 66.360 114.255 66.530 114.865 ;
        RECT 66.700 114.475 67.030 114.910 ;
        RECT 67.270 114.785 67.470 115.165 ;
        RECT 68.215 115.080 68.450 115.650 ;
        RECT 68.625 115.640 68.915 116.805 ;
        RECT 71.045 116.175 71.215 116.675 ;
        RECT 71.385 116.345 71.715 116.845 ;
        RECT 71.045 116.005 71.710 116.175 ;
        RECT 70.960 115.185 71.310 115.835 ;
        RECT 67.220 114.515 67.470 114.785 ;
        RECT 67.705 114.255 68.025 114.715 ;
        RECT 68.195 114.425 68.450 115.080 ;
        RECT 71.480 115.015 71.710 116.005 ;
        RECT 68.625 114.255 68.915 114.980 ;
        RECT 71.045 114.845 71.710 115.015 ;
        RECT 71.045 114.555 71.215 114.845 ;
        RECT 71.385 114.295 71.715 114.675 ;
        RECT 71.885 114.555 72.070 116.675 ;
        RECT 72.310 116.385 72.575 116.845 ;
        RECT 72.745 116.250 72.995 116.675 ;
        RECT 73.205 116.400 74.310 116.570 ;
        RECT 72.690 116.120 72.995 116.250 ;
        RECT 72.240 114.925 72.520 115.875 ;
        RECT 72.690 115.015 72.860 116.120 ;
        RECT 73.030 115.335 73.270 115.930 ;
        RECT 73.440 115.865 73.970 116.230 ;
        RECT 73.440 115.165 73.610 115.865 ;
        RECT 74.140 115.785 74.310 116.400 ;
        RECT 74.480 116.045 74.650 116.845 ;
        RECT 74.820 116.345 75.070 116.675 ;
        RECT 75.295 116.375 76.180 116.545 ;
        RECT 74.140 115.695 74.650 115.785 ;
        RECT 72.690 114.885 72.915 115.015 ;
        RECT 73.085 114.945 73.610 115.165 ;
        RECT 73.780 115.525 74.650 115.695 ;
        RECT 72.325 114.295 72.575 114.755 ;
        RECT 72.745 114.745 72.915 114.885 ;
        RECT 73.780 114.745 73.950 115.525 ;
        RECT 74.480 115.455 74.650 115.525 ;
        RECT 74.160 115.275 74.360 115.305 ;
        RECT 74.820 115.275 74.990 116.345 ;
        RECT 75.160 115.455 75.350 116.175 ;
        RECT 74.160 114.975 74.990 115.275 ;
        RECT 75.520 115.245 75.840 116.205 ;
        RECT 72.745 114.575 73.080 114.745 ;
        RECT 73.275 114.575 73.950 114.745 ;
        RECT 74.270 114.295 74.640 114.795 ;
        RECT 74.820 114.745 74.990 114.975 ;
        RECT 75.375 114.915 75.840 115.245 ;
        RECT 76.010 115.535 76.180 116.375 ;
        RECT 76.360 116.345 76.675 116.845 ;
        RECT 76.910 116.115 77.250 116.675 ;
        RECT 76.350 115.740 77.250 116.115 ;
        RECT 77.420 115.835 77.590 116.845 ;
        RECT 77.060 115.535 77.250 115.740 ;
        RECT 77.760 115.785 78.090 116.630 ;
        RECT 78.280 115.925 78.610 116.655 ;
        RECT 77.760 115.705 78.170 115.785 ;
        RECT 77.935 115.655 78.170 115.705 ;
        RECT 76.010 115.205 76.890 115.535 ;
        RECT 77.060 115.205 77.810 115.535 ;
        RECT 76.010 114.745 76.180 115.205 ;
        RECT 77.060 115.035 77.260 115.205 ;
        RECT 77.980 115.075 78.170 115.655 ;
        RECT 77.925 115.035 78.170 115.075 ;
        RECT 74.820 114.575 75.225 114.745 ;
        RECT 75.395 114.575 76.180 114.745 ;
        RECT 76.455 114.295 76.665 114.825 ;
        RECT 76.930 114.510 77.260 115.035 ;
        RECT 77.770 114.950 78.170 115.035 ;
        RECT 78.340 115.535 78.610 115.925 ;
        RECT 78.800 115.705 79.015 116.845 ;
        RECT 79.185 115.690 79.520 116.675 ;
        RECT 78.340 115.205 79.115 115.535 ;
        RECT 77.430 114.295 77.600 114.905 ;
        RECT 77.770 114.515 78.100 114.950 ;
        RECT 78.340 114.825 78.540 115.205 ;
        RECT 79.285 115.120 79.520 115.690 ;
        RECT 79.695 115.680 79.985 116.845 ;
        RECT 82.575 116.215 82.745 116.715 ;
        RECT 82.915 116.385 83.245 116.885 ;
        RECT 82.575 116.045 83.240 116.215 ;
        RECT 82.490 115.225 82.840 115.875 ;
        RECT 78.290 114.555 78.540 114.825 ;
        RECT 78.775 114.295 79.095 114.755 ;
        RECT 79.265 114.465 79.520 115.120 ;
        RECT 83.010 115.055 83.240 116.045 ;
        RECT 79.695 114.295 79.985 115.020 ;
        RECT 82.575 114.885 83.240 115.055 ;
        RECT 82.575 114.595 82.745 114.885 ;
        RECT 82.915 114.335 83.245 114.715 ;
        RECT 83.415 114.595 83.600 116.715 ;
        RECT 83.840 116.425 84.105 116.885 ;
        RECT 84.275 116.290 84.525 116.715 ;
        RECT 84.735 116.440 85.840 116.610 ;
        RECT 84.220 116.160 84.525 116.290 ;
        RECT 83.770 114.965 84.050 115.915 ;
        RECT 84.220 115.055 84.390 116.160 ;
        RECT 84.560 115.375 84.800 115.970 ;
        RECT 84.970 115.905 85.500 116.270 ;
        RECT 84.970 115.205 85.140 115.905 ;
        RECT 85.670 115.825 85.840 116.440 ;
        RECT 86.010 116.085 86.180 116.885 ;
        RECT 86.350 116.385 86.600 116.715 ;
        RECT 86.825 116.415 87.710 116.585 ;
        RECT 85.670 115.735 86.180 115.825 ;
        RECT 84.220 114.925 84.445 115.055 ;
        RECT 84.615 114.985 85.140 115.205 ;
        RECT 85.310 115.565 86.180 115.735 ;
        RECT 83.855 114.335 84.105 114.795 ;
        RECT 84.275 114.785 84.445 114.925 ;
        RECT 85.310 114.785 85.480 115.565 ;
        RECT 86.010 115.495 86.180 115.565 ;
        RECT 85.690 115.315 85.890 115.345 ;
        RECT 86.350 115.315 86.520 116.385 ;
        RECT 86.690 115.495 86.880 116.215 ;
        RECT 85.690 115.015 86.520 115.315 ;
        RECT 87.050 115.285 87.370 116.245 ;
        RECT 84.275 114.615 84.610 114.785 ;
        RECT 84.805 114.615 85.480 114.785 ;
        RECT 85.800 114.335 86.170 114.835 ;
        RECT 86.350 114.785 86.520 115.015 ;
        RECT 86.905 114.955 87.370 115.285 ;
        RECT 87.540 115.575 87.710 116.415 ;
        RECT 87.890 116.385 88.205 116.885 ;
        RECT 88.440 116.155 88.780 116.715 ;
        RECT 87.880 115.780 88.780 116.155 ;
        RECT 88.950 115.875 89.120 116.885 ;
        RECT 88.590 115.575 88.780 115.780 ;
        RECT 89.290 115.825 89.620 116.670 ;
        RECT 89.810 115.965 90.140 116.695 ;
        RECT 89.290 115.745 89.700 115.825 ;
        RECT 89.465 115.695 89.700 115.745 ;
        RECT 87.540 115.245 88.420 115.575 ;
        RECT 88.590 115.245 89.340 115.575 ;
        RECT 87.540 114.785 87.710 115.245 ;
        RECT 88.590 115.075 88.790 115.245 ;
        RECT 89.510 115.115 89.700 115.695 ;
        RECT 89.455 115.075 89.700 115.115 ;
        RECT 86.350 114.615 86.755 114.785 ;
        RECT 86.925 114.615 87.710 114.785 ;
        RECT 87.985 114.335 88.195 114.865 ;
        RECT 88.460 114.550 88.790 115.075 ;
        RECT 89.300 114.990 89.700 115.075 ;
        RECT 89.870 115.575 90.140 115.965 ;
        RECT 90.330 115.745 90.545 116.885 ;
        RECT 90.715 115.730 91.050 116.715 ;
        RECT 89.870 115.245 90.645 115.575 ;
        RECT 88.960 114.335 89.130 114.945 ;
        RECT 89.300 114.555 89.630 114.990 ;
        RECT 89.870 114.865 90.070 115.245 ;
        RECT 90.815 115.160 91.050 115.730 ;
        RECT 91.225 115.720 91.515 116.885 ;
        RECT 89.820 114.595 90.070 114.865 ;
        RECT 90.305 114.335 90.625 114.795 ;
        RECT 90.795 114.505 91.050 115.160 ;
        RECT 91.225 114.335 91.515 115.060 ;
        RECT 59.800 114.085 69.000 114.255 ;
        RECT 70.870 114.125 80.070 114.295 ;
        RECT 82.400 114.165 91.600 114.335 ;
        RECT 47.150 88.885 48.910 89.055 ;
        RECT 47.480 88.085 47.810 88.715 ;
        RECT 47.480 87.485 47.710 88.085 ;
        RECT 47.980 88.065 48.210 88.885 ;
        RECT 48.535 88.160 48.825 88.885 ;
        RECT 81.335 88.335 83.105 88.505 ;
        RECT 85.665 88.345 87.475 88.515 ;
        RECT 77.405 88.145 79.215 88.315 ;
        RECT 47.880 87.655 48.210 87.895 ;
        RECT 47.480 86.505 47.810 87.485 ;
        RECT 47.980 86.335 48.190 87.475 ;
        RECT 48.535 86.335 48.825 87.500 ;
        RECT 77.490 87.420 77.780 88.145 ;
        RECT 78.165 87.345 78.495 87.975 ;
        RECT 47.150 86.165 48.910 86.335 ;
        RECT 77.490 85.595 77.780 86.760 ;
        RECT 78.165 86.745 78.395 87.345 ;
        RECT 78.665 87.325 78.895 88.145 ;
        RECT 81.420 87.610 81.710 88.335 ;
        RECT 82.055 87.535 82.385 88.165 ;
        RECT 78.565 86.915 78.895 87.155 ;
        RECT 78.165 85.765 78.495 86.745 ;
        RECT 78.665 85.595 78.875 86.735 ;
        RECT 81.420 85.785 81.710 86.950 ;
        RECT 82.055 86.935 82.285 87.535 ;
        RECT 82.555 87.515 82.785 88.335 ;
        RECT 85.750 87.620 86.040 88.345 ;
        RECT 86.425 87.545 86.755 88.175 ;
        RECT 82.455 87.105 82.785 87.345 ;
        RECT 82.055 85.955 82.385 86.935 ;
        RECT 82.555 85.785 82.765 86.925 ;
        RECT 85.750 85.795 86.040 86.960 ;
        RECT 86.425 86.945 86.655 87.545 ;
        RECT 86.925 87.525 87.155 88.345 ;
        RECT 89.555 88.295 91.315 88.465 ;
        RECT 95.135 88.305 96.925 88.475 ;
        RECT 99.465 88.315 101.295 88.485 ;
        RECT 89.640 87.570 89.930 88.295 ;
        RECT 90.265 87.495 90.595 88.125 ;
        RECT 86.825 87.115 87.155 87.355 ;
        RECT 86.425 85.965 86.755 86.945 ;
        RECT 86.925 85.795 87.135 86.935 ;
        RECT 81.335 85.615 83.105 85.785 ;
        RECT 85.665 85.625 87.475 85.795 ;
        RECT 89.640 85.745 89.930 86.910 ;
        RECT 90.265 86.895 90.495 87.495 ;
        RECT 90.765 87.475 90.995 88.295 ;
        RECT 95.220 87.580 95.510 88.305 ;
        RECT 95.875 87.505 96.205 88.135 ;
        RECT 90.665 87.065 90.995 87.305 ;
        RECT 90.265 85.915 90.595 86.895 ;
        RECT 90.765 85.745 90.975 86.885 ;
        RECT 95.220 85.755 95.510 86.920 ;
        RECT 95.875 86.905 96.105 87.505 ;
        RECT 96.375 87.485 96.605 88.305 ;
        RECT 99.550 87.590 99.840 88.315 ;
        RECT 100.245 87.515 100.575 88.145 ;
        RECT 96.275 87.075 96.605 87.315 ;
        RECT 95.875 85.925 96.205 86.905 ;
        RECT 96.375 85.755 96.585 86.895 ;
        RECT 99.550 85.765 99.840 86.930 ;
        RECT 100.245 86.915 100.475 87.515 ;
        RECT 100.745 87.495 100.975 88.315 ;
        RECT 103.315 88.265 105.135 88.435 ;
        RECT 103.400 87.540 103.690 88.265 ;
        RECT 104.085 87.465 104.415 88.095 ;
        RECT 100.645 87.085 100.975 87.325 ;
        RECT 100.245 85.935 100.575 86.915 ;
        RECT 100.745 85.765 100.955 86.905 ;
        RECT 77.405 85.425 79.215 85.595 ;
        RECT 89.555 85.575 91.315 85.745 ;
        RECT 95.135 85.585 96.925 85.755 ;
        RECT 99.465 85.595 101.295 85.765 ;
        RECT 103.400 85.715 103.690 86.880 ;
        RECT 104.085 86.865 104.315 87.465 ;
        RECT 104.585 87.445 104.815 88.265 ;
        RECT 106.825 88.255 108.665 88.425 ;
        RECT 110.745 88.265 112.575 88.435 ;
        RECT 107.155 87.455 107.485 88.085 ;
        RECT 104.485 87.035 104.815 87.275 ;
        RECT 104.085 85.885 104.415 86.865 ;
        RECT 107.155 86.855 107.385 87.455 ;
        RECT 107.655 87.435 107.885 88.255 ;
        RECT 108.290 87.530 108.580 88.255 ;
        RECT 110.830 87.540 111.120 88.265 ;
        RECT 111.525 87.465 111.855 88.095 ;
        RECT 107.555 87.025 107.885 87.265 ;
        RECT 104.585 85.715 104.795 86.855 ;
        RECT 107.155 85.875 107.485 86.855 ;
        RECT 103.315 85.545 105.135 85.715 ;
        RECT 107.655 85.705 107.865 86.845 ;
        RECT 108.290 85.705 108.580 86.870 ;
        RECT 110.830 85.715 111.120 86.880 ;
        RECT 111.525 86.865 111.755 87.465 ;
        RECT 112.025 87.445 112.255 88.265 ;
        RECT 115.035 88.215 116.865 88.385 ;
        RECT 115.365 87.415 115.695 88.045 ;
        RECT 111.925 87.035 112.255 87.275 ;
        RECT 111.525 85.885 111.855 86.865 ;
        RECT 112.025 85.715 112.235 86.855 ;
        RECT 115.365 86.815 115.595 87.415 ;
        RECT 115.865 87.395 116.095 88.215 ;
        RECT 116.490 87.490 116.780 88.215 ;
        RECT 115.765 86.985 116.095 87.225 ;
        RECT 115.365 85.835 115.695 86.815 ;
        RECT 106.825 85.535 108.665 85.705 ;
        RECT 110.745 85.545 112.575 85.715 ;
        RECT 115.865 85.665 116.075 86.805 ;
        RECT 116.490 85.665 116.780 86.830 ;
        RECT 115.035 85.495 116.865 85.665 ;
        RECT 81.230 83.385 83.060 83.555 ;
        RECT 21.880 82.845 25.560 83.015 ;
        RECT 46.210 82.865 49.890 83.035 ;
        RECT 21.965 81.680 22.255 82.845 ;
        RECT 22.425 81.995 22.805 82.675 ;
        RECT 23.395 81.995 23.565 82.845 ;
        RECT 23.735 82.165 24.065 82.675 ;
        RECT 24.235 82.335 24.405 82.845 ;
        RECT 24.575 82.165 24.975 82.675 ;
        RECT 23.735 81.995 24.975 82.165 ;
        RECT 22.425 81.035 22.595 81.995 ;
        RECT 22.765 81.655 24.070 81.825 ;
        RECT 25.155 81.745 25.475 82.675 ;
        RECT 22.765 81.205 23.010 81.655 ;
        RECT 23.180 81.285 23.730 81.485 ;
        RECT 23.900 81.455 24.070 81.655 ;
        RECT 24.845 81.575 25.475 81.745 ;
        RECT 46.295 81.700 46.585 82.865 ;
        RECT 46.755 82.015 47.135 82.695 ;
        RECT 47.725 82.015 47.895 82.865 ;
        RECT 48.065 82.185 48.395 82.695 ;
        RECT 48.565 82.355 48.735 82.865 ;
        RECT 48.905 82.185 49.305 82.695 ;
        RECT 48.065 82.015 49.305 82.185 ;
        RECT 23.900 81.285 24.275 81.455 ;
        RECT 24.445 81.035 24.675 81.535 ;
        RECT 21.965 80.295 22.255 81.020 ;
        RECT 22.425 80.865 24.675 81.035 ;
        RECT 22.475 80.295 22.805 80.685 ;
        RECT 22.975 80.545 23.145 80.865 ;
        RECT 24.845 80.695 25.015 81.575 ;
        RECT 23.315 80.295 23.645 80.685 ;
        RECT 24.060 80.525 25.015 80.695 ;
        RECT 25.185 80.295 25.475 81.130 ;
        RECT 46.755 81.055 46.925 82.015 ;
        RECT 47.095 81.675 48.400 81.845 ;
        RECT 49.485 81.765 49.805 82.695 ;
        RECT 81.315 82.220 81.605 83.385 ;
        RECT 82.020 82.245 82.230 83.385 ;
        RECT 85.520 83.335 87.350 83.505 ;
        RECT 89.430 83.345 91.270 83.515 ;
        RECT 82.400 82.235 82.730 83.215 ;
        RECT 82.000 81.825 82.330 82.065 ;
        RECT 47.095 81.225 47.340 81.675 ;
        RECT 47.510 81.305 48.060 81.505 ;
        RECT 48.230 81.475 48.400 81.675 ;
        RECT 49.175 81.595 49.805 81.765 ;
        RECT 48.230 81.305 48.605 81.475 ;
        RECT 48.775 81.055 49.005 81.555 ;
        RECT 46.295 80.315 46.585 81.040 ;
        RECT 46.755 80.885 49.005 81.055 ;
        RECT 46.805 80.315 47.135 80.705 ;
        RECT 47.305 80.565 47.475 80.885 ;
        RECT 49.175 80.715 49.345 81.595 ;
        RECT 47.645 80.315 47.975 80.705 ;
        RECT 48.390 80.545 49.345 80.715 ;
        RECT 49.515 80.315 49.805 81.150 ;
        RECT 81.315 80.835 81.605 81.560 ;
        RECT 82.000 80.835 82.230 81.655 ;
        RECT 82.500 81.635 82.730 82.235 ;
        RECT 85.860 82.195 86.070 83.335 ;
        RECT 86.240 82.185 86.570 83.165 ;
        RECT 85.840 81.775 86.170 82.015 ;
        RECT 82.400 81.005 82.730 81.635 ;
        RECT 81.230 80.665 83.060 80.835 ;
        RECT 85.840 80.785 86.070 81.605 ;
        RECT 86.340 81.585 86.570 82.185 ;
        RECT 86.975 82.170 87.265 83.335 ;
        RECT 89.515 82.180 89.805 83.345 ;
        RECT 90.230 82.205 90.440 83.345 ;
        RECT 92.960 83.335 94.780 83.505 ;
        RECT 90.610 82.195 90.940 83.175 ;
        RECT 93.300 82.195 93.510 83.335 ;
        RECT 90.210 81.785 90.540 82.025 ;
        RECT 86.240 80.955 86.570 81.585 ;
        RECT 86.975 80.785 87.265 81.510 ;
        RECT 89.515 80.795 89.805 81.520 ;
        RECT 90.210 80.795 90.440 81.615 ;
        RECT 90.710 81.595 90.940 82.195 ;
        RECT 93.680 82.185 94.010 83.165 ;
        RECT 93.280 81.775 93.610 82.015 ;
        RECT 90.610 80.965 90.940 81.595 ;
        RECT 85.520 80.615 87.350 80.785 ;
        RECT 89.430 80.625 91.270 80.795 ;
        RECT 93.280 80.785 93.510 81.605 ;
        RECT 93.780 81.585 94.010 82.185 ;
        RECT 94.405 82.170 94.695 83.335 ;
        RECT 96.800 83.285 98.630 83.455 ;
        RECT 101.170 83.295 102.960 83.465 ;
        RECT 106.780 83.305 108.540 83.475 ;
        RECT 97.140 82.145 97.350 83.285 ;
        RECT 97.520 82.135 97.850 83.115 ;
        RECT 97.120 81.725 97.450 81.965 ;
        RECT 93.680 80.955 94.010 81.585 ;
        RECT 94.405 80.785 94.695 81.510 ;
        RECT 92.960 80.615 94.780 80.785 ;
        RECT 97.120 80.735 97.350 81.555 ;
        RECT 97.620 81.535 97.850 82.135 ;
        RECT 98.255 82.120 98.545 83.285 ;
        RECT 101.510 82.155 101.720 83.295 ;
        RECT 101.890 82.145 102.220 83.125 ;
        RECT 101.490 81.735 101.820 81.975 ;
        RECT 97.520 80.905 97.850 81.535 ;
        RECT 98.255 80.735 98.545 81.460 ;
        RECT 101.490 80.745 101.720 81.565 ;
        RECT 101.990 81.545 102.220 82.145 ;
        RECT 102.585 82.130 102.875 83.295 ;
        RECT 107.120 82.165 107.330 83.305 ;
        RECT 107.500 82.155 107.830 83.135 ;
        RECT 107.100 81.745 107.430 81.985 ;
        RECT 101.890 80.915 102.220 81.545 ;
        RECT 102.585 80.745 102.875 81.470 ;
        RECT 107.100 80.755 107.330 81.575 ;
        RECT 107.600 81.555 107.830 82.155 ;
        RECT 108.165 82.140 108.455 83.305 ;
        RECT 110.620 83.255 112.430 83.425 ;
        RECT 114.990 83.265 116.760 83.435 ;
        RECT 110.960 82.115 111.170 83.255 ;
        RECT 111.340 82.105 111.670 83.085 ;
        RECT 110.940 81.695 111.270 81.935 ;
        RECT 107.500 80.925 107.830 81.555 ;
        RECT 108.165 80.755 108.455 81.480 ;
        RECT 96.800 80.565 98.630 80.735 ;
        RECT 101.170 80.575 102.960 80.745 ;
        RECT 106.780 80.585 108.540 80.755 ;
        RECT 110.940 80.705 111.170 81.525 ;
        RECT 111.440 81.505 111.670 82.105 ;
        RECT 112.055 82.090 112.345 83.255 ;
        RECT 115.330 82.125 115.540 83.265 ;
        RECT 115.710 82.115 116.040 83.095 ;
        RECT 115.310 81.705 115.640 81.945 ;
        RECT 111.340 80.875 111.670 81.505 ;
        RECT 112.055 80.705 112.345 81.430 ;
        RECT 115.310 80.715 115.540 81.535 ;
        RECT 115.810 81.515 116.040 82.115 ;
        RECT 116.385 82.100 116.675 83.265 ;
        RECT 115.710 80.885 116.040 81.515 ;
        RECT 116.385 80.715 116.675 81.440 ;
        RECT 110.620 80.535 112.430 80.705 ;
        RECT 114.990 80.545 116.760 80.715 ;
        RECT 21.880 80.125 25.560 80.295 ;
        RECT 46.210 80.145 49.890 80.315 ;
        RECT 22.380 79.125 25.130 79.295 ;
        RECT 46.710 79.145 49.460 79.315 ;
        RECT 22.465 77.960 22.755 79.125 ;
        RECT 23.115 78.455 23.395 79.125 ;
        RECT 23.565 78.235 23.865 78.785 ;
        RECT 24.065 78.405 24.395 79.125 ;
        RECT 24.585 78.405 25.045 78.955 ;
        RECT 33.040 78.575 36.720 78.745 ;
        RECT 22.930 77.815 23.195 78.175 ;
        RECT 23.565 78.065 24.505 78.235 ;
        RECT 24.335 77.815 24.505 78.065 ;
        RECT 22.930 77.565 23.605 77.815 ;
        RECT 23.825 77.565 24.165 77.815 ;
        RECT 24.335 77.485 24.625 77.815 ;
        RECT 24.335 77.395 24.505 77.485 ;
        RECT 22.465 76.575 22.755 77.300 ;
        RECT 23.115 77.205 24.505 77.395 ;
        RECT 23.115 76.845 23.445 77.205 ;
        RECT 24.795 77.035 25.045 78.405 ;
        RECT 33.130 78.195 33.465 78.575 ;
        RECT 24.065 76.575 24.315 77.035 ;
        RECT 24.485 76.745 25.045 77.035 ;
        RECT 33.125 76.705 33.365 78.015 ;
        RECT 33.635 77.605 33.885 78.405 ;
        RECT 34.105 77.855 34.435 78.575 ;
        RECT 34.620 77.605 34.870 78.405 ;
        RECT 35.335 77.775 35.665 78.575 ;
        RECT 35.835 78.145 36.175 78.405 ;
        RECT 33.535 77.435 35.725 77.605 ;
        RECT 22.380 76.405 25.130 76.575 ;
        RECT 33.535 76.525 33.705 77.435 ;
        RECT 35.410 77.265 35.725 77.435 ;
        RECT 28.750 76.075 31.510 76.245 ;
        RECT 33.210 76.195 33.705 76.525 ;
        RECT 33.925 76.300 34.275 77.265 ;
        RECT 34.455 76.295 34.755 77.265 ;
        RECT 34.935 76.295 35.215 77.265 ;
        RECT 35.410 77.015 35.740 77.265 ;
        RECT 29.035 75.405 29.315 76.075 ;
        RECT 21.930 75.025 25.610 75.195 ;
        RECT 29.485 75.185 29.785 75.735 ;
        RECT 29.985 75.355 30.315 76.075 ;
        RECT 30.505 75.355 30.965 75.905 ;
        RECT 22.015 73.860 22.305 75.025 ;
        RECT 22.475 74.175 22.855 74.855 ;
        RECT 23.445 74.175 23.615 75.025 ;
        RECT 23.785 74.345 24.115 74.855 ;
        RECT 24.285 74.515 24.455 75.025 ;
        RECT 24.625 74.345 25.025 74.855 ;
        RECT 23.785 74.175 25.025 74.345 ;
        RECT 22.475 73.215 22.645 74.175 ;
        RECT 22.815 73.835 24.120 74.005 ;
        RECT 25.205 73.925 25.525 74.855 ;
        RECT 28.850 74.765 29.115 75.125 ;
        RECT 29.485 75.015 30.425 75.185 ;
        RECT 30.255 74.765 30.425 75.015 ;
        RECT 28.850 74.515 29.525 74.765 ;
        RECT 29.745 74.515 30.085 74.765 ;
        RECT 30.255 74.435 30.545 74.765 ;
        RECT 30.255 74.345 30.425 74.435 ;
        RECT 22.815 73.385 23.060 73.835 ;
        RECT 23.230 73.465 23.780 73.665 ;
        RECT 23.950 73.635 24.120 73.835 ;
        RECT 24.895 73.755 25.525 73.925 ;
        RECT 29.035 74.155 30.425 74.345 ;
        RECT 29.035 73.795 29.365 74.155 ;
        RECT 30.715 73.985 30.965 75.355 ;
        RECT 31.135 74.910 31.425 76.075 ;
        RECT 35.395 76.025 35.665 76.825 ;
        RECT 35.915 76.745 36.175 78.145 ;
        RECT 36.345 77.410 36.635 78.575 ;
        RECT 46.795 77.980 47.085 79.145 ;
        RECT 47.445 78.475 47.725 79.145 ;
        RECT 47.895 78.255 48.195 78.805 ;
        RECT 48.395 78.425 48.725 79.145 ;
        RECT 48.915 78.425 49.375 78.975 ;
        RECT 57.370 78.595 61.050 78.765 ;
        RECT 47.260 77.835 47.525 78.195 ;
        RECT 47.895 78.085 48.835 78.255 ;
        RECT 48.665 77.835 48.835 78.085 ;
        RECT 47.260 77.585 47.935 77.835 ;
        RECT 48.155 77.585 48.495 77.835 ;
        RECT 48.665 77.505 48.955 77.835 ;
        RECT 48.665 77.415 48.835 77.505 ;
        RECT 35.835 76.235 36.175 76.745 ;
        RECT 36.345 76.025 36.635 76.750 ;
        RECT 46.795 76.595 47.085 77.320 ;
        RECT 47.445 77.225 48.835 77.415 ;
        RECT 47.445 76.865 47.775 77.225 ;
        RECT 49.125 77.055 49.375 78.425 ;
        RECT 57.460 78.215 57.795 78.595 ;
        RECT 48.395 76.595 48.645 77.055 ;
        RECT 48.815 76.765 49.375 77.055 ;
        RECT 57.455 76.725 57.695 78.035 ;
        RECT 57.965 77.625 58.215 78.425 ;
        RECT 58.435 77.875 58.765 78.595 ;
        RECT 58.950 77.625 59.200 78.425 ;
        RECT 59.665 77.795 59.995 78.595 ;
        RECT 60.165 78.165 60.505 78.425 ;
        RECT 57.865 77.455 60.055 77.625 ;
        RECT 46.710 76.425 49.460 76.595 ;
        RECT 57.865 76.545 58.035 77.455 ;
        RECT 59.740 77.285 60.055 77.455 ;
        RECT 53.080 76.095 55.840 76.265 ;
        RECT 57.540 76.215 58.035 76.545 ;
        RECT 58.255 76.320 58.605 77.285 ;
        RECT 58.785 76.315 59.085 77.285 ;
        RECT 59.265 76.315 59.545 77.285 ;
        RECT 59.740 77.035 60.070 77.285 ;
        RECT 33.040 75.855 36.720 76.025 ;
        RECT 53.365 75.425 53.645 76.095 ;
        RECT 46.260 75.045 49.940 75.215 ;
        RECT 53.815 75.205 54.115 75.755 ;
        RECT 54.315 75.375 54.645 76.095 ;
        RECT 54.835 75.375 55.295 75.925 ;
        RECT 23.950 73.465 24.325 73.635 ;
        RECT 24.495 73.215 24.725 73.715 ;
        RECT 22.015 72.475 22.305 73.200 ;
        RECT 22.475 73.045 24.725 73.215 ;
        RECT 22.525 72.475 22.855 72.865 ;
        RECT 23.025 72.725 23.195 73.045 ;
        RECT 24.895 72.875 25.065 73.755 ;
        RECT 29.985 73.525 30.235 73.985 ;
        RECT 30.405 73.695 30.965 73.985 ;
        RECT 31.135 73.525 31.425 74.250 ;
        RECT 46.345 73.880 46.635 75.045 ;
        RECT 46.805 74.195 47.185 74.875 ;
        RECT 47.775 74.195 47.945 75.045 ;
        RECT 48.115 74.365 48.445 74.875 ;
        RECT 48.615 74.535 48.785 75.045 ;
        RECT 48.955 74.365 49.355 74.875 ;
        RECT 48.115 74.195 49.355 74.365 ;
        RECT 28.750 73.355 31.510 73.525 ;
        RECT 23.365 72.475 23.695 72.865 ;
        RECT 24.110 72.705 25.065 72.875 ;
        RECT 25.235 72.475 25.525 73.310 ;
        RECT 46.805 73.235 46.975 74.195 ;
        RECT 47.145 73.855 48.450 74.025 ;
        RECT 49.535 73.945 49.855 74.875 ;
        RECT 53.180 74.785 53.445 75.145 ;
        RECT 53.815 75.035 54.755 75.205 ;
        RECT 54.585 74.785 54.755 75.035 ;
        RECT 53.180 74.535 53.855 74.785 ;
        RECT 54.075 74.535 54.415 74.785 ;
        RECT 54.585 74.455 54.875 74.785 ;
        RECT 54.585 74.365 54.755 74.455 ;
        RECT 47.145 73.405 47.390 73.855 ;
        RECT 47.560 73.485 48.110 73.685 ;
        RECT 48.280 73.655 48.450 73.855 ;
        RECT 49.225 73.775 49.855 73.945 ;
        RECT 53.365 74.175 54.755 74.365 ;
        RECT 53.365 73.815 53.695 74.175 ;
        RECT 55.045 74.005 55.295 75.375 ;
        RECT 55.465 74.930 55.755 76.095 ;
        RECT 59.725 76.045 59.995 76.845 ;
        RECT 60.245 76.765 60.505 78.165 ;
        RECT 60.675 77.430 60.965 78.595 ;
        RECT 60.165 76.255 60.505 76.765 ;
        RECT 60.675 76.045 60.965 76.770 ;
        RECT 57.370 75.875 61.050 76.045 ;
        RECT 48.280 73.485 48.655 73.655 ;
        RECT 48.825 73.235 49.055 73.735 ;
        RECT 46.345 72.495 46.635 73.220 ;
        RECT 46.805 73.065 49.055 73.235 ;
        RECT 46.855 72.495 47.185 72.885 ;
        RECT 47.355 72.745 47.525 73.065 ;
        RECT 49.225 72.895 49.395 73.775 ;
        RECT 54.315 73.545 54.565 74.005 ;
        RECT 54.735 73.715 55.295 74.005 ;
        RECT 55.465 73.545 55.755 74.270 ;
        RECT 117.420 74.075 127.540 74.245 ;
        RECT 53.080 73.375 55.840 73.545 ;
        RECT 117.595 73.405 117.765 73.905 ;
        RECT 117.935 73.695 118.265 74.075 ;
        RECT 118.435 73.735 119.965 73.905 ;
        RECT 118.435 73.575 118.605 73.735 ;
        RECT 118.955 73.405 119.125 73.565 ;
        RECT 47.695 72.495 48.025 72.885 ;
        RECT 48.440 72.725 49.395 72.895 ;
        RECT 49.565 72.495 49.855 73.330 ;
        RECT 117.595 73.235 119.125 73.405 ;
        RECT 119.295 73.395 119.625 73.565 ;
        RECT 119.295 73.065 119.465 73.395 ;
        RECT 119.795 73.235 119.965 73.735 ;
        RECT 120.135 73.065 120.485 73.905 ;
        RECT 120.655 73.695 120.985 74.075 ;
        RECT 121.245 73.735 122.255 73.905 ;
        RECT 21.930 72.305 25.610 72.475 ;
        RECT 46.260 72.325 49.940 72.495 ;
        RECT 117.570 72.435 117.915 73.055 ;
        RECT 118.225 72.435 118.660 73.055 ;
        RECT 118.830 72.895 119.465 73.065 ;
        RECT 118.830 72.375 119.000 72.895 ;
        RECT 119.680 72.835 120.485 73.065 ;
        RECT 119.680 72.725 120.040 72.835 ;
        RECT 119.500 72.545 120.040 72.725 ;
        RECT 117.595 72.075 118.605 72.245 ;
        RECT 117.595 71.700 117.765 72.075 ;
        RECT 117.935 71.525 118.265 71.905 ;
        RECT 118.435 71.865 118.605 72.075 ;
        RECT 118.830 72.205 119.120 72.375 ;
        RECT 118.830 72.035 119.170 72.205 ;
        RECT 119.340 71.865 119.510 72.200 ;
        RECT 119.680 71.870 120.040 72.545 ;
        RECT 120.685 72.435 120.985 73.435 ;
        RECT 121.245 73.225 121.415 73.735 ;
        RECT 121.585 73.055 121.915 73.565 ;
        RECT 122.085 73.525 122.255 73.735 ;
        RECT 122.480 73.695 122.810 74.075 ;
        RECT 122.980 73.525 123.150 73.905 ;
        RECT 123.400 73.695 123.750 74.075 ;
        RECT 123.920 73.575 124.105 73.905 ;
        RECT 122.085 73.355 123.150 73.525 ;
        RECT 121.155 72.885 121.915 73.055 ;
        RECT 121.155 72.360 121.325 72.885 ;
        RECT 121.710 72.705 121.880 72.715 ;
        RECT 121.495 72.545 121.880 72.705 ;
        RECT 121.495 72.535 121.825 72.545 ;
        RECT 122.220 72.495 122.465 73.115 ;
        RECT 122.670 72.495 123.000 73.115 ;
        RECT 123.475 72.435 123.765 73.115 ;
        RECT 123.935 72.715 124.105 73.575 ;
        RECT 124.400 73.575 124.610 73.905 ;
        RECT 124.780 73.735 126.065 73.905 ;
        RECT 124.780 73.695 125.110 73.735 ;
        RECT 123.935 72.545 124.225 72.715 ;
        RECT 121.155 72.285 121.470 72.360 ;
        RECT 118.435 71.695 119.510 71.865 ;
        RECT 120.220 71.525 120.510 72.245 ;
        RECT 120.800 71.865 120.970 72.235 ;
        RECT 121.140 72.035 121.470 72.285 ;
        RECT 121.640 72.325 121.810 72.365 ;
        RECT 121.640 72.155 123.160 72.325 ;
        RECT 121.640 72.035 121.810 72.155 ;
        RECT 122.045 71.865 122.400 71.905 ;
        RECT 120.800 71.695 122.400 71.865 ;
        RECT 122.570 71.525 122.740 71.985 ;
        RECT 122.915 71.735 123.160 72.155 ;
        RECT 123.935 72.095 124.105 72.545 ;
        RECT 124.400 72.375 124.570 73.575 ;
        RECT 125.265 73.425 125.595 73.565 ;
        RECT 124.810 73.195 125.595 73.425 ;
        RECT 125.895 73.275 126.065 73.735 ;
        RECT 126.235 73.695 126.565 74.075 ;
        RECT 124.400 72.205 124.640 72.375 ;
        RECT 123.430 71.525 123.760 71.905 ;
        RECT 123.930 71.765 124.105 72.095 ;
        RECT 124.810 72.025 124.980 73.195 ;
        RECT 125.895 73.105 126.545 73.275 ;
        RECT 125.610 72.545 126.065 72.715 ;
        RECT 125.390 72.365 125.800 72.375 ;
        RECT 125.390 72.205 125.805 72.365 ;
        RECT 126.375 72.325 126.545 73.105 ;
        RECT 125.630 72.035 125.805 72.205 ;
        RECT 125.975 72.155 126.545 72.325 ;
        RECT 124.450 71.855 124.980 72.025 ;
        RECT 125.150 71.865 125.320 72.025 ;
        RECT 125.975 71.865 126.145 72.155 ;
        RECT 124.450 71.695 124.620 71.855 ;
        RECT 125.150 71.695 126.145 71.865 ;
        RECT 126.315 71.525 126.485 71.985 ;
        RECT 126.735 71.695 126.995 73.905 ;
        RECT 127.165 72.910 127.455 74.075 ;
        RECT 127.165 71.525 127.455 72.250 ;
        RECT 22.430 71.305 25.180 71.475 ;
        RECT 22.515 70.140 22.805 71.305 ;
        RECT 23.165 70.635 23.445 71.305 ;
        RECT 23.615 70.415 23.915 70.965 ;
        RECT 24.115 70.585 24.445 71.305 ;
        RECT 28.660 71.245 32.340 71.415 ;
        RECT 24.635 70.585 25.095 71.135 ;
        RECT 22.980 69.995 23.245 70.355 ;
        RECT 23.615 70.245 24.555 70.415 ;
        RECT 24.385 69.995 24.555 70.245 ;
        RECT 22.980 69.745 23.655 69.995 ;
        RECT 23.875 69.745 24.215 69.995 ;
        RECT 24.385 69.665 24.675 69.995 ;
        RECT 24.385 69.575 24.555 69.665 ;
        RECT 22.515 68.755 22.805 69.480 ;
        RECT 23.165 69.385 24.555 69.575 ;
        RECT 23.165 69.025 23.495 69.385 ;
        RECT 24.845 69.215 25.095 70.585 ;
        RECT 28.745 70.080 29.035 71.245 ;
        RECT 29.210 70.865 29.545 71.245 ;
        RECT 24.115 68.755 24.365 69.215 ;
        RECT 24.535 68.925 25.095 69.215 ;
        RECT 22.430 68.585 25.180 68.755 ;
        RECT 28.745 68.695 29.035 69.420 ;
        RECT 29.205 69.375 29.445 70.685 ;
        RECT 29.715 70.275 29.965 71.075 ;
        RECT 30.185 70.525 30.515 71.245 ;
        RECT 30.700 70.275 30.950 71.075 ;
        RECT 31.415 70.445 31.745 71.245 ;
        RECT 38.610 71.165 41.830 71.335 ;
        RECT 46.750 71.325 49.510 71.495 ;
        RECT 31.915 70.815 32.255 71.075 ;
        RECT 29.615 70.105 31.805 70.275 ;
        RECT 29.615 69.195 29.785 70.105 ;
        RECT 31.490 69.935 31.805 70.105 ;
        RECT 29.290 68.865 29.785 69.195 ;
        RECT 30.005 68.970 30.355 69.935 ;
        RECT 30.535 68.965 30.835 69.935 ;
        RECT 31.015 68.965 31.295 69.935 ;
        RECT 31.490 69.685 31.820 69.935 ;
        RECT 31.475 68.695 31.745 69.495 ;
        RECT 31.995 69.415 32.255 70.815 ;
        RECT 38.700 70.655 40.355 70.945 ;
        RECT 38.700 70.315 40.290 70.485 ;
        RECT 40.525 70.365 40.805 71.165 ;
        RECT 38.700 70.025 39.020 70.315 ;
        RECT 40.120 70.195 40.290 70.315 ;
        RECT 31.915 68.905 32.255 69.415 ;
        RECT 33.970 69.375 36.710 69.545 ;
        RECT 28.660 68.525 32.340 68.695 ;
        RECT 34.240 68.405 34.630 68.580 ;
        RECT 35.115 68.575 35.445 69.375 ;
        RECT 35.615 68.585 36.150 69.205 ;
        RECT 34.240 68.235 35.665 68.405 ;
        RECT 34.115 67.505 34.470 68.065 ;
        RECT 34.640 67.335 34.810 68.235 ;
        RECT 34.980 67.505 35.245 68.065 ;
        RECT 35.495 67.735 35.665 68.235 ;
        RECT 35.835 67.565 36.150 68.585 ;
        RECT 36.335 68.210 36.625 69.375 ;
        RECT 38.700 69.285 39.050 69.855 ;
        RECT 39.220 69.525 39.930 70.145 ;
        RECT 40.120 70.025 40.845 70.195 ;
        RECT 41.015 70.025 41.285 70.995 ;
        RECT 40.675 69.855 40.845 70.025 ;
        RECT 40.100 69.525 40.505 69.855 ;
        RECT 40.675 69.525 40.945 69.855 ;
        RECT 40.675 69.355 40.845 69.525 ;
        RECT 39.235 69.185 40.845 69.355 ;
        RECT 41.115 69.290 41.285 70.025 ;
        RECT 41.455 70.000 41.745 71.165 ;
        RECT 46.835 70.160 47.125 71.325 ;
        RECT 47.495 70.655 47.775 71.325 ;
        RECT 47.945 70.435 48.245 70.985 ;
        RECT 48.445 70.605 48.775 71.325 ;
        RECT 52.990 71.265 56.670 71.435 ;
        RECT 117.420 71.355 127.540 71.525 ;
        RECT 48.965 70.605 49.425 71.155 ;
        RECT 47.310 70.015 47.575 70.375 ;
        RECT 47.945 70.265 48.885 70.435 ;
        RECT 48.715 70.015 48.885 70.265 ;
        RECT 47.310 69.765 47.985 70.015 ;
        RECT 48.205 69.765 48.545 70.015 ;
        RECT 48.715 69.685 49.005 70.015 ;
        RECT 48.715 69.595 48.885 69.685 ;
        RECT 38.705 68.615 39.035 69.115 ;
        RECT 39.235 68.835 39.405 69.185 ;
        RECT 39.605 68.615 39.935 69.015 ;
        RECT 40.105 68.835 40.275 69.185 ;
        RECT 40.445 68.615 40.825 69.015 ;
        RECT 41.015 68.945 41.285 69.290 ;
        RECT 41.455 68.615 41.745 69.340 ;
        RECT 46.835 68.775 47.125 69.500 ;
        RECT 47.495 69.405 48.885 69.595 ;
        RECT 47.495 69.045 47.825 69.405 ;
        RECT 49.175 69.235 49.425 70.605 ;
        RECT 53.075 70.100 53.365 71.265 ;
        RECT 53.540 70.885 53.875 71.265 ;
        RECT 48.445 68.775 48.695 69.235 ;
        RECT 48.865 68.945 49.425 69.235 ;
        RECT 38.610 68.445 41.830 68.615 ;
        RECT 46.750 68.605 49.510 68.775 ;
        RECT 53.075 68.715 53.365 69.440 ;
        RECT 53.535 69.395 53.775 70.705 ;
        RECT 54.045 70.295 54.295 71.095 ;
        RECT 54.515 70.545 54.845 71.265 ;
        RECT 55.030 70.295 55.280 71.095 ;
        RECT 55.745 70.465 56.075 71.265 ;
        RECT 62.940 71.185 66.160 71.355 ;
        RECT 56.245 70.835 56.585 71.095 ;
        RECT 53.945 70.125 56.135 70.295 ;
        RECT 53.945 69.215 54.115 70.125 ;
        RECT 55.820 69.955 56.135 70.125 ;
        RECT 53.620 68.885 54.115 69.215 ;
        RECT 54.335 68.990 54.685 69.955 ;
        RECT 54.865 68.985 55.165 69.955 ;
        RECT 55.345 68.985 55.625 69.955 ;
        RECT 55.820 69.705 56.150 69.955 ;
        RECT 55.805 68.715 56.075 69.515 ;
        RECT 56.325 69.435 56.585 70.835 ;
        RECT 63.030 70.675 64.685 70.965 ;
        RECT 63.030 70.335 64.620 70.505 ;
        RECT 64.855 70.385 65.135 71.185 ;
        RECT 63.030 70.045 63.350 70.335 ;
        RECT 64.450 70.215 64.620 70.335 ;
        RECT 56.245 68.925 56.585 69.435 ;
        RECT 58.300 69.395 61.050 69.565 ;
        RECT 52.990 68.545 56.670 68.715 ;
        RECT 58.570 68.425 58.960 68.600 ;
        RECT 59.445 68.595 59.775 69.395 ;
        RECT 59.945 68.605 60.480 69.225 ;
        RECT 58.570 68.255 59.995 68.425 ;
        RECT 29.280 67.035 32.040 67.205 ;
        RECT 21.890 66.685 25.570 66.855 ;
        RECT 21.975 65.520 22.265 66.685 ;
        RECT 22.435 65.835 22.815 66.515 ;
        RECT 23.405 65.835 23.575 66.685 ;
        RECT 23.745 66.005 24.075 66.515 ;
        RECT 24.245 66.175 24.415 66.685 ;
        RECT 24.585 66.005 24.985 66.515 ;
        RECT 23.745 65.835 24.985 66.005 ;
        RECT 22.435 64.875 22.605 65.835 ;
        RECT 22.775 65.495 24.080 65.665 ;
        RECT 25.165 65.585 25.485 66.515 ;
        RECT 29.365 65.870 29.655 67.035 ;
        RECT 29.825 66.480 30.430 67.035 ;
        RECT 30.605 66.525 31.085 66.865 ;
        RECT 30.730 66.490 30.910 66.525 ;
        RECT 31.255 66.490 31.510 67.035 ;
        RECT 29.825 66.380 30.440 66.480 ;
        RECT 30.255 66.355 30.440 66.380 ;
        RECT 29.825 65.760 30.085 66.210 ;
        RECT 30.255 66.110 30.585 66.355 ;
        RECT 30.755 66.035 31.510 66.285 ;
        RECT 31.680 66.165 31.955 66.865 ;
        RECT 34.220 66.825 34.460 67.335 ;
        RECT 34.640 67.005 34.920 67.335 ;
        RECT 35.150 66.825 35.365 67.335 ;
        RECT 35.535 66.995 36.150 67.565 ;
        RECT 36.335 66.825 36.625 67.550 ;
        RECT 58.445 67.525 58.800 68.085 ;
        RECT 58.970 67.355 59.140 68.255 ;
        RECT 59.310 67.525 59.575 68.085 ;
        RECT 59.825 67.755 59.995 68.255 ;
        RECT 60.165 67.585 60.480 68.605 ;
        RECT 60.675 68.230 60.965 69.395 ;
        RECT 63.030 69.305 63.380 69.875 ;
        RECT 63.550 69.545 64.260 70.165 ;
        RECT 64.450 70.045 65.175 70.215 ;
        RECT 65.345 70.045 65.615 71.015 ;
        RECT 65.005 69.875 65.175 70.045 ;
        RECT 64.430 69.545 64.835 69.875 ;
        RECT 65.005 69.545 65.275 69.875 ;
        RECT 65.005 69.375 65.175 69.545 ;
        RECT 63.565 69.205 65.175 69.375 ;
        RECT 65.445 69.310 65.615 70.045 ;
        RECT 65.785 70.020 66.075 71.185 ;
        RECT 63.035 68.635 63.365 69.135 ;
        RECT 63.565 68.855 63.735 69.205 ;
        RECT 63.935 68.635 64.265 69.035 ;
        RECT 64.435 68.855 64.605 69.205 ;
        RECT 64.775 68.635 65.155 69.035 ;
        RECT 65.345 68.965 65.615 69.310 ;
        RECT 65.785 68.635 66.075 69.360 ;
        RECT 62.940 68.465 66.160 68.635 ;
        RECT 53.610 67.055 56.370 67.225 ;
        RECT 33.970 66.655 36.710 66.825 ;
        RECT 46.220 66.705 49.900 66.875 ;
        RECT 30.740 66.000 31.510 66.035 ;
        RECT 30.725 65.990 31.510 66.000 ;
        RECT 30.720 65.975 31.615 65.990 ;
        RECT 30.700 65.960 31.615 65.975 ;
        RECT 30.680 65.950 31.615 65.960 ;
        RECT 30.655 65.940 31.615 65.950 ;
        RECT 30.585 65.910 31.615 65.940 ;
        RECT 30.565 65.880 31.615 65.910 ;
        RECT 30.545 65.850 31.615 65.880 ;
        RECT 30.515 65.825 31.615 65.850 ;
        RECT 30.480 65.790 31.615 65.825 ;
        RECT 30.450 65.785 31.615 65.790 ;
        RECT 30.450 65.780 30.840 65.785 ;
        RECT 30.450 65.770 30.815 65.780 ;
        RECT 30.450 65.765 30.800 65.770 ;
        RECT 30.450 65.760 30.785 65.765 ;
        RECT 29.825 65.755 30.785 65.760 ;
        RECT 29.825 65.745 30.775 65.755 ;
        RECT 29.825 65.740 30.765 65.745 ;
        RECT 29.825 65.730 30.755 65.740 ;
        RECT 29.825 65.720 30.750 65.730 ;
        RECT 29.825 65.715 30.745 65.720 ;
        RECT 29.825 65.700 30.735 65.715 ;
        RECT 29.825 65.685 30.730 65.700 ;
        RECT 29.825 65.660 30.720 65.685 ;
        RECT 29.825 65.590 30.715 65.660 ;
        RECT 22.775 65.045 23.020 65.495 ;
        RECT 23.190 65.125 23.740 65.325 ;
        RECT 23.910 65.295 24.080 65.495 ;
        RECT 24.855 65.415 25.485 65.585 ;
        RECT 23.910 65.125 24.285 65.295 ;
        RECT 24.455 64.875 24.685 65.375 ;
        RECT 21.975 64.135 22.265 64.860 ;
        RECT 22.435 64.705 24.685 64.875 ;
        RECT 22.485 64.135 22.815 64.525 ;
        RECT 22.985 64.385 23.155 64.705 ;
        RECT 24.855 64.535 25.025 65.415 ;
        RECT 23.325 64.135 23.655 64.525 ;
        RECT 24.070 64.365 25.025 64.535 ;
        RECT 25.195 64.135 25.485 64.970 ;
        RECT 29.365 64.485 29.655 65.210 ;
        RECT 29.825 65.035 30.375 65.420 ;
        RECT 30.545 64.865 30.715 65.590 ;
        RECT 29.825 64.695 30.715 64.865 ;
        RECT 30.885 65.190 31.215 65.615 ;
        RECT 31.385 65.390 31.615 65.785 ;
        RECT 30.885 65.160 31.160 65.190 ;
        RECT 30.885 64.705 31.105 65.160 ;
        RECT 31.785 65.135 31.955 66.165 ;
        RECT 46.305 65.540 46.595 66.705 ;
        RECT 46.765 65.855 47.145 66.535 ;
        RECT 47.735 65.855 47.905 66.705 ;
        RECT 48.075 66.025 48.405 66.535 ;
        RECT 48.575 66.195 48.745 66.705 ;
        RECT 48.915 66.025 49.315 66.535 ;
        RECT 48.075 65.855 49.315 66.025 ;
        RECT 31.275 64.485 31.525 65.025 ;
        RECT 31.695 64.655 31.955 65.135 ;
        RECT 46.765 64.895 46.935 65.855 ;
        RECT 47.105 65.515 48.410 65.685 ;
        RECT 49.495 65.605 49.815 66.535 ;
        RECT 53.695 65.890 53.985 67.055 ;
        RECT 54.155 66.500 54.760 67.055 ;
        RECT 54.935 66.545 55.415 66.885 ;
        RECT 55.060 66.510 55.240 66.545 ;
        RECT 55.585 66.510 55.840 67.055 ;
        RECT 54.155 66.400 54.770 66.500 ;
        RECT 54.585 66.375 54.770 66.400 ;
        RECT 54.155 65.780 54.415 66.230 ;
        RECT 54.585 66.130 54.915 66.375 ;
        RECT 55.085 66.055 55.840 66.305 ;
        RECT 56.010 66.185 56.285 66.885 ;
        RECT 58.550 66.845 58.790 67.355 ;
        RECT 58.970 67.025 59.250 67.355 ;
        RECT 59.480 66.845 59.695 67.355 ;
        RECT 59.865 67.015 60.480 67.585 ;
        RECT 60.675 66.845 60.965 67.570 ;
        RECT 58.300 66.675 61.050 66.845 ;
        RECT 55.070 66.020 55.840 66.055 ;
        RECT 55.055 66.010 55.840 66.020 ;
        RECT 55.050 65.995 55.945 66.010 ;
        RECT 55.030 65.980 55.945 65.995 ;
        RECT 55.010 65.970 55.945 65.980 ;
        RECT 54.985 65.960 55.945 65.970 ;
        RECT 54.915 65.930 55.945 65.960 ;
        RECT 54.895 65.900 55.945 65.930 ;
        RECT 54.875 65.870 55.945 65.900 ;
        RECT 54.845 65.845 55.945 65.870 ;
        RECT 54.810 65.810 55.945 65.845 ;
        RECT 54.780 65.805 55.945 65.810 ;
        RECT 54.780 65.800 55.170 65.805 ;
        RECT 54.780 65.790 55.145 65.800 ;
        RECT 54.780 65.785 55.130 65.790 ;
        RECT 54.780 65.780 55.115 65.785 ;
        RECT 54.155 65.775 55.115 65.780 ;
        RECT 54.155 65.765 55.105 65.775 ;
        RECT 54.155 65.760 55.095 65.765 ;
        RECT 54.155 65.750 55.085 65.760 ;
        RECT 54.155 65.740 55.080 65.750 ;
        RECT 54.155 65.735 55.075 65.740 ;
        RECT 54.155 65.720 55.065 65.735 ;
        RECT 54.155 65.705 55.060 65.720 ;
        RECT 54.155 65.680 55.050 65.705 ;
        RECT 54.155 65.610 55.045 65.680 ;
        RECT 47.105 65.065 47.350 65.515 ;
        RECT 47.520 65.145 48.070 65.345 ;
        RECT 48.240 65.315 48.410 65.515 ;
        RECT 49.185 65.435 49.815 65.605 ;
        RECT 48.240 65.145 48.615 65.315 ;
        RECT 48.785 64.895 49.015 65.395 ;
        RECT 29.280 64.315 32.040 64.485 ;
        RECT 46.305 64.155 46.595 64.880 ;
        RECT 46.765 64.725 49.015 64.895 ;
        RECT 46.815 64.155 47.145 64.545 ;
        RECT 47.315 64.405 47.485 64.725 ;
        RECT 49.185 64.555 49.355 65.435 ;
        RECT 47.655 64.155 47.985 64.545 ;
        RECT 48.400 64.385 49.355 64.555 ;
        RECT 49.525 64.155 49.815 64.990 ;
        RECT 53.695 64.505 53.985 65.230 ;
        RECT 54.155 65.055 54.705 65.440 ;
        RECT 54.875 64.885 55.045 65.610 ;
        RECT 54.155 64.715 55.045 64.885 ;
        RECT 55.215 65.210 55.545 65.635 ;
        RECT 55.715 65.410 55.945 65.805 ;
        RECT 55.215 65.180 55.490 65.210 ;
        RECT 55.215 64.725 55.435 65.180 ;
        RECT 56.115 65.155 56.285 66.185 ;
        RECT 55.605 64.505 55.855 65.045 ;
        RECT 56.025 64.675 56.285 65.155 ;
        RECT 53.610 64.335 56.370 64.505 ;
        RECT 21.890 63.965 25.570 64.135 ;
        RECT 46.220 63.985 49.900 64.155 ;
        RECT 22.390 62.965 25.140 63.135 ;
        RECT 46.710 62.985 49.470 63.155 ;
        RECT 22.475 61.800 22.765 62.965 ;
        RECT 23.125 62.295 23.405 62.965 ;
        RECT 23.575 62.075 23.875 62.625 ;
        RECT 24.075 62.245 24.405 62.965 ;
        RECT 24.595 62.245 25.055 62.795 ;
        RECT 22.940 61.655 23.205 62.015 ;
        RECT 23.575 61.905 24.515 62.075 ;
        RECT 24.345 61.655 24.515 61.905 ;
        RECT 22.940 61.405 23.615 61.655 ;
        RECT 23.835 61.405 24.175 61.655 ;
        RECT 24.345 61.325 24.635 61.655 ;
        RECT 24.345 61.235 24.515 61.325 ;
        RECT 22.475 60.415 22.765 61.140 ;
        RECT 23.125 61.045 24.515 61.235 ;
        RECT 23.125 60.685 23.455 61.045 ;
        RECT 24.805 60.875 25.055 62.245 ;
        RECT 29.260 61.935 32.020 62.105 ;
        RECT 24.075 60.415 24.325 60.875 ;
        RECT 24.495 60.585 25.055 60.875 ;
        RECT 29.345 60.770 29.635 61.935 ;
        RECT 30.005 61.265 30.285 61.935 ;
        RECT 30.455 61.045 30.755 61.595 ;
        RECT 30.955 61.215 31.285 61.935 ;
        RECT 46.795 61.820 47.085 62.985 ;
        RECT 47.455 62.315 47.735 62.985 ;
        RECT 47.905 62.095 48.205 62.645 ;
        RECT 48.405 62.265 48.735 62.985 ;
        RECT 48.925 62.265 49.385 62.815 ;
        RECT 31.475 61.215 31.935 61.765 ;
        RECT 47.270 61.675 47.535 62.035 ;
        RECT 47.905 61.925 48.845 62.095 ;
        RECT 48.675 61.675 48.845 61.925 ;
        RECT 47.270 61.425 47.945 61.675 ;
        RECT 48.165 61.425 48.505 61.675 ;
        RECT 48.675 61.345 48.965 61.675 ;
        RECT 48.675 61.255 48.845 61.345 ;
        RECT 29.820 60.625 30.085 60.985 ;
        RECT 30.455 60.875 31.395 61.045 ;
        RECT 31.225 60.625 31.395 60.875 ;
        RECT 22.390 60.245 25.140 60.415 ;
        RECT 29.820 60.375 30.495 60.625 ;
        RECT 30.715 60.375 31.055 60.625 ;
        RECT 31.225 60.295 31.515 60.625 ;
        RECT 31.225 60.205 31.395 60.295 ;
        RECT 29.345 59.385 29.635 60.110 ;
        RECT 30.005 60.015 31.395 60.205 ;
        RECT 30.005 59.655 30.335 60.015 ;
        RECT 31.685 59.845 31.935 61.215 ;
        RECT 46.795 60.435 47.085 61.160 ;
        RECT 47.455 61.065 48.845 61.255 ;
        RECT 47.455 60.705 47.785 61.065 ;
        RECT 49.135 60.895 49.385 62.265 ;
        RECT 53.590 61.955 56.350 62.125 ;
        RECT 48.405 60.435 48.655 60.895 ;
        RECT 48.825 60.605 49.385 60.895 ;
        RECT 53.675 60.790 53.965 61.955 ;
        RECT 54.335 61.285 54.615 61.955 ;
        RECT 54.785 61.065 55.085 61.615 ;
        RECT 55.285 61.235 55.615 61.955 ;
        RECT 55.805 61.235 56.265 61.785 ;
        RECT 54.150 60.645 54.415 61.005 ;
        RECT 54.785 60.895 55.725 61.065 ;
        RECT 55.555 60.645 55.725 60.895 ;
        RECT 46.710 60.265 49.470 60.435 ;
        RECT 54.150 60.395 54.825 60.645 ;
        RECT 55.045 60.395 55.385 60.645 ;
        RECT 55.555 60.315 55.845 60.645 ;
        RECT 55.555 60.225 55.725 60.315 ;
        RECT 30.955 59.385 31.205 59.845 ;
        RECT 31.375 59.555 31.935 59.845 ;
        RECT 53.675 59.405 53.965 60.130 ;
        RECT 54.335 60.035 55.725 60.225 ;
        RECT 54.335 59.675 54.665 60.035 ;
        RECT 56.015 59.865 56.265 61.235 ;
        RECT 55.285 59.405 55.535 59.865 ;
        RECT 55.705 59.575 56.265 59.865 ;
        RECT 29.260 59.215 32.020 59.385 ;
        RECT 53.590 59.235 56.350 59.405 ;
        RECT 21.940 58.865 25.620 59.035 ;
        RECT 46.270 58.885 49.950 59.055 ;
        RECT 22.025 57.700 22.315 58.865 ;
        RECT 22.485 58.015 22.865 58.695 ;
        RECT 23.455 58.015 23.625 58.865 ;
        RECT 23.795 58.185 24.125 58.695 ;
        RECT 24.295 58.355 24.465 58.865 ;
        RECT 24.635 58.185 25.035 58.695 ;
        RECT 23.795 58.015 25.035 58.185 ;
        RECT 22.485 57.055 22.655 58.015 ;
        RECT 22.825 57.675 24.130 57.845 ;
        RECT 25.215 57.765 25.535 58.695 ;
        RECT 22.825 57.225 23.070 57.675 ;
        RECT 23.240 57.305 23.790 57.505 ;
        RECT 23.960 57.475 24.130 57.675 ;
        RECT 24.905 57.595 25.535 57.765 ;
        RECT 46.355 57.720 46.645 58.885 ;
        RECT 46.815 58.035 47.195 58.715 ;
        RECT 47.785 58.035 47.955 58.885 ;
        RECT 48.125 58.205 48.455 58.715 ;
        RECT 48.625 58.375 48.795 58.885 ;
        RECT 48.965 58.205 49.365 58.715 ;
        RECT 48.125 58.035 49.365 58.205 ;
        RECT 23.960 57.305 24.335 57.475 ;
        RECT 24.505 57.055 24.735 57.555 ;
        RECT 22.025 56.315 22.315 57.040 ;
        RECT 22.485 56.885 24.735 57.055 ;
        RECT 22.535 56.315 22.865 56.705 ;
        RECT 23.035 56.565 23.205 56.885 ;
        RECT 24.905 56.715 25.075 57.595 ;
        RECT 23.375 56.315 23.705 56.705 ;
        RECT 24.120 56.545 25.075 56.715 ;
        RECT 25.245 56.315 25.535 57.150 ;
        RECT 46.815 57.075 46.985 58.035 ;
        RECT 47.155 57.695 48.460 57.865 ;
        RECT 49.545 57.785 49.865 58.715 ;
        RECT 47.155 57.245 47.400 57.695 ;
        RECT 47.570 57.325 48.120 57.525 ;
        RECT 48.290 57.495 48.460 57.695 ;
        RECT 49.235 57.615 49.865 57.785 ;
        RECT 48.290 57.325 48.665 57.495 ;
        RECT 48.835 57.075 49.065 57.575 ;
        RECT 46.355 56.335 46.645 57.060 ;
        RECT 46.815 56.905 49.065 57.075 ;
        RECT 46.865 56.335 47.195 56.725 ;
        RECT 47.365 56.585 47.535 56.905 ;
        RECT 49.235 56.735 49.405 57.615 ;
        RECT 47.705 56.335 48.035 56.725 ;
        RECT 48.450 56.565 49.405 56.735 ;
        RECT 49.575 56.335 49.865 57.170 ;
        RECT 21.940 56.145 25.620 56.315 ;
        RECT 46.270 56.165 49.950 56.335 ;
        RECT 22.430 55.145 25.190 55.315 ;
        RECT 46.760 55.165 49.520 55.335 ;
        RECT 22.515 53.980 22.805 55.145 ;
        RECT 23.175 54.475 23.455 55.145 ;
        RECT 23.625 54.255 23.925 54.805 ;
        RECT 24.125 54.425 24.455 55.145 ;
        RECT 24.645 54.425 25.105 54.975 ;
        RECT 22.990 53.835 23.255 54.195 ;
        RECT 23.625 54.085 24.565 54.255 ;
        RECT 24.395 53.835 24.565 54.085 ;
        RECT 22.990 53.585 23.665 53.835 ;
        RECT 23.885 53.585 24.225 53.835 ;
        RECT 24.395 53.505 24.685 53.835 ;
        RECT 24.395 53.415 24.565 53.505 ;
        RECT 22.515 52.595 22.805 53.320 ;
        RECT 23.175 53.225 24.565 53.415 ;
        RECT 23.175 52.865 23.505 53.225 ;
        RECT 24.855 53.055 25.105 54.425 ;
        RECT 46.845 54.000 47.135 55.165 ;
        RECT 47.505 54.495 47.785 55.165 ;
        RECT 47.955 54.275 48.255 54.825 ;
        RECT 48.455 54.445 48.785 55.165 ;
        RECT 48.975 54.445 49.435 54.995 ;
        RECT 47.320 53.855 47.585 54.215 ;
        RECT 47.955 54.105 48.895 54.275 ;
        RECT 48.725 53.855 48.895 54.105 ;
        RECT 47.320 53.605 47.995 53.855 ;
        RECT 48.215 53.605 48.555 53.855 ;
        RECT 48.725 53.525 49.015 53.855 ;
        RECT 48.725 53.435 48.895 53.525 ;
        RECT 24.125 52.595 24.375 53.055 ;
        RECT 24.545 52.765 25.105 53.055 ;
        RECT 46.845 52.615 47.135 53.340 ;
        RECT 47.505 53.245 48.895 53.435 ;
        RECT 47.505 52.885 47.835 53.245 ;
        RECT 49.185 53.075 49.435 54.445 ;
        RECT 48.455 52.615 48.705 53.075 ;
        RECT 48.875 52.785 49.435 53.075 ;
        RECT 22.430 52.425 25.190 52.595 ;
        RECT 46.760 52.445 49.520 52.615 ;
        RECT 30.560 32.915 32.350 33.085 ;
        RECT 30.890 32.115 31.220 32.745 ;
        RECT 30.890 31.515 31.120 32.115 ;
        RECT 31.390 32.095 31.620 32.915 ;
        RECT 31.975 32.190 32.265 32.915 ;
        RECT 31.290 31.685 31.620 31.925 ;
        RECT 30.890 30.535 31.220 31.515 ;
        RECT 31.390 30.365 31.600 31.505 ;
        RECT 31.975 30.365 32.265 31.530 ;
        RECT 30.560 30.195 32.350 30.365 ;
        RECT 49.640 29.755 57.450 29.925 ;
        RECT 49.725 29.030 50.015 29.755 ;
        RECT 50.210 29.030 50.610 29.585 ;
        RECT 50.855 29.395 51.185 29.755 ;
        RECT 51.355 29.335 52.365 29.585 ;
        RECT 51.355 29.225 51.525 29.335 ;
        RECT 52.195 29.245 52.365 29.335 ;
        RECT 50.785 29.055 51.525 29.225 ;
        RECT 52.700 29.225 52.870 29.585 ;
        RECT 53.040 29.395 53.370 29.755 ;
        RECT 53.540 29.225 53.710 29.585 ;
        RECT 53.880 29.350 54.210 29.755 ;
        RECT 8.730 27.655 16.540 27.825 ;
        RECT 8.815 26.930 9.105 27.655 ;
        RECT 9.300 26.930 9.700 27.485 ;
        RECT 9.945 27.295 10.275 27.655 ;
        RECT 10.445 27.235 11.455 27.485 ;
        RECT 10.445 27.125 10.615 27.235 ;
        RECT 11.285 27.145 11.455 27.235 ;
        RECT 9.875 26.955 10.615 27.125 ;
        RECT 11.790 27.125 11.960 27.485 ;
        RECT 12.130 27.295 12.460 27.655 ;
        RECT 12.630 27.125 12.800 27.485 ;
        RECT 12.970 27.250 13.300 27.655 ;
        RECT 8.815 25.105 9.105 26.270 ;
        RECT 9.300 26.255 9.630 26.930 ;
        RECT 9.875 26.745 10.045 26.955 ;
        RECT 9.800 26.415 10.045 26.745 ;
        RECT 11.080 26.785 11.575 26.975 ;
        RECT 11.790 26.955 12.800 27.125 ;
        RECT 13.570 27.125 13.740 27.485 ;
        RECT 13.910 27.295 14.240 27.655 ;
        RECT 14.410 27.125 14.580 27.485 ;
        RECT 13.570 26.955 14.580 27.125 ;
        RECT 14.830 27.105 15.430 27.485 ;
        RECT 15.695 27.275 16.025 27.655 ;
        RECT 19.400 27.615 27.210 27.785 ;
        RECT 29.150 27.615 36.970 27.785 ;
        RECT 39.160 27.645 46.980 27.815 ;
        RECT 14.830 26.935 16.025 27.105 ;
        RECT 14.830 26.805 15.070 26.935 ;
        RECT 10.215 26.465 10.655 26.705 ;
        RECT 11.080 26.615 11.745 26.785 ;
        RECT 11.915 26.465 12.290 26.785 ;
        RECT 12.585 26.490 13.750 26.775 ;
        RECT 15.855 26.745 16.025 26.935 ;
        RECT 16.195 26.910 16.455 27.485 ;
        RECT 9.300 25.275 9.700 26.255 ;
        RECT 9.875 25.805 10.045 26.415 ;
        RECT 10.485 25.975 10.905 26.295 ;
        RECT 12.585 26.225 12.755 26.490 ;
        RECT 11.135 26.055 12.755 26.225 ;
        RECT 9.875 25.635 10.540 25.805 ;
        RECT 11.135 25.785 11.385 26.055 ;
        RECT 12.980 25.975 13.340 26.305 ;
        RECT 13.580 26.145 13.750 26.490 ;
        RECT 13.920 26.380 14.310 26.710 ;
        RECT 14.500 26.465 14.870 26.635 ;
        RECT 15.300 26.465 15.630 26.745 ;
        RECT 14.500 26.145 14.670 26.465 ;
        RECT 15.460 26.415 15.630 26.465 ;
        RECT 15.855 26.415 16.110 26.745 ;
        RECT 13.580 25.975 14.670 26.145 ;
        RECT 14.840 25.860 15.240 26.295 ;
        RECT 15.855 26.115 16.025 26.415 ;
        RECT 16.280 26.255 16.455 26.910 ;
        RECT 19.485 26.890 19.775 27.615 ;
        RECT 19.970 26.890 20.370 27.445 ;
        RECT 20.615 27.255 20.945 27.615 ;
        RECT 21.115 27.195 22.125 27.445 ;
        RECT 21.115 27.085 21.285 27.195 ;
        RECT 21.955 27.105 22.125 27.195 ;
        RECT 20.545 26.915 21.285 27.085 ;
        RECT 22.460 27.085 22.630 27.445 ;
        RECT 22.800 27.255 23.130 27.615 ;
        RECT 23.300 27.085 23.470 27.445 ;
        RECT 23.640 27.210 23.970 27.615 ;
        RECT 10.370 25.615 10.540 25.635 ;
        RECT 11.790 25.635 12.800 25.805 ;
        RECT 9.870 25.105 10.200 25.465 ;
        RECT 10.370 25.275 11.455 25.615 ;
        RECT 11.790 25.275 11.960 25.635 ;
        RECT 12.130 25.105 12.460 25.465 ;
        RECT 12.630 25.275 12.800 25.635 ;
        RECT 13.505 25.635 14.580 25.805 ;
        RECT 15.435 25.795 16.025 26.115 ;
        RECT 15.435 25.675 15.605 25.795 ;
        RECT 12.970 25.105 13.300 25.485 ;
        RECT 13.505 25.275 13.740 25.635 ;
        RECT 13.910 25.105 14.240 25.465 ;
        RECT 14.410 25.275 14.580 25.635 ;
        RECT 14.830 25.275 15.605 25.675 ;
        RECT 15.775 25.105 16.025 25.590 ;
        RECT 16.195 25.275 16.455 26.255 ;
        RECT 8.730 24.935 16.540 25.105 ;
        RECT 19.485 25.065 19.775 26.230 ;
        RECT 19.970 26.215 20.300 26.890 ;
        RECT 20.545 26.705 20.715 26.915 ;
        RECT 20.470 26.375 20.715 26.705 ;
        RECT 21.750 26.745 22.245 26.935 ;
        RECT 22.460 26.915 23.470 27.085 ;
        RECT 24.240 27.085 24.410 27.445 ;
        RECT 24.580 27.255 24.910 27.615 ;
        RECT 25.080 27.085 25.250 27.445 ;
        RECT 24.240 26.915 25.250 27.085 ;
        RECT 25.500 27.065 26.100 27.445 ;
        RECT 26.365 27.235 26.695 27.615 ;
        RECT 25.500 26.895 26.695 27.065 ;
        RECT 25.500 26.765 25.740 26.895 ;
        RECT 20.885 26.425 21.325 26.665 ;
        RECT 21.750 26.575 22.415 26.745 ;
        RECT 22.585 26.425 22.960 26.745 ;
        RECT 23.255 26.450 24.420 26.735 ;
        RECT 26.525 26.705 26.695 26.895 ;
        RECT 26.865 26.870 27.125 27.445 ;
        RECT 29.235 26.890 29.525 27.615 ;
        RECT 29.730 26.890 30.130 27.445 ;
        RECT 30.375 27.255 30.705 27.615 ;
        RECT 30.875 27.195 31.885 27.445 ;
        RECT 30.875 27.085 31.045 27.195 ;
        RECT 31.715 27.105 31.885 27.195 ;
        RECT 30.305 26.915 31.045 27.085 ;
        RECT 32.220 27.085 32.390 27.445 ;
        RECT 32.560 27.255 32.890 27.615 ;
        RECT 33.060 27.085 33.230 27.445 ;
        RECT 33.400 27.210 33.730 27.615 ;
        RECT 19.970 25.235 20.370 26.215 ;
        RECT 20.545 25.765 20.715 26.375 ;
        RECT 21.155 25.935 21.575 26.255 ;
        RECT 23.255 26.185 23.425 26.450 ;
        RECT 21.805 26.015 23.425 26.185 ;
        RECT 20.545 25.595 21.210 25.765 ;
        RECT 21.805 25.745 22.055 26.015 ;
        RECT 23.650 25.935 24.010 26.265 ;
        RECT 24.250 26.105 24.420 26.450 ;
        RECT 24.590 26.340 24.980 26.670 ;
        RECT 25.170 26.425 25.540 26.595 ;
        RECT 25.970 26.425 26.300 26.705 ;
        RECT 25.170 26.105 25.340 26.425 ;
        RECT 26.130 26.375 26.300 26.425 ;
        RECT 26.525 26.375 26.780 26.705 ;
        RECT 24.250 25.935 25.340 26.105 ;
        RECT 25.510 25.820 25.910 26.255 ;
        RECT 26.525 26.075 26.695 26.375 ;
        RECT 26.950 26.215 27.125 26.870 ;
        RECT 21.040 25.575 21.210 25.595 ;
        RECT 22.460 25.595 23.470 25.765 ;
        RECT 20.540 25.065 20.870 25.425 ;
        RECT 21.040 25.235 22.125 25.575 ;
        RECT 22.460 25.235 22.630 25.595 ;
        RECT 22.800 25.065 23.130 25.425 ;
        RECT 23.300 25.235 23.470 25.595 ;
        RECT 24.175 25.595 25.250 25.765 ;
        RECT 26.105 25.755 26.695 26.075 ;
        RECT 26.105 25.635 26.275 25.755 ;
        RECT 23.640 25.065 23.970 25.445 ;
        RECT 24.175 25.235 24.410 25.595 ;
        RECT 24.580 25.065 24.910 25.425 ;
        RECT 25.080 25.235 25.250 25.595 ;
        RECT 25.500 25.235 26.275 25.635 ;
        RECT 26.445 25.065 26.695 25.550 ;
        RECT 26.865 25.235 27.125 26.215 ;
        RECT 29.235 25.065 29.525 26.230 ;
        RECT 29.730 26.215 30.060 26.890 ;
        RECT 30.305 26.705 30.475 26.915 ;
        RECT 30.230 26.375 30.475 26.705 ;
        RECT 31.510 26.745 32.005 26.935 ;
        RECT 32.220 26.915 33.230 27.085 ;
        RECT 34.000 27.085 34.170 27.445 ;
        RECT 34.340 27.255 34.670 27.615 ;
        RECT 34.840 27.085 35.010 27.445 ;
        RECT 34.000 26.915 35.010 27.085 ;
        RECT 35.260 27.065 35.860 27.445 ;
        RECT 36.125 27.235 36.455 27.615 ;
        RECT 35.260 26.895 36.455 27.065 ;
        RECT 35.260 26.765 35.500 26.895 ;
        RECT 30.645 26.425 31.085 26.665 ;
        RECT 31.510 26.575 32.175 26.745 ;
        RECT 32.345 26.425 32.720 26.745 ;
        RECT 33.015 26.450 34.180 26.735 ;
        RECT 36.285 26.705 36.455 26.895 ;
        RECT 36.625 26.870 36.885 27.445 ;
        RECT 39.245 26.920 39.535 27.645 ;
        RECT 39.740 26.920 40.140 27.475 ;
        RECT 40.385 27.285 40.715 27.645 ;
        RECT 40.885 27.225 41.895 27.475 ;
        RECT 40.885 27.115 41.055 27.225 ;
        RECT 41.725 27.135 41.895 27.225 ;
        RECT 40.315 26.945 41.055 27.115 ;
        RECT 42.230 27.115 42.400 27.475 ;
        RECT 42.570 27.285 42.900 27.645 ;
        RECT 43.070 27.115 43.240 27.475 ;
        RECT 43.410 27.240 43.740 27.645 ;
        RECT 29.730 25.235 30.130 26.215 ;
        RECT 30.305 25.765 30.475 26.375 ;
        RECT 30.915 25.935 31.335 26.255 ;
        RECT 33.015 26.185 33.185 26.450 ;
        RECT 31.565 26.015 33.185 26.185 ;
        RECT 30.305 25.595 30.970 25.765 ;
        RECT 31.565 25.745 31.815 26.015 ;
        RECT 33.410 25.935 33.770 26.265 ;
        RECT 34.010 26.105 34.180 26.450 ;
        RECT 34.350 26.340 34.740 26.670 ;
        RECT 34.930 26.425 35.300 26.595 ;
        RECT 35.730 26.425 36.060 26.705 ;
        RECT 34.930 26.105 35.100 26.425 ;
        RECT 35.890 26.375 36.060 26.425 ;
        RECT 36.285 26.375 36.540 26.705 ;
        RECT 34.010 25.935 35.100 26.105 ;
        RECT 35.270 25.820 35.670 26.255 ;
        RECT 36.285 26.075 36.455 26.375 ;
        RECT 36.710 26.215 36.885 26.870 ;
        RECT 30.800 25.575 30.970 25.595 ;
        RECT 32.220 25.595 33.230 25.765 ;
        RECT 30.300 25.065 30.630 25.425 ;
        RECT 30.800 25.235 31.885 25.575 ;
        RECT 32.220 25.235 32.390 25.595 ;
        RECT 32.560 25.065 32.890 25.425 ;
        RECT 33.060 25.235 33.230 25.595 ;
        RECT 33.935 25.595 35.010 25.765 ;
        RECT 35.865 25.755 36.455 26.075 ;
        RECT 35.865 25.635 36.035 25.755 ;
        RECT 33.400 25.065 33.730 25.445 ;
        RECT 33.935 25.235 34.170 25.595 ;
        RECT 34.340 25.065 34.670 25.425 ;
        RECT 34.840 25.235 35.010 25.595 ;
        RECT 35.260 25.235 36.035 25.635 ;
        RECT 36.205 25.065 36.455 25.550 ;
        RECT 36.625 25.235 36.885 26.215 ;
        RECT 39.245 25.095 39.535 26.260 ;
        RECT 39.740 26.245 40.070 26.920 ;
        RECT 40.315 26.735 40.485 26.945 ;
        RECT 40.240 26.405 40.485 26.735 ;
        RECT 41.520 26.775 42.015 26.965 ;
        RECT 42.230 26.945 43.240 27.115 ;
        RECT 44.010 27.115 44.180 27.475 ;
        RECT 44.350 27.285 44.680 27.645 ;
        RECT 44.850 27.115 45.020 27.475 ;
        RECT 44.010 26.945 45.020 27.115 ;
        RECT 45.270 27.095 45.870 27.475 ;
        RECT 46.135 27.265 46.465 27.645 ;
        RECT 45.270 26.925 46.465 27.095 ;
        RECT 45.270 26.795 45.510 26.925 ;
        RECT 40.655 26.455 41.095 26.695 ;
        RECT 41.520 26.605 42.185 26.775 ;
        RECT 42.355 26.455 42.730 26.775 ;
        RECT 43.025 26.480 44.190 26.765 ;
        RECT 46.295 26.735 46.465 26.925 ;
        RECT 46.635 26.900 46.895 27.475 ;
        RECT 49.725 27.205 50.015 28.370 ;
        RECT 50.210 28.355 50.540 29.030 ;
        RECT 50.785 28.845 50.955 29.055 ;
        RECT 50.710 28.515 50.955 28.845 ;
        RECT 51.990 28.885 52.485 29.075 ;
        RECT 52.700 29.055 53.710 29.225 ;
        RECT 54.480 29.225 54.650 29.585 ;
        RECT 54.820 29.395 55.150 29.755 ;
        RECT 55.320 29.225 55.490 29.585 ;
        RECT 54.480 29.055 55.490 29.225 ;
        RECT 55.740 29.205 56.340 29.585 ;
        RECT 56.605 29.375 56.935 29.755 ;
        RECT 59.940 29.695 67.760 29.865 ;
        RECT 69.730 29.735 77.550 29.905 ;
        RECT 79.710 29.765 87.520 29.935 ;
        RECT 55.740 29.035 56.935 29.205 ;
        RECT 55.740 28.905 55.980 29.035 ;
        RECT 51.125 28.565 51.565 28.805 ;
        RECT 51.990 28.715 52.655 28.885 ;
        RECT 52.825 28.565 53.200 28.885 ;
        RECT 53.495 28.590 54.660 28.875 ;
        RECT 56.765 28.845 56.935 29.035 ;
        RECT 57.105 29.010 57.365 29.585 ;
        RECT 50.210 27.375 50.610 28.355 ;
        RECT 50.785 27.905 50.955 28.515 ;
        RECT 51.395 28.075 51.815 28.395 ;
        RECT 53.495 28.325 53.665 28.590 ;
        RECT 52.045 28.155 53.665 28.325 ;
        RECT 50.785 27.735 51.450 27.905 ;
        RECT 52.045 27.885 52.295 28.155 ;
        RECT 53.890 28.075 54.250 28.405 ;
        RECT 54.490 28.245 54.660 28.590 ;
        RECT 54.830 28.480 55.220 28.810 ;
        RECT 55.410 28.565 55.780 28.735 ;
        RECT 56.210 28.565 56.540 28.845 ;
        RECT 55.410 28.245 55.580 28.565 ;
        RECT 56.370 28.515 56.540 28.565 ;
        RECT 56.765 28.515 57.020 28.845 ;
        RECT 54.490 28.075 55.580 28.245 ;
        RECT 55.750 27.960 56.150 28.395 ;
        RECT 56.765 28.215 56.935 28.515 ;
        RECT 57.190 28.355 57.365 29.010 ;
        RECT 60.025 28.970 60.315 29.695 ;
        RECT 60.520 28.970 60.920 29.525 ;
        RECT 61.165 29.335 61.495 29.695 ;
        RECT 61.665 29.275 62.675 29.525 ;
        RECT 61.665 29.165 61.835 29.275 ;
        RECT 62.505 29.185 62.675 29.275 ;
        RECT 61.095 28.995 61.835 29.165 ;
        RECT 63.010 29.165 63.180 29.525 ;
        RECT 63.350 29.335 63.680 29.695 ;
        RECT 63.850 29.165 64.020 29.525 ;
        RECT 64.190 29.290 64.520 29.695 ;
        RECT 51.280 27.715 51.450 27.735 ;
        RECT 52.700 27.735 53.710 27.905 ;
        RECT 50.780 27.205 51.110 27.565 ;
        RECT 51.280 27.375 52.365 27.715 ;
        RECT 52.700 27.375 52.870 27.735 ;
        RECT 53.040 27.205 53.370 27.565 ;
        RECT 53.540 27.375 53.710 27.735 ;
        RECT 54.415 27.735 55.490 27.905 ;
        RECT 56.345 27.895 56.935 28.215 ;
        RECT 56.345 27.775 56.515 27.895 ;
        RECT 53.880 27.205 54.210 27.585 ;
        RECT 54.415 27.375 54.650 27.735 ;
        RECT 54.820 27.205 55.150 27.565 ;
        RECT 55.320 27.375 55.490 27.735 ;
        RECT 55.740 27.375 56.515 27.775 ;
        RECT 56.685 27.205 56.935 27.690 ;
        RECT 57.105 27.375 57.365 28.355 ;
        RECT 49.640 27.035 57.450 27.205 ;
        RECT 60.025 27.145 60.315 28.310 ;
        RECT 60.520 28.295 60.850 28.970 ;
        RECT 61.095 28.785 61.265 28.995 ;
        RECT 61.020 28.455 61.265 28.785 ;
        RECT 62.300 28.825 62.795 29.015 ;
        RECT 63.010 28.995 64.020 29.165 ;
        RECT 64.790 29.165 64.960 29.525 ;
        RECT 65.130 29.335 65.460 29.695 ;
        RECT 65.630 29.165 65.800 29.525 ;
        RECT 64.790 28.995 65.800 29.165 ;
        RECT 66.050 29.145 66.650 29.525 ;
        RECT 66.915 29.315 67.245 29.695 ;
        RECT 66.050 28.975 67.245 29.145 ;
        RECT 66.050 28.845 66.290 28.975 ;
        RECT 61.435 28.505 61.875 28.745 ;
        RECT 62.300 28.655 62.965 28.825 ;
        RECT 63.135 28.505 63.510 28.825 ;
        RECT 63.805 28.530 64.970 28.815 ;
        RECT 67.075 28.785 67.245 28.975 ;
        RECT 67.415 28.950 67.675 29.525 ;
        RECT 69.815 29.010 70.105 29.735 ;
        RECT 70.310 29.010 70.710 29.565 ;
        RECT 70.955 29.375 71.285 29.735 ;
        RECT 71.455 29.315 72.465 29.565 ;
        RECT 71.455 29.205 71.625 29.315 ;
        RECT 72.295 29.225 72.465 29.315 ;
        RECT 70.885 29.035 71.625 29.205 ;
        RECT 72.800 29.205 72.970 29.565 ;
        RECT 73.140 29.375 73.470 29.735 ;
        RECT 73.640 29.205 73.810 29.565 ;
        RECT 73.980 29.330 74.310 29.735 ;
        RECT 60.520 27.315 60.920 28.295 ;
        RECT 61.095 27.845 61.265 28.455 ;
        RECT 61.705 28.015 62.125 28.335 ;
        RECT 63.805 28.265 63.975 28.530 ;
        RECT 62.355 28.095 63.975 28.265 ;
        RECT 61.095 27.675 61.760 27.845 ;
        RECT 62.355 27.825 62.605 28.095 ;
        RECT 64.200 28.015 64.560 28.345 ;
        RECT 64.800 28.185 64.970 28.530 ;
        RECT 65.140 28.420 65.530 28.750 ;
        RECT 65.720 28.505 66.090 28.675 ;
        RECT 66.520 28.505 66.850 28.785 ;
        RECT 65.720 28.185 65.890 28.505 ;
        RECT 66.680 28.455 66.850 28.505 ;
        RECT 67.075 28.455 67.330 28.785 ;
        RECT 64.800 28.015 65.890 28.185 ;
        RECT 66.060 27.900 66.460 28.335 ;
        RECT 67.075 28.155 67.245 28.455 ;
        RECT 67.500 28.295 67.675 28.950 ;
        RECT 61.590 27.655 61.760 27.675 ;
        RECT 63.010 27.675 64.020 27.845 ;
        RECT 61.090 27.145 61.420 27.505 ;
        RECT 61.590 27.315 62.675 27.655 ;
        RECT 63.010 27.315 63.180 27.675 ;
        RECT 63.350 27.145 63.680 27.505 ;
        RECT 63.850 27.315 64.020 27.675 ;
        RECT 64.725 27.675 65.800 27.845 ;
        RECT 66.655 27.835 67.245 28.155 ;
        RECT 66.655 27.715 66.825 27.835 ;
        RECT 64.190 27.145 64.520 27.525 ;
        RECT 64.725 27.315 64.960 27.675 ;
        RECT 65.130 27.145 65.460 27.505 ;
        RECT 65.630 27.315 65.800 27.675 ;
        RECT 66.050 27.315 66.825 27.715 ;
        RECT 66.995 27.145 67.245 27.630 ;
        RECT 67.415 27.315 67.675 28.295 ;
        RECT 69.815 27.185 70.105 28.350 ;
        RECT 70.310 28.335 70.640 29.010 ;
        RECT 70.885 28.825 71.055 29.035 ;
        RECT 70.810 28.495 71.055 28.825 ;
        RECT 72.090 28.865 72.585 29.055 ;
        RECT 72.800 29.035 73.810 29.205 ;
        RECT 74.580 29.205 74.750 29.565 ;
        RECT 74.920 29.375 75.250 29.735 ;
        RECT 75.420 29.205 75.590 29.565 ;
        RECT 74.580 29.035 75.590 29.205 ;
        RECT 75.840 29.185 76.440 29.565 ;
        RECT 76.705 29.355 77.035 29.735 ;
        RECT 75.840 29.015 77.035 29.185 ;
        RECT 75.840 28.885 76.080 29.015 ;
        RECT 71.225 28.545 71.665 28.785 ;
        RECT 72.090 28.695 72.755 28.865 ;
        RECT 72.925 28.545 73.300 28.865 ;
        RECT 73.595 28.570 74.760 28.855 ;
        RECT 76.865 28.825 77.035 29.015 ;
        RECT 77.205 28.990 77.465 29.565 ;
        RECT 79.795 29.040 80.085 29.765 ;
        RECT 80.280 29.040 80.680 29.595 ;
        RECT 80.925 29.405 81.255 29.765 ;
        RECT 81.425 29.345 82.435 29.595 ;
        RECT 81.425 29.235 81.595 29.345 ;
        RECT 82.265 29.255 82.435 29.345 ;
        RECT 80.855 29.065 81.595 29.235 ;
        RECT 82.770 29.235 82.940 29.595 ;
        RECT 83.110 29.405 83.440 29.765 ;
        RECT 83.610 29.235 83.780 29.595 ;
        RECT 83.950 29.360 84.280 29.765 ;
        RECT 70.310 27.355 70.710 28.335 ;
        RECT 70.885 27.885 71.055 28.495 ;
        RECT 71.495 28.055 71.915 28.375 ;
        RECT 73.595 28.305 73.765 28.570 ;
        RECT 72.145 28.135 73.765 28.305 ;
        RECT 70.885 27.715 71.550 27.885 ;
        RECT 72.145 27.865 72.395 28.135 ;
        RECT 73.990 28.055 74.350 28.385 ;
        RECT 74.590 28.225 74.760 28.570 ;
        RECT 74.930 28.460 75.320 28.790 ;
        RECT 75.510 28.545 75.880 28.715 ;
        RECT 76.310 28.545 76.640 28.825 ;
        RECT 75.510 28.225 75.680 28.545 ;
        RECT 76.470 28.495 76.640 28.545 ;
        RECT 76.865 28.495 77.120 28.825 ;
        RECT 74.590 28.055 75.680 28.225 ;
        RECT 75.850 27.940 76.250 28.375 ;
        RECT 76.865 28.195 77.035 28.495 ;
        RECT 77.290 28.335 77.465 28.990 ;
        RECT 71.380 27.695 71.550 27.715 ;
        RECT 72.800 27.715 73.810 27.885 ;
        RECT 70.880 27.185 71.210 27.545 ;
        RECT 71.380 27.355 72.465 27.695 ;
        RECT 72.800 27.355 72.970 27.715 ;
        RECT 73.140 27.185 73.470 27.545 ;
        RECT 73.640 27.355 73.810 27.715 ;
        RECT 74.515 27.715 75.590 27.885 ;
        RECT 76.445 27.875 77.035 28.195 ;
        RECT 76.445 27.755 76.615 27.875 ;
        RECT 73.980 27.185 74.310 27.565 ;
        RECT 74.515 27.355 74.750 27.715 ;
        RECT 74.920 27.185 75.250 27.545 ;
        RECT 75.420 27.355 75.590 27.715 ;
        RECT 75.840 27.355 76.615 27.755 ;
        RECT 76.785 27.185 77.035 27.670 ;
        RECT 77.205 27.355 77.465 28.335 ;
        RECT 79.795 27.215 80.085 28.380 ;
        RECT 80.280 28.365 80.610 29.040 ;
        RECT 80.855 28.855 81.025 29.065 ;
        RECT 80.780 28.525 81.025 28.855 ;
        RECT 82.060 28.895 82.555 29.085 ;
        RECT 82.770 29.065 83.780 29.235 ;
        RECT 84.550 29.235 84.720 29.595 ;
        RECT 84.890 29.405 85.220 29.765 ;
        RECT 85.390 29.235 85.560 29.595 ;
        RECT 84.550 29.065 85.560 29.235 ;
        RECT 85.810 29.215 86.410 29.595 ;
        RECT 86.675 29.385 87.005 29.765 ;
        RECT 85.810 29.045 87.005 29.215 ;
        RECT 85.810 28.915 86.050 29.045 ;
        RECT 81.195 28.575 81.635 28.815 ;
        RECT 82.060 28.725 82.725 28.895 ;
        RECT 82.895 28.575 83.270 28.895 ;
        RECT 83.565 28.600 84.730 28.885 ;
        RECT 86.835 28.855 87.005 29.045 ;
        RECT 87.175 29.020 87.435 29.595 ;
        RECT 80.280 27.385 80.680 28.365 ;
        RECT 80.855 27.915 81.025 28.525 ;
        RECT 81.465 28.085 81.885 28.405 ;
        RECT 83.565 28.335 83.735 28.600 ;
        RECT 82.115 28.165 83.735 28.335 ;
        RECT 80.855 27.745 81.520 27.915 ;
        RECT 82.115 27.895 82.365 28.165 ;
        RECT 83.960 28.085 84.320 28.415 ;
        RECT 84.560 28.255 84.730 28.600 ;
        RECT 84.900 28.490 85.290 28.820 ;
        RECT 85.480 28.575 85.850 28.745 ;
        RECT 86.280 28.575 86.610 28.855 ;
        RECT 85.480 28.255 85.650 28.575 ;
        RECT 86.440 28.525 86.610 28.575 ;
        RECT 86.835 28.525 87.090 28.855 ;
        RECT 84.560 28.085 85.650 28.255 ;
        RECT 85.820 27.970 86.220 28.405 ;
        RECT 86.835 28.225 87.005 28.525 ;
        RECT 87.260 28.365 87.435 29.020 ;
        RECT 81.350 27.725 81.520 27.745 ;
        RECT 82.770 27.745 83.780 27.915 ;
        RECT 80.850 27.215 81.180 27.575 ;
        RECT 81.350 27.385 82.435 27.725 ;
        RECT 82.770 27.385 82.940 27.745 ;
        RECT 83.110 27.215 83.440 27.575 ;
        RECT 83.610 27.385 83.780 27.745 ;
        RECT 84.485 27.745 85.560 27.915 ;
        RECT 86.415 27.905 87.005 28.225 ;
        RECT 86.415 27.785 86.585 27.905 ;
        RECT 83.950 27.215 84.280 27.595 ;
        RECT 84.485 27.385 84.720 27.745 ;
        RECT 84.890 27.215 85.220 27.575 ;
        RECT 85.390 27.385 85.560 27.745 ;
        RECT 85.810 27.385 86.585 27.785 ;
        RECT 86.755 27.215 87.005 27.700 ;
        RECT 87.175 27.385 87.435 28.365 ;
        RECT 59.940 26.975 67.760 27.145 ;
        RECT 69.730 27.015 77.550 27.185 ;
        RECT 79.710 27.045 87.520 27.215 ;
        RECT 39.740 25.265 40.140 26.245 ;
        RECT 40.315 25.795 40.485 26.405 ;
        RECT 40.925 25.965 41.345 26.285 ;
        RECT 43.025 26.215 43.195 26.480 ;
        RECT 41.575 26.045 43.195 26.215 ;
        RECT 40.315 25.625 40.980 25.795 ;
        RECT 41.575 25.775 41.825 26.045 ;
        RECT 43.420 25.965 43.780 26.295 ;
        RECT 44.020 26.135 44.190 26.480 ;
        RECT 44.360 26.370 44.750 26.700 ;
        RECT 44.940 26.455 45.310 26.625 ;
        RECT 45.740 26.455 46.070 26.735 ;
        RECT 44.940 26.135 45.110 26.455 ;
        RECT 45.900 26.405 46.070 26.455 ;
        RECT 46.295 26.405 46.550 26.735 ;
        RECT 44.020 25.965 45.110 26.135 ;
        RECT 45.280 25.850 45.680 26.285 ;
        RECT 46.295 26.105 46.465 26.405 ;
        RECT 46.720 26.245 46.895 26.900 ;
        RECT 91.510 26.895 96.110 27.065 ;
        RECT 40.810 25.605 40.980 25.625 ;
        RECT 42.230 25.625 43.240 25.795 ;
        RECT 40.310 25.095 40.640 25.455 ;
        RECT 40.810 25.265 41.895 25.605 ;
        RECT 42.230 25.265 42.400 25.625 ;
        RECT 42.570 25.095 42.900 25.455 ;
        RECT 43.070 25.265 43.240 25.625 ;
        RECT 43.945 25.625 45.020 25.795 ;
        RECT 45.875 25.785 46.465 26.105 ;
        RECT 45.875 25.665 46.045 25.785 ;
        RECT 43.410 25.095 43.740 25.475 ;
        RECT 43.945 25.265 44.180 25.625 ;
        RECT 44.350 25.095 44.680 25.455 ;
        RECT 44.850 25.265 45.020 25.625 ;
        RECT 45.270 25.265 46.045 25.665 ;
        RECT 46.215 25.095 46.465 25.580 ;
        RECT 46.635 25.265 46.895 26.245 ;
        RECT 91.870 26.085 92.115 26.690 ;
        RECT 92.335 26.360 92.845 26.895 ;
        RECT 91.595 25.915 92.825 26.085 ;
        RECT 50.230 25.385 58.050 25.555 ;
        RECT 19.400 24.895 27.210 25.065 ;
        RECT 29.150 24.895 36.970 25.065 ;
        RECT 39.160 24.925 46.980 25.095 ;
        RECT 50.350 24.660 50.750 25.215 ;
        RECT 50.995 25.025 51.325 25.385 ;
        RECT 51.495 24.965 52.505 25.215 ;
        RECT 51.495 24.855 51.665 24.965 ;
        RECT 52.335 24.875 52.505 24.965 ;
        RECT 50.925 24.685 51.665 24.855 ;
        RECT 52.840 24.855 53.010 25.215 ;
        RECT 53.180 25.025 53.510 25.385 ;
        RECT 53.680 24.855 53.850 25.215 ;
        RECT 54.020 24.980 54.350 25.385 ;
        RECT 50.350 23.985 50.680 24.660 ;
        RECT 50.925 24.475 51.095 24.685 ;
        RECT 50.850 24.145 51.095 24.475 ;
        RECT 52.130 24.515 52.625 24.705 ;
        RECT 52.840 24.685 53.850 24.855 ;
        RECT 54.620 24.855 54.790 25.215 ;
        RECT 54.960 25.025 55.290 25.385 ;
        RECT 55.460 24.855 55.630 25.215 ;
        RECT 54.620 24.685 55.630 24.855 ;
        RECT 55.880 24.835 56.480 25.215 ;
        RECT 56.745 25.005 57.075 25.385 ;
        RECT 55.880 24.665 57.075 24.835 ;
        RECT 55.880 24.535 56.120 24.665 ;
        RECT 51.265 24.195 51.705 24.435 ;
        RECT 52.130 24.345 52.795 24.515 ;
        RECT 52.965 24.195 53.340 24.515 ;
        RECT 53.635 24.220 54.800 24.505 ;
        RECT 56.905 24.475 57.075 24.665 ;
        RECT 57.245 24.640 57.505 25.215 ;
        RECT 57.675 24.660 57.965 25.385 ;
        RECT 61.140 25.165 68.940 25.335 ;
        RECT 50.350 23.005 50.750 23.985 ;
        RECT 50.925 23.535 51.095 24.145 ;
        RECT 51.535 23.705 51.955 24.025 ;
        RECT 53.635 23.955 53.805 24.220 ;
        RECT 52.185 23.785 53.805 23.955 ;
        RECT 50.925 23.365 51.590 23.535 ;
        RECT 52.185 23.515 52.435 23.785 ;
        RECT 54.030 23.705 54.390 24.035 ;
        RECT 54.630 23.875 54.800 24.220 ;
        RECT 54.970 24.110 55.360 24.440 ;
        RECT 55.550 24.195 55.920 24.365 ;
        RECT 56.350 24.195 56.680 24.475 ;
        RECT 55.550 23.875 55.720 24.195 ;
        RECT 56.510 24.145 56.680 24.195 ;
        RECT 56.905 24.145 57.160 24.475 ;
        RECT 54.630 23.705 55.720 23.875 ;
        RECT 55.890 23.590 56.290 24.025 ;
        RECT 56.905 23.845 57.075 24.145 ;
        RECT 57.330 23.985 57.505 24.640 ;
        RECT 61.225 24.440 61.515 25.165 ;
        RECT 61.700 24.440 62.100 24.995 ;
        RECT 62.345 24.805 62.675 25.165 ;
        RECT 62.845 24.745 63.855 24.995 ;
        RECT 62.845 24.635 63.015 24.745 ;
        RECT 63.685 24.655 63.855 24.745 ;
        RECT 62.275 24.465 63.015 24.635 ;
        RECT 64.190 24.635 64.360 24.995 ;
        RECT 64.530 24.805 64.860 25.165 ;
        RECT 65.030 24.635 65.200 24.995 ;
        RECT 65.370 24.760 65.700 25.165 ;
        RECT 51.420 23.345 51.590 23.365 ;
        RECT 52.840 23.365 53.850 23.535 ;
        RECT 50.920 22.835 51.250 23.195 ;
        RECT 51.420 23.005 52.505 23.345 ;
        RECT 52.840 23.005 53.010 23.365 ;
        RECT 53.180 22.835 53.510 23.195 ;
        RECT 53.680 23.005 53.850 23.365 ;
        RECT 54.555 23.365 55.630 23.535 ;
        RECT 56.485 23.525 57.075 23.845 ;
        RECT 56.485 23.405 56.655 23.525 ;
        RECT 54.020 22.835 54.350 23.215 ;
        RECT 54.555 23.005 54.790 23.365 ;
        RECT 54.960 22.835 55.290 23.195 ;
        RECT 55.460 23.005 55.630 23.365 ;
        RECT 55.880 23.005 56.655 23.405 ;
        RECT 56.825 22.835 57.075 23.320 ;
        RECT 57.245 23.005 57.505 23.985 ;
        RECT 57.675 22.835 57.965 24.000 ;
        RECT 50.230 22.665 58.050 22.835 ;
        RECT 61.225 22.615 61.515 23.780 ;
        RECT 61.700 23.765 62.030 24.440 ;
        RECT 62.275 24.255 62.445 24.465 ;
        RECT 62.200 23.925 62.445 24.255 ;
        RECT 63.480 24.295 63.975 24.485 ;
        RECT 64.190 24.465 65.200 24.635 ;
        RECT 65.970 24.635 66.140 24.995 ;
        RECT 66.310 24.805 66.640 25.165 ;
        RECT 66.810 24.635 66.980 24.995 ;
        RECT 65.970 24.465 66.980 24.635 ;
        RECT 67.230 24.615 67.830 24.995 ;
        RECT 68.095 24.785 68.425 25.165 ;
        RECT 71.140 25.135 78.950 25.305 ;
        RECT 67.230 24.445 68.425 24.615 ;
        RECT 67.230 24.315 67.470 24.445 ;
        RECT 62.615 23.975 63.055 24.215 ;
        RECT 63.480 24.125 64.145 24.295 ;
        RECT 64.315 23.975 64.690 24.295 ;
        RECT 64.985 24.000 66.150 24.285 ;
        RECT 68.255 24.255 68.425 24.445 ;
        RECT 68.595 24.420 68.855 24.995 ;
        RECT 61.700 22.785 62.100 23.765 ;
        RECT 62.275 23.315 62.445 23.925 ;
        RECT 62.885 23.485 63.305 23.805 ;
        RECT 64.985 23.735 65.155 24.000 ;
        RECT 63.535 23.565 65.155 23.735 ;
        RECT 62.275 23.145 62.940 23.315 ;
        RECT 63.535 23.295 63.785 23.565 ;
        RECT 65.380 23.485 65.740 23.815 ;
        RECT 65.980 23.655 66.150 24.000 ;
        RECT 66.320 23.890 66.710 24.220 ;
        RECT 66.900 23.975 67.270 24.145 ;
        RECT 67.700 23.975 68.030 24.255 ;
        RECT 66.900 23.655 67.070 23.975 ;
        RECT 67.860 23.925 68.030 23.975 ;
        RECT 68.255 23.925 68.510 24.255 ;
        RECT 65.980 23.485 67.070 23.655 ;
        RECT 67.240 23.370 67.640 23.805 ;
        RECT 68.255 23.625 68.425 23.925 ;
        RECT 68.680 23.765 68.855 24.420 ;
        RECT 71.225 24.410 71.515 25.135 ;
        RECT 71.710 24.410 72.110 24.965 ;
        RECT 72.355 24.775 72.685 25.135 ;
        RECT 72.855 24.715 73.865 24.965 ;
        RECT 72.855 24.605 73.025 24.715 ;
        RECT 73.695 24.625 73.865 24.715 ;
        RECT 72.285 24.435 73.025 24.605 ;
        RECT 74.200 24.605 74.370 24.965 ;
        RECT 74.540 24.775 74.870 25.135 ;
        RECT 75.040 24.605 75.210 24.965 ;
        RECT 75.380 24.730 75.710 25.135 ;
        RECT 62.770 23.125 62.940 23.145 ;
        RECT 64.190 23.145 65.200 23.315 ;
        RECT 62.270 22.615 62.600 22.975 ;
        RECT 62.770 22.785 63.855 23.125 ;
        RECT 64.190 22.785 64.360 23.145 ;
        RECT 64.530 22.615 64.860 22.975 ;
        RECT 65.030 22.785 65.200 23.145 ;
        RECT 65.905 23.145 66.980 23.315 ;
        RECT 67.835 23.305 68.425 23.625 ;
        RECT 67.835 23.185 68.005 23.305 ;
        RECT 65.370 22.615 65.700 22.995 ;
        RECT 65.905 22.785 66.140 23.145 ;
        RECT 66.310 22.615 66.640 22.975 ;
        RECT 66.810 22.785 66.980 23.145 ;
        RECT 67.230 22.785 68.005 23.185 ;
        RECT 68.175 22.615 68.425 23.100 ;
        RECT 68.595 22.785 68.855 23.765 ;
        RECT 61.140 22.445 68.940 22.615 ;
        RECT 71.225 22.585 71.515 23.750 ;
        RECT 71.710 23.735 72.040 24.410 ;
        RECT 72.285 24.225 72.455 24.435 ;
        RECT 72.210 23.895 72.455 24.225 ;
        RECT 73.490 24.265 73.985 24.455 ;
        RECT 74.200 24.435 75.210 24.605 ;
        RECT 75.980 24.605 76.150 24.965 ;
        RECT 76.320 24.775 76.650 25.135 ;
        RECT 76.820 24.605 76.990 24.965 ;
        RECT 75.980 24.435 76.990 24.605 ;
        RECT 77.240 24.585 77.840 24.965 ;
        RECT 78.105 24.755 78.435 25.135 ;
        RECT 81.260 25.045 89.060 25.215 ;
        RECT 91.595 25.105 91.935 25.915 ;
        RECT 92.105 25.350 92.855 25.540 ;
        RECT 77.240 24.415 78.435 24.585 ;
        RECT 77.240 24.285 77.480 24.415 ;
        RECT 72.625 23.945 73.065 24.185 ;
        RECT 73.490 24.095 74.155 24.265 ;
        RECT 74.325 23.945 74.700 24.265 ;
        RECT 74.995 23.970 76.160 24.255 ;
        RECT 78.265 24.225 78.435 24.415 ;
        RECT 78.605 24.390 78.865 24.965 ;
        RECT 71.710 22.755 72.110 23.735 ;
        RECT 72.285 23.285 72.455 23.895 ;
        RECT 72.895 23.455 73.315 23.775 ;
        RECT 74.995 23.705 75.165 23.970 ;
        RECT 73.545 23.535 75.165 23.705 ;
        RECT 72.285 23.115 72.950 23.285 ;
        RECT 73.545 23.265 73.795 23.535 ;
        RECT 75.390 23.455 75.750 23.785 ;
        RECT 75.990 23.625 76.160 23.970 ;
        RECT 76.330 23.860 76.720 24.190 ;
        RECT 76.910 23.945 77.280 24.115 ;
        RECT 77.710 23.945 78.040 24.225 ;
        RECT 76.910 23.625 77.080 23.945 ;
        RECT 77.870 23.895 78.040 23.945 ;
        RECT 78.265 23.895 78.520 24.225 ;
        RECT 75.990 23.455 77.080 23.625 ;
        RECT 77.250 23.340 77.650 23.775 ;
        RECT 78.265 23.595 78.435 23.895 ;
        RECT 78.690 23.735 78.865 24.390 ;
        RECT 81.345 24.320 81.635 25.045 ;
        RECT 81.820 24.320 82.220 24.875 ;
        RECT 82.465 24.685 82.795 25.045 ;
        RECT 82.965 24.625 83.975 24.875 ;
        RECT 82.965 24.515 83.135 24.625 ;
        RECT 83.805 24.535 83.975 24.625 ;
        RECT 82.395 24.345 83.135 24.515 ;
        RECT 84.310 24.515 84.480 24.875 ;
        RECT 84.650 24.685 84.980 25.045 ;
        RECT 85.150 24.515 85.320 24.875 ;
        RECT 85.490 24.640 85.820 25.045 ;
        RECT 72.780 23.095 72.950 23.115 ;
        RECT 74.200 23.115 75.210 23.285 ;
        RECT 72.280 22.585 72.610 22.945 ;
        RECT 72.780 22.755 73.865 23.095 ;
        RECT 74.200 22.755 74.370 23.115 ;
        RECT 74.540 22.585 74.870 22.945 ;
        RECT 75.040 22.755 75.210 23.115 ;
        RECT 75.915 23.115 76.990 23.285 ;
        RECT 77.845 23.275 78.435 23.595 ;
        RECT 77.845 23.155 78.015 23.275 ;
        RECT 75.380 22.585 75.710 22.965 ;
        RECT 75.915 22.755 76.150 23.115 ;
        RECT 76.320 22.585 76.650 22.945 ;
        RECT 76.820 22.755 76.990 23.115 ;
        RECT 77.240 22.755 78.015 23.155 ;
        RECT 78.185 22.585 78.435 23.070 ;
        RECT 78.605 22.755 78.865 23.735 ;
        RECT 71.140 22.415 78.950 22.585 ;
        RECT 81.345 22.495 81.635 23.660 ;
        RECT 81.820 23.645 82.150 24.320 ;
        RECT 82.395 24.135 82.565 24.345 ;
        RECT 82.320 23.805 82.565 24.135 ;
        RECT 83.600 24.175 84.095 24.365 ;
        RECT 84.310 24.345 85.320 24.515 ;
        RECT 86.090 24.515 86.260 24.875 ;
        RECT 86.430 24.685 86.760 25.045 ;
        RECT 86.930 24.515 87.100 24.875 ;
        RECT 86.090 24.345 87.100 24.515 ;
        RECT 87.350 24.495 87.950 24.875 ;
        RECT 88.215 24.665 88.545 25.045 ;
        RECT 87.350 24.325 88.545 24.495 ;
        RECT 87.350 24.195 87.590 24.325 ;
        RECT 82.735 23.855 83.175 24.095 ;
        RECT 83.600 24.005 84.265 24.175 ;
        RECT 84.435 23.855 84.810 24.175 ;
        RECT 85.105 23.880 86.270 24.165 ;
        RECT 88.375 24.135 88.545 24.325 ;
        RECT 88.715 24.300 88.975 24.875 ;
        RECT 91.595 24.695 92.110 25.105 ;
        RECT 92.345 24.345 92.515 25.105 ;
        RECT 92.685 24.685 92.855 25.350 ;
        RECT 93.025 25.365 93.215 26.725 ;
        RECT 93.385 25.565 93.660 26.725 ;
        RECT 93.850 26.360 94.380 26.725 ;
        RECT 94.805 26.495 95.135 26.895 ;
        RECT 94.205 26.325 94.380 26.360 ;
        RECT 93.865 25.365 94.035 26.165 ;
        RECT 93.025 25.195 94.035 25.365 ;
        RECT 94.205 26.155 95.135 26.325 ;
        RECT 95.305 26.155 95.560 26.725 ;
        RECT 95.735 26.170 96.025 26.895 ;
        RECT 94.205 25.025 94.375 26.155 ;
        RECT 94.965 25.985 95.135 26.155 ;
        RECT 93.250 24.855 94.375 25.025 ;
        RECT 94.545 25.655 94.740 25.985 ;
        RECT 94.965 25.655 95.220 25.985 ;
        RECT 94.545 24.685 94.715 25.655 ;
        RECT 95.390 25.485 95.560 26.155 ;
        RECT 92.685 24.515 94.715 24.685 ;
        RECT 94.885 24.345 95.055 25.485 ;
        RECT 95.225 24.515 95.560 25.485 ;
        RECT 95.735 24.345 96.025 25.510 ;
        RECT 81.820 22.665 82.220 23.645 ;
        RECT 82.395 23.195 82.565 23.805 ;
        RECT 83.005 23.365 83.425 23.685 ;
        RECT 85.105 23.615 85.275 23.880 ;
        RECT 83.655 23.445 85.275 23.615 ;
        RECT 82.395 23.025 83.060 23.195 ;
        RECT 83.655 23.175 83.905 23.445 ;
        RECT 85.500 23.365 85.860 23.695 ;
        RECT 86.100 23.535 86.270 23.880 ;
        RECT 86.440 23.770 86.830 24.100 ;
        RECT 87.020 23.855 87.390 24.025 ;
        RECT 87.820 23.855 88.150 24.135 ;
        RECT 87.020 23.535 87.190 23.855 ;
        RECT 87.980 23.805 88.150 23.855 ;
        RECT 88.375 23.805 88.630 24.135 ;
        RECT 86.100 23.365 87.190 23.535 ;
        RECT 87.360 23.250 87.760 23.685 ;
        RECT 88.375 23.505 88.545 23.805 ;
        RECT 88.800 23.645 88.975 24.300 ;
        RECT 91.510 24.175 96.110 24.345 ;
        RECT 82.890 23.005 83.060 23.025 ;
        RECT 84.310 23.025 85.320 23.195 ;
        RECT 82.390 22.495 82.720 22.855 ;
        RECT 82.890 22.665 83.975 23.005 ;
        RECT 84.310 22.665 84.480 23.025 ;
        RECT 84.650 22.495 84.980 22.855 ;
        RECT 85.150 22.665 85.320 23.025 ;
        RECT 86.025 23.025 87.100 23.195 ;
        RECT 87.955 23.185 88.545 23.505 ;
        RECT 87.955 23.065 88.125 23.185 ;
        RECT 85.490 22.495 85.820 22.875 ;
        RECT 86.025 22.665 86.260 23.025 ;
        RECT 86.430 22.495 86.760 22.855 ;
        RECT 86.930 22.665 87.100 23.025 ;
        RECT 87.350 22.665 88.125 23.065 ;
        RECT 88.295 22.495 88.545 22.980 ;
        RECT 88.715 22.665 88.975 23.645 ;
        RECT 81.260 22.325 89.060 22.495 ;
        RECT 29.970 16.615 31.790 16.785 ;
        RECT 30.055 15.890 30.345 16.615 ;
        RECT 30.740 15.815 31.070 16.445 ;
        RECT 30.055 14.065 30.345 15.230 ;
        RECT 30.740 15.215 30.970 15.815 ;
        RECT 31.240 15.795 31.470 16.615 ;
        RECT 31.140 15.385 31.470 15.625 ;
        RECT 30.740 14.235 31.070 15.215 ;
        RECT 31.240 14.065 31.450 15.205 ;
        RECT 29.970 13.895 31.790 14.065 ;
        RECT 8.580 11.355 16.390 11.525 ;
        RECT 8.665 10.630 8.955 11.355 ;
        RECT 9.150 10.630 9.550 11.185 ;
        RECT 9.795 10.995 10.125 11.355 ;
        RECT 10.295 10.935 11.305 11.185 ;
        RECT 10.295 10.825 10.465 10.935 ;
        RECT 11.135 10.845 11.305 10.935 ;
        RECT 9.725 10.655 10.465 10.825 ;
        RECT 11.640 10.825 11.810 11.185 ;
        RECT 11.980 10.995 12.310 11.355 ;
        RECT 12.480 10.825 12.650 11.185 ;
        RECT 12.820 10.950 13.150 11.355 ;
        RECT 8.665 8.805 8.955 9.970 ;
        RECT 9.150 9.955 9.480 10.630 ;
        RECT 9.725 10.445 9.895 10.655 ;
        RECT 9.650 10.115 9.895 10.445 ;
        RECT 10.930 10.485 11.425 10.675 ;
        RECT 11.640 10.655 12.650 10.825 ;
        RECT 13.420 10.825 13.590 11.185 ;
        RECT 13.760 10.995 14.090 11.355 ;
        RECT 14.260 10.825 14.430 11.185 ;
        RECT 13.420 10.655 14.430 10.825 ;
        RECT 14.680 10.805 15.280 11.185 ;
        RECT 15.545 10.975 15.875 11.355 ;
        RECT 18.930 11.335 26.740 11.505 ;
        RECT 28.710 11.335 36.500 11.505 ;
        RECT 38.700 11.365 46.510 11.535 ;
        RECT 48.480 11.365 56.270 11.535 ;
        RECT 58.420 11.365 66.230 11.535 ;
        RECT 68.190 11.365 75.990 11.535 ;
        RECT 78.500 11.365 86.310 11.535 ;
        RECT 14.680 10.635 15.875 10.805 ;
        RECT 14.680 10.505 14.920 10.635 ;
        RECT 10.065 10.165 10.505 10.405 ;
        RECT 10.930 10.315 11.595 10.485 ;
        RECT 11.765 10.165 12.140 10.485 ;
        RECT 12.435 10.190 13.600 10.475 ;
        RECT 15.705 10.445 15.875 10.635 ;
        RECT 16.045 10.610 16.305 11.185 ;
        RECT 19.015 10.610 19.305 11.335 ;
        RECT 19.500 10.610 19.900 11.165 ;
        RECT 20.145 10.975 20.475 11.335 ;
        RECT 20.645 10.915 21.655 11.165 ;
        RECT 20.645 10.805 20.815 10.915 ;
        RECT 21.485 10.825 21.655 10.915 ;
        RECT 20.075 10.635 20.815 10.805 ;
        RECT 21.990 10.805 22.160 11.165 ;
        RECT 22.330 10.975 22.660 11.335 ;
        RECT 22.830 10.805 23.000 11.165 ;
        RECT 23.170 10.930 23.500 11.335 ;
        RECT 9.150 8.975 9.550 9.955 ;
        RECT 9.725 9.505 9.895 10.115 ;
        RECT 10.335 9.675 10.755 9.995 ;
        RECT 12.435 9.925 12.605 10.190 ;
        RECT 10.985 9.755 12.605 9.925 ;
        RECT 9.725 9.335 10.390 9.505 ;
        RECT 10.985 9.485 11.235 9.755 ;
        RECT 12.830 9.675 13.190 10.005 ;
        RECT 13.430 9.845 13.600 10.190 ;
        RECT 13.770 10.080 14.160 10.410 ;
        RECT 14.350 10.165 14.720 10.335 ;
        RECT 15.150 10.165 15.480 10.445 ;
        RECT 14.350 9.845 14.520 10.165 ;
        RECT 15.310 10.115 15.480 10.165 ;
        RECT 15.705 10.115 15.960 10.445 ;
        RECT 13.430 9.675 14.520 9.845 ;
        RECT 14.690 9.560 15.090 9.995 ;
        RECT 15.705 9.815 15.875 10.115 ;
        RECT 16.130 9.955 16.305 10.610 ;
        RECT 10.220 9.315 10.390 9.335 ;
        RECT 11.640 9.335 12.650 9.505 ;
        RECT 9.720 8.805 10.050 9.165 ;
        RECT 10.220 8.975 11.305 9.315 ;
        RECT 11.640 8.975 11.810 9.335 ;
        RECT 11.980 8.805 12.310 9.165 ;
        RECT 12.480 8.975 12.650 9.335 ;
        RECT 13.355 9.335 14.430 9.505 ;
        RECT 15.285 9.495 15.875 9.815 ;
        RECT 15.285 9.375 15.455 9.495 ;
        RECT 12.820 8.805 13.150 9.185 ;
        RECT 13.355 8.975 13.590 9.335 ;
        RECT 13.760 8.805 14.090 9.165 ;
        RECT 14.260 8.975 14.430 9.335 ;
        RECT 14.680 8.975 15.455 9.375 ;
        RECT 15.625 8.805 15.875 9.290 ;
        RECT 16.045 8.975 16.305 9.955 ;
        RECT 8.580 8.635 16.390 8.805 ;
        RECT 19.015 8.785 19.305 9.950 ;
        RECT 19.500 9.935 19.830 10.610 ;
        RECT 20.075 10.425 20.245 10.635 ;
        RECT 20.000 10.095 20.245 10.425 ;
        RECT 21.280 10.465 21.775 10.655 ;
        RECT 21.990 10.635 23.000 10.805 ;
        RECT 23.770 10.805 23.940 11.165 ;
        RECT 24.110 10.975 24.440 11.335 ;
        RECT 24.610 10.805 24.780 11.165 ;
        RECT 23.770 10.635 24.780 10.805 ;
        RECT 25.030 10.785 25.630 11.165 ;
        RECT 25.895 10.955 26.225 11.335 ;
        RECT 25.030 10.615 26.225 10.785 ;
        RECT 25.030 10.485 25.270 10.615 ;
        RECT 20.415 10.145 20.855 10.385 ;
        RECT 21.280 10.295 21.945 10.465 ;
        RECT 22.115 10.145 22.490 10.465 ;
        RECT 22.785 10.170 23.950 10.455 ;
        RECT 26.055 10.425 26.225 10.615 ;
        RECT 26.395 10.590 26.655 11.165 ;
        RECT 28.795 10.610 29.085 11.335 ;
        RECT 29.260 10.610 29.660 11.165 ;
        RECT 29.905 10.975 30.235 11.335 ;
        RECT 30.405 10.915 31.415 11.165 ;
        RECT 30.405 10.805 30.575 10.915 ;
        RECT 31.245 10.825 31.415 10.915 ;
        RECT 29.835 10.635 30.575 10.805 ;
        RECT 31.750 10.805 31.920 11.165 ;
        RECT 32.090 10.975 32.420 11.335 ;
        RECT 32.590 10.805 32.760 11.165 ;
        RECT 32.930 10.930 33.260 11.335 ;
        RECT 19.500 8.955 19.900 9.935 ;
        RECT 20.075 9.485 20.245 10.095 ;
        RECT 20.685 9.655 21.105 9.975 ;
        RECT 22.785 9.905 22.955 10.170 ;
        RECT 21.335 9.735 22.955 9.905 ;
        RECT 20.075 9.315 20.740 9.485 ;
        RECT 21.335 9.465 21.585 9.735 ;
        RECT 23.180 9.655 23.540 9.985 ;
        RECT 23.780 9.825 23.950 10.170 ;
        RECT 24.120 10.060 24.510 10.390 ;
        RECT 24.700 10.145 25.070 10.315 ;
        RECT 25.500 10.145 25.830 10.425 ;
        RECT 24.700 9.825 24.870 10.145 ;
        RECT 25.660 10.095 25.830 10.145 ;
        RECT 26.055 10.095 26.310 10.425 ;
        RECT 23.780 9.655 24.870 9.825 ;
        RECT 25.040 9.540 25.440 9.975 ;
        RECT 26.055 9.795 26.225 10.095 ;
        RECT 26.480 9.935 26.655 10.590 ;
        RECT 20.570 9.295 20.740 9.315 ;
        RECT 21.990 9.315 23.000 9.485 ;
        RECT 20.070 8.785 20.400 9.145 ;
        RECT 20.570 8.955 21.655 9.295 ;
        RECT 21.990 8.955 22.160 9.315 ;
        RECT 22.330 8.785 22.660 9.145 ;
        RECT 22.830 8.955 23.000 9.315 ;
        RECT 23.705 9.315 24.780 9.485 ;
        RECT 25.635 9.475 26.225 9.795 ;
        RECT 25.635 9.355 25.805 9.475 ;
        RECT 23.170 8.785 23.500 9.165 ;
        RECT 23.705 8.955 23.940 9.315 ;
        RECT 24.110 8.785 24.440 9.145 ;
        RECT 24.610 8.955 24.780 9.315 ;
        RECT 25.030 8.955 25.805 9.355 ;
        RECT 25.975 8.785 26.225 9.270 ;
        RECT 26.395 8.955 26.655 9.935 ;
        RECT 28.795 8.785 29.085 9.950 ;
        RECT 29.260 9.935 29.590 10.610 ;
        RECT 29.835 10.425 30.005 10.635 ;
        RECT 29.760 10.095 30.005 10.425 ;
        RECT 31.040 10.465 31.535 10.655 ;
        RECT 31.750 10.635 32.760 10.805 ;
        RECT 33.530 10.805 33.700 11.165 ;
        RECT 33.870 10.975 34.200 11.335 ;
        RECT 34.370 10.805 34.540 11.165 ;
        RECT 33.530 10.635 34.540 10.805 ;
        RECT 34.790 10.785 35.390 11.165 ;
        RECT 35.655 10.955 35.985 11.335 ;
        RECT 34.790 10.615 35.985 10.785 ;
        RECT 34.790 10.485 35.030 10.615 ;
        RECT 30.175 10.145 30.615 10.385 ;
        RECT 31.040 10.295 31.705 10.465 ;
        RECT 31.875 10.145 32.250 10.465 ;
        RECT 32.545 10.170 33.710 10.455 ;
        RECT 35.815 10.425 35.985 10.615 ;
        RECT 36.155 10.590 36.415 11.165 ;
        RECT 38.785 10.640 39.075 11.365 ;
        RECT 39.270 10.640 39.670 11.195 ;
        RECT 39.915 11.005 40.245 11.365 ;
        RECT 40.415 10.945 41.425 11.195 ;
        RECT 40.415 10.835 40.585 10.945 ;
        RECT 41.255 10.855 41.425 10.945 ;
        RECT 39.845 10.665 40.585 10.835 ;
        RECT 41.760 10.835 41.930 11.195 ;
        RECT 42.100 11.005 42.430 11.365 ;
        RECT 42.600 10.835 42.770 11.195 ;
        RECT 42.940 10.960 43.270 11.365 ;
        RECT 29.260 8.955 29.660 9.935 ;
        RECT 29.835 9.485 30.005 10.095 ;
        RECT 30.445 9.655 30.865 9.975 ;
        RECT 32.545 9.905 32.715 10.170 ;
        RECT 31.095 9.735 32.715 9.905 ;
        RECT 29.835 9.315 30.500 9.485 ;
        RECT 31.095 9.465 31.345 9.735 ;
        RECT 32.940 9.655 33.300 9.985 ;
        RECT 33.540 9.825 33.710 10.170 ;
        RECT 33.880 10.060 34.270 10.390 ;
        RECT 34.460 10.145 34.830 10.315 ;
        RECT 35.260 10.145 35.590 10.425 ;
        RECT 34.460 9.825 34.630 10.145 ;
        RECT 35.420 10.095 35.590 10.145 ;
        RECT 35.815 10.095 36.070 10.425 ;
        RECT 33.540 9.655 34.630 9.825 ;
        RECT 34.800 9.540 35.200 9.975 ;
        RECT 35.815 9.795 35.985 10.095 ;
        RECT 36.240 9.935 36.415 10.590 ;
        RECT 30.330 9.295 30.500 9.315 ;
        RECT 31.750 9.315 32.760 9.485 ;
        RECT 29.830 8.785 30.160 9.145 ;
        RECT 30.330 8.955 31.415 9.295 ;
        RECT 31.750 8.955 31.920 9.315 ;
        RECT 32.090 8.785 32.420 9.145 ;
        RECT 32.590 8.955 32.760 9.315 ;
        RECT 33.465 9.315 34.540 9.485 ;
        RECT 35.395 9.475 35.985 9.795 ;
        RECT 35.395 9.355 35.565 9.475 ;
        RECT 32.930 8.785 33.260 9.165 ;
        RECT 33.465 8.955 33.700 9.315 ;
        RECT 33.870 8.785 34.200 9.145 ;
        RECT 34.370 8.955 34.540 9.315 ;
        RECT 34.790 8.955 35.565 9.355 ;
        RECT 35.735 8.785 35.985 9.270 ;
        RECT 36.155 8.955 36.415 9.935 ;
        RECT 38.785 8.815 39.075 9.980 ;
        RECT 39.270 9.965 39.600 10.640 ;
        RECT 39.845 10.455 40.015 10.665 ;
        RECT 39.770 10.125 40.015 10.455 ;
        RECT 41.050 10.495 41.545 10.685 ;
        RECT 41.760 10.665 42.770 10.835 ;
        RECT 43.540 10.835 43.710 11.195 ;
        RECT 43.880 11.005 44.210 11.365 ;
        RECT 44.380 10.835 44.550 11.195 ;
        RECT 43.540 10.665 44.550 10.835 ;
        RECT 44.800 10.815 45.400 11.195 ;
        RECT 45.665 10.985 45.995 11.365 ;
        RECT 44.800 10.645 45.995 10.815 ;
        RECT 44.800 10.515 45.040 10.645 ;
        RECT 40.185 10.175 40.625 10.415 ;
        RECT 41.050 10.325 41.715 10.495 ;
        RECT 41.885 10.175 42.260 10.495 ;
        RECT 42.555 10.200 43.720 10.485 ;
        RECT 45.825 10.455 45.995 10.645 ;
        RECT 46.165 10.620 46.425 11.195 ;
        RECT 48.565 10.640 48.855 11.365 ;
        RECT 49.030 10.640 49.430 11.195 ;
        RECT 49.675 11.005 50.005 11.365 ;
        RECT 50.175 10.945 51.185 11.195 ;
        RECT 50.175 10.835 50.345 10.945 ;
        RECT 51.015 10.855 51.185 10.945 ;
        RECT 49.605 10.665 50.345 10.835 ;
        RECT 51.520 10.835 51.690 11.195 ;
        RECT 51.860 11.005 52.190 11.365 ;
        RECT 52.360 10.835 52.530 11.195 ;
        RECT 52.700 10.960 53.030 11.365 ;
        RECT 39.270 8.985 39.670 9.965 ;
        RECT 39.845 9.515 40.015 10.125 ;
        RECT 40.455 9.685 40.875 10.005 ;
        RECT 42.555 9.935 42.725 10.200 ;
        RECT 41.105 9.765 42.725 9.935 ;
        RECT 39.845 9.345 40.510 9.515 ;
        RECT 41.105 9.495 41.355 9.765 ;
        RECT 42.950 9.685 43.310 10.015 ;
        RECT 43.550 9.855 43.720 10.200 ;
        RECT 43.890 10.090 44.280 10.420 ;
        RECT 44.470 10.175 44.840 10.345 ;
        RECT 45.270 10.175 45.600 10.455 ;
        RECT 44.470 9.855 44.640 10.175 ;
        RECT 45.430 10.125 45.600 10.175 ;
        RECT 45.825 10.125 46.080 10.455 ;
        RECT 43.550 9.685 44.640 9.855 ;
        RECT 44.810 9.570 45.210 10.005 ;
        RECT 45.825 9.825 45.995 10.125 ;
        RECT 46.250 9.965 46.425 10.620 ;
        RECT 40.340 9.325 40.510 9.345 ;
        RECT 41.760 9.345 42.770 9.515 ;
        RECT 39.840 8.815 40.170 9.175 ;
        RECT 40.340 8.985 41.425 9.325 ;
        RECT 41.760 8.985 41.930 9.345 ;
        RECT 42.100 8.815 42.430 9.175 ;
        RECT 42.600 8.985 42.770 9.345 ;
        RECT 43.475 9.345 44.550 9.515 ;
        RECT 45.405 9.505 45.995 9.825 ;
        RECT 45.405 9.385 45.575 9.505 ;
        RECT 42.940 8.815 43.270 9.195 ;
        RECT 43.475 8.985 43.710 9.345 ;
        RECT 43.880 8.815 44.210 9.175 ;
        RECT 44.380 8.985 44.550 9.345 ;
        RECT 44.800 8.985 45.575 9.385 ;
        RECT 45.745 8.815 45.995 9.300 ;
        RECT 46.165 8.985 46.425 9.965 ;
        RECT 48.565 8.815 48.855 9.980 ;
        RECT 49.030 9.965 49.360 10.640 ;
        RECT 49.605 10.455 49.775 10.665 ;
        RECT 49.530 10.125 49.775 10.455 ;
        RECT 50.810 10.495 51.305 10.685 ;
        RECT 51.520 10.665 52.530 10.835 ;
        RECT 53.300 10.835 53.470 11.195 ;
        RECT 53.640 11.005 53.970 11.365 ;
        RECT 54.140 10.835 54.310 11.195 ;
        RECT 53.300 10.665 54.310 10.835 ;
        RECT 54.560 10.815 55.160 11.195 ;
        RECT 55.425 10.985 55.755 11.365 ;
        RECT 54.560 10.645 55.755 10.815 ;
        RECT 54.560 10.515 54.800 10.645 ;
        RECT 49.945 10.175 50.385 10.415 ;
        RECT 50.810 10.325 51.475 10.495 ;
        RECT 51.645 10.175 52.020 10.495 ;
        RECT 52.315 10.200 53.480 10.485 ;
        RECT 55.585 10.455 55.755 10.645 ;
        RECT 55.925 10.620 56.185 11.195 ;
        RECT 58.505 10.640 58.795 11.365 ;
        RECT 58.990 10.640 59.390 11.195 ;
        RECT 59.635 11.005 59.965 11.365 ;
        RECT 60.135 10.945 61.145 11.195 ;
        RECT 60.135 10.835 60.305 10.945 ;
        RECT 60.975 10.855 61.145 10.945 ;
        RECT 59.565 10.665 60.305 10.835 ;
        RECT 61.480 10.835 61.650 11.195 ;
        RECT 61.820 11.005 62.150 11.365 ;
        RECT 62.320 10.835 62.490 11.195 ;
        RECT 62.660 10.960 62.990 11.365 ;
        RECT 49.030 8.985 49.430 9.965 ;
        RECT 49.605 9.515 49.775 10.125 ;
        RECT 50.215 9.685 50.635 10.005 ;
        RECT 52.315 9.935 52.485 10.200 ;
        RECT 50.865 9.765 52.485 9.935 ;
        RECT 49.605 9.345 50.270 9.515 ;
        RECT 50.865 9.495 51.115 9.765 ;
        RECT 52.710 9.685 53.070 10.015 ;
        RECT 53.310 9.855 53.480 10.200 ;
        RECT 53.650 10.090 54.040 10.420 ;
        RECT 54.230 10.175 54.600 10.345 ;
        RECT 55.030 10.175 55.360 10.455 ;
        RECT 54.230 9.855 54.400 10.175 ;
        RECT 55.190 10.125 55.360 10.175 ;
        RECT 55.585 10.125 55.840 10.455 ;
        RECT 53.310 9.685 54.400 9.855 ;
        RECT 54.570 9.570 54.970 10.005 ;
        RECT 55.585 9.825 55.755 10.125 ;
        RECT 56.010 9.965 56.185 10.620 ;
        RECT 50.100 9.325 50.270 9.345 ;
        RECT 51.520 9.345 52.530 9.515 ;
        RECT 49.600 8.815 49.930 9.175 ;
        RECT 50.100 8.985 51.185 9.325 ;
        RECT 51.520 8.985 51.690 9.345 ;
        RECT 51.860 8.815 52.190 9.175 ;
        RECT 52.360 8.985 52.530 9.345 ;
        RECT 53.235 9.345 54.310 9.515 ;
        RECT 55.165 9.505 55.755 9.825 ;
        RECT 55.165 9.385 55.335 9.505 ;
        RECT 52.700 8.815 53.030 9.195 ;
        RECT 53.235 8.985 53.470 9.345 ;
        RECT 53.640 8.815 53.970 9.175 ;
        RECT 54.140 8.985 54.310 9.345 ;
        RECT 54.560 8.985 55.335 9.385 ;
        RECT 55.505 8.815 55.755 9.300 ;
        RECT 55.925 8.985 56.185 9.965 ;
        RECT 58.505 8.815 58.795 9.980 ;
        RECT 58.990 9.965 59.320 10.640 ;
        RECT 59.565 10.455 59.735 10.665 ;
        RECT 59.490 10.125 59.735 10.455 ;
        RECT 60.770 10.495 61.265 10.685 ;
        RECT 61.480 10.665 62.490 10.835 ;
        RECT 63.260 10.835 63.430 11.195 ;
        RECT 63.600 11.005 63.930 11.365 ;
        RECT 64.100 10.835 64.270 11.195 ;
        RECT 63.260 10.665 64.270 10.835 ;
        RECT 64.520 10.815 65.120 11.195 ;
        RECT 65.385 10.985 65.715 11.365 ;
        RECT 64.520 10.645 65.715 10.815 ;
        RECT 64.520 10.515 64.760 10.645 ;
        RECT 59.905 10.175 60.345 10.415 ;
        RECT 60.770 10.325 61.435 10.495 ;
        RECT 61.605 10.175 61.980 10.495 ;
        RECT 62.275 10.200 63.440 10.485 ;
        RECT 65.545 10.455 65.715 10.645 ;
        RECT 65.885 10.620 66.145 11.195 ;
        RECT 68.275 10.640 68.565 11.365 ;
        RECT 68.750 10.640 69.150 11.195 ;
        RECT 69.395 11.005 69.725 11.365 ;
        RECT 69.895 10.945 70.905 11.195 ;
        RECT 69.895 10.835 70.065 10.945 ;
        RECT 70.735 10.855 70.905 10.945 ;
        RECT 69.325 10.665 70.065 10.835 ;
        RECT 71.240 10.835 71.410 11.195 ;
        RECT 71.580 11.005 71.910 11.365 ;
        RECT 72.080 10.835 72.250 11.195 ;
        RECT 72.420 10.960 72.750 11.365 ;
        RECT 58.990 8.985 59.390 9.965 ;
        RECT 59.565 9.515 59.735 10.125 ;
        RECT 60.175 9.685 60.595 10.005 ;
        RECT 62.275 9.935 62.445 10.200 ;
        RECT 60.825 9.765 62.445 9.935 ;
        RECT 59.565 9.345 60.230 9.515 ;
        RECT 60.825 9.495 61.075 9.765 ;
        RECT 62.670 9.685 63.030 10.015 ;
        RECT 63.270 9.855 63.440 10.200 ;
        RECT 63.610 10.090 64.000 10.420 ;
        RECT 64.190 10.175 64.560 10.345 ;
        RECT 64.990 10.175 65.320 10.455 ;
        RECT 64.190 9.855 64.360 10.175 ;
        RECT 65.150 10.125 65.320 10.175 ;
        RECT 65.545 10.125 65.800 10.455 ;
        RECT 63.270 9.685 64.360 9.855 ;
        RECT 64.530 9.570 64.930 10.005 ;
        RECT 65.545 9.825 65.715 10.125 ;
        RECT 65.970 9.965 66.145 10.620 ;
        RECT 60.060 9.325 60.230 9.345 ;
        RECT 61.480 9.345 62.490 9.515 ;
        RECT 59.560 8.815 59.890 9.175 ;
        RECT 60.060 8.985 61.145 9.325 ;
        RECT 61.480 8.985 61.650 9.345 ;
        RECT 61.820 8.815 62.150 9.175 ;
        RECT 62.320 8.985 62.490 9.345 ;
        RECT 63.195 9.345 64.270 9.515 ;
        RECT 65.125 9.505 65.715 9.825 ;
        RECT 65.125 9.385 65.295 9.505 ;
        RECT 62.660 8.815 62.990 9.195 ;
        RECT 63.195 8.985 63.430 9.345 ;
        RECT 63.600 8.815 63.930 9.175 ;
        RECT 64.100 8.985 64.270 9.345 ;
        RECT 64.520 8.985 65.295 9.385 ;
        RECT 65.465 8.815 65.715 9.300 ;
        RECT 65.885 8.985 66.145 9.965 ;
        RECT 68.275 8.815 68.565 9.980 ;
        RECT 68.750 9.965 69.080 10.640 ;
        RECT 69.325 10.455 69.495 10.665 ;
        RECT 69.250 10.125 69.495 10.455 ;
        RECT 70.530 10.495 71.025 10.685 ;
        RECT 71.240 10.665 72.250 10.835 ;
        RECT 73.020 10.835 73.190 11.195 ;
        RECT 73.360 11.005 73.690 11.365 ;
        RECT 73.860 10.835 74.030 11.195 ;
        RECT 73.020 10.665 74.030 10.835 ;
        RECT 74.280 10.815 74.880 11.195 ;
        RECT 75.145 10.985 75.475 11.365 ;
        RECT 74.280 10.645 75.475 10.815 ;
        RECT 74.280 10.515 74.520 10.645 ;
        RECT 69.665 10.175 70.105 10.415 ;
        RECT 70.530 10.325 71.195 10.495 ;
        RECT 71.365 10.175 71.740 10.495 ;
        RECT 72.035 10.200 73.200 10.485 ;
        RECT 75.305 10.455 75.475 10.645 ;
        RECT 75.645 10.620 75.905 11.195 ;
        RECT 78.585 10.640 78.875 11.365 ;
        RECT 79.070 10.640 79.470 11.195 ;
        RECT 79.715 11.005 80.045 11.365 ;
        RECT 80.215 10.945 81.225 11.195 ;
        RECT 80.215 10.835 80.385 10.945 ;
        RECT 81.055 10.855 81.225 10.945 ;
        RECT 79.645 10.665 80.385 10.835 ;
        RECT 81.560 10.835 81.730 11.195 ;
        RECT 81.900 11.005 82.230 11.365 ;
        RECT 82.400 10.835 82.570 11.195 ;
        RECT 82.740 10.960 83.070 11.365 ;
        RECT 68.750 8.985 69.150 9.965 ;
        RECT 69.325 9.515 69.495 10.125 ;
        RECT 69.935 9.685 70.355 10.005 ;
        RECT 72.035 9.935 72.205 10.200 ;
        RECT 70.585 9.765 72.205 9.935 ;
        RECT 69.325 9.345 69.990 9.515 ;
        RECT 70.585 9.495 70.835 9.765 ;
        RECT 72.430 9.685 72.790 10.015 ;
        RECT 73.030 9.855 73.200 10.200 ;
        RECT 73.370 10.090 73.760 10.420 ;
        RECT 73.950 10.175 74.320 10.345 ;
        RECT 74.750 10.175 75.080 10.455 ;
        RECT 73.950 9.855 74.120 10.175 ;
        RECT 74.910 10.125 75.080 10.175 ;
        RECT 75.305 10.125 75.560 10.455 ;
        RECT 73.030 9.685 74.120 9.855 ;
        RECT 74.290 9.570 74.690 10.005 ;
        RECT 75.305 9.825 75.475 10.125 ;
        RECT 75.730 9.965 75.905 10.620 ;
        RECT 69.820 9.325 69.990 9.345 ;
        RECT 71.240 9.345 72.250 9.515 ;
        RECT 69.320 8.815 69.650 9.175 ;
        RECT 69.820 8.985 70.905 9.325 ;
        RECT 71.240 8.985 71.410 9.345 ;
        RECT 71.580 8.815 71.910 9.175 ;
        RECT 72.080 8.985 72.250 9.345 ;
        RECT 72.955 9.345 74.030 9.515 ;
        RECT 74.885 9.505 75.475 9.825 ;
        RECT 74.885 9.385 75.055 9.505 ;
        RECT 72.420 8.815 72.750 9.195 ;
        RECT 72.955 8.985 73.190 9.345 ;
        RECT 73.360 8.815 73.690 9.175 ;
        RECT 73.860 8.985 74.030 9.345 ;
        RECT 74.280 8.985 75.055 9.385 ;
        RECT 75.225 8.815 75.475 9.300 ;
        RECT 75.645 8.985 75.905 9.965 ;
        RECT 78.585 8.815 78.875 9.980 ;
        RECT 79.070 9.965 79.400 10.640 ;
        RECT 79.645 10.455 79.815 10.665 ;
        RECT 79.570 10.125 79.815 10.455 ;
        RECT 80.850 10.495 81.345 10.685 ;
        RECT 81.560 10.665 82.570 10.835 ;
        RECT 83.340 10.835 83.510 11.195 ;
        RECT 83.680 11.005 84.010 11.365 ;
        RECT 84.180 10.835 84.350 11.195 ;
        RECT 83.340 10.665 84.350 10.835 ;
        RECT 84.600 10.815 85.200 11.195 ;
        RECT 85.465 10.985 85.795 11.365 ;
        RECT 84.600 10.645 85.795 10.815 ;
        RECT 84.600 10.515 84.840 10.645 ;
        RECT 79.985 10.175 80.425 10.415 ;
        RECT 80.850 10.325 81.515 10.495 ;
        RECT 81.685 10.175 82.060 10.495 ;
        RECT 82.355 10.200 83.520 10.485 ;
        RECT 85.625 10.455 85.795 10.645 ;
        RECT 85.965 10.620 86.225 11.195 ;
        RECT 79.070 8.985 79.470 9.965 ;
        RECT 79.645 9.515 79.815 10.125 ;
        RECT 80.255 9.685 80.675 10.005 ;
        RECT 82.355 9.935 82.525 10.200 ;
        RECT 80.905 9.765 82.525 9.935 ;
        RECT 79.645 9.345 80.310 9.515 ;
        RECT 80.905 9.495 81.155 9.765 ;
        RECT 82.750 9.685 83.110 10.015 ;
        RECT 83.350 9.855 83.520 10.200 ;
        RECT 83.690 10.090 84.080 10.420 ;
        RECT 84.270 10.175 84.640 10.345 ;
        RECT 85.070 10.175 85.400 10.455 ;
        RECT 84.270 9.855 84.440 10.175 ;
        RECT 85.230 10.125 85.400 10.175 ;
        RECT 85.625 10.125 85.880 10.455 ;
        RECT 83.350 9.685 84.440 9.855 ;
        RECT 84.610 9.570 85.010 10.005 ;
        RECT 85.625 9.825 85.795 10.125 ;
        RECT 86.050 9.965 86.225 10.620 ;
        RECT 80.140 9.325 80.310 9.345 ;
        RECT 81.560 9.345 82.570 9.515 ;
        RECT 79.640 8.815 79.970 9.175 ;
        RECT 80.140 8.985 81.225 9.325 ;
        RECT 81.560 8.985 81.730 9.345 ;
        RECT 81.900 8.815 82.230 9.175 ;
        RECT 82.400 8.985 82.570 9.345 ;
        RECT 83.275 9.345 84.350 9.515 ;
        RECT 85.205 9.505 85.795 9.825 ;
        RECT 85.205 9.385 85.375 9.505 ;
        RECT 82.740 8.815 83.070 9.195 ;
        RECT 83.275 8.985 83.510 9.345 ;
        RECT 83.680 8.815 84.010 9.175 ;
        RECT 84.180 8.985 84.350 9.345 ;
        RECT 84.600 8.985 85.375 9.385 ;
        RECT 85.545 8.815 85.795 9.300 ;
        RECT 85.965 8.985 86.225 9.965 ;
        RECT 18.930 8.615 26.740 8.785 ;
        RECT 28.710 8.615 36.500 8.785 ;
        RECT 38.700 8.645 46.510 8.815 ;
        RECT 48.480 8.645 56.270 8.815 ;
        RECT 58.420 8.645 66.230 8.815 ;
        RECT 68.190 8.645 75.990 8.815 ;
        RECT 78.500 8.645 86.310 8.815 ;
      LAYER met1 ;
        RECT 92.950 219.140 95.640 220.840 ;
        RECT 92.740 209.740 93.220 217.550 ;
        RECT 94.330 216.220 94.680 219.140 ;
        RECT 92.660 201.180 93.140 207.620 ;
        RECT 94.280 206.730 94.690 210.250 ;
        RECT 95.460 209.740 95.940 217.550 ;
        RECT 92.700 194.040 93.180 198.640 ;
        RECT 94.230 197.770 94.570 202.550 ;
        RECT 95.380 201.180 95.860 207.620 ;
        RECT 92.770 188.650 93.250 192.330 ;
        RECT 94.320 191.420 94.730 195.570 ;
        RECT 95.420 194.040 95.900 198.640 ;
        RECT 92.830 183.820 93.310 186.560 ;
        RECT 94.360 185.990 94.670 189.770 ;
        RECT 95.490 188.650 95.970 192.330 ;
        RECT 94.350 185.720 94.760 185.990 ;
        RECT 94.430 184.340 94.750 184.640 ;
        RECT 92.870 180.300 93.350 182.140 ;
        RECT 94.490 181.180 94.720 184.340 ;
        RECT 95.550 183.820 96.030 186.560 ;
        RECT 94.450 180.880 94.770 181.180 ;
        RECT 94.480 180.400 94.790 180.730 ;
        RECT 94.555 179.395 94.765 180.400 ;
        RECT 95.590 180.300 96.070 182.140 ;
        RECT 94.350 179.185 94.765 179.395 ;
        RECT 92.090 166.930 92.570 176.130 ;
        RECT 93.160 175.510 93.680 175.630 ;
        RECT 93.160 175.260 93.770 175.510 ;
        RECT 93.160 175.250 93.680 175.260 ;
        RECT 93.305 173.020 93.660 175.250 ;
        RECT 94.350 174.170 94.560 179.185 ;
        RECT 94.230 173.870 94.670 174.170 ;
        RECT 93.305 172.665 94.335 173.020 ;
        RECT 93.405 171.605 93.635 171.895 ;
        RECT 93.065 171.170 93.295 171.460 ;
        RECT 93.110 169.890 93.250 171.170 ;
        RECT 93.065 169.600 93.295 169.890 ;
        RECT 93.110 167.790 93.250 169.600 ;
        RECT 93.450 169.375 93.590 171.605 ;
        RECT 93.405 169.085 93.635 169.375 ;
        RECT 93.450 168.185 93.590 169.085 ;
        RECT 93.980 168.300 94.335 172.665 ;
        RECT 93.405 167.895 93.635 168.185 ;
        RECT 93.065 167.500 93.295 167.790 ;
        RECT 93.575 166.390 94.305 167.385 ;
        RECT 94.810 166.930 95.290 176.130 ;
        RECT 93.570 166.080 94.305 166.390 ;
        RECT 92.130 155.400 92.610 164.600 ;
        RECT 93.570 164.100 93.920 166.080 ;
        RECT 93.200 164.000 93.920 164.100 ;
        RECT 93.200 163.730 94.375 164.000 ;
        RECT 93.200 163.720 93.720 163.730 ;
        RECT 93.445 160.075 93.675 160.365 ;
        RECT 93.105 159.640 93.335 159.930 ;
        RECT 93.150 158.360 93.290 159.640 ;
        RECT 93.105 158.070 93.335 158.360 ;
        RECT 93.150 156.260 93.290 158.070 ;
        RECT 93.490 157.845 93.630 160.075 ;
        RECT 93.445 157.555 93.675 157.845 ;
        RECT 93.490 156.655 93.630 157.555 ;
        RECT 94.020 156.770 94.375 163.730 ;
        RECT 93.445 156.365 93.675 156.655 ;
        RECT 93.105 155.970 93.335 156.260 ;
        RECT 93.615 154.410 94.345 155.855 ;
        RECT 94.850 155.400 95.330 164.600 ;
        RECT 93.600 153.890 94.345 154.410 ;
        RECT 92.170 144.330 92.650 153.530 ;
        RECT 93.600 153.030 93.770 153.890 ;
        RECT 93.240 152.910 93.770 153.030 ;
        RECT 94.060 152.910 94.415 152.930 ;
        RECT 93.240 152.660 94.415 152.910 ;
        RECT 93.240 152.650 93.760 152.660 ;
        RECT 93.485 149.005 93.715 149.295 ;
        RECT 93.145 148.570 93.375 148.860 ;
        RECT 93.190 147.290 93.330 148.570 ;
        RECT 93.145 147.000 93.375 147.290 ;
        RECT 93.190 145.190 93.330 147.000 ;
        RECT 93.530 146.775 93.670 149.005 ;
        RECT 93.485 146.485 93.715 146.775 ;
        RECT 93.530 145.585 93.670 146.485 ;
        RECT 94.060 145.700 94.415 152.660 ;
        RECT 93.485 145.295 93.715 145.585 ;
        RECT 93.145 144.900 93.375 145.190 ;
        RECT 93.655 143.710 94.385 144.785 ;
        RECT 94.890 144.330 95.370 153.530 ;
        RECT 93.650 143.040 94.385 143.710 ;
        RECT 92.080 133.330 92.560 142.530 ;
        RECT 93.650 142.030 93.830 143.040 ;
        RECT 93.150 141.910 93.830 142.030 ;
        RECT 93.970 141.910 94.325 141.930 ;
        RECT 93.150 141.660 94.325 141.910 ;
        RECT 93.150 141.650 93.670 141.660 ;
        RECT 93.395 138.005 93.625 138.295 ;
        RECT 93.055 137.570 93.285 137.860 ;
        RECT 93.100 136.290 93.240 137.570 ;
        RECT 93.055 136.000 93.285 136.290 ;
        RECT 93.100 134.190 93.240 136.000 ;
        RECT 93.440 135.775 93.580 138.005 ;
        RECT 93.395 135.485 93.625 135.775 ;
        RECT 93.440 134.585 93.580 135.485 ;
        RECT 93.970 134.700 94.325 141.660 ;
        RECT 93.395 134.295 93.625 134.585 ;
        RECT 93.055 133.900 93.285 134.190 ;
        RECT 93.565 132.340 94.295 133.785 ;
        RECT 94.800 133.330 95.280 142.530 ;
        RECT 93.550 131.820 94.295 132.340 ;
        RECT 92.120 122.260 92.600 131.460 ;
        RECT 93.550 130.960 93.720 131.820 ;
        RECT 93.190 130.840 93.720 130.960 ;
        RECT 94.010 130.840 94.365 130.860 ;
        RECT 93.190 130.590 94.365 130.840 ;
        RECT 93.190 130.580 93.710 130.590 ;
        RECT 93.435 126.935 93.665 127.225 ;
        RECT 93.095 126.500 93.325 126.790 ;
        RECT 93.140 125.220 93.280 126.500 ;
        RECT 93.095 124.930 93.325 125.220 ;
        RECT 93.140 123.120 93.280 124.930 ;
        RECT 93.480 124.705 93.620 126.935 ;
        RECT 93.435 124.415 93.665 124.705 ;
        RECT 93.480 123.515 93.620 124.415 ;
        RECT 94.010 123.630 94.365 130.590 ;
        RECT 93.435 123.225 93.665 123.515 ;
        RECT 93.095 122.830 93.325 123.120 ;
        RECT 93.605 121.710 94.335 122.715 ;
        RECT 94.840 122.260 95.320 131.460 ;
        RECT 37.730 116.700 46.930 117.180 ;
        RECT 48.800 116.740 58.000 117.220 ;
        RECT 59.800 116.650 69.000 117.130 ;
        RECT 70.870 116.690 80.070 117.170 ;
        RECT 82.400 116.730 91.600 117.210 ;
        RECT 38.300 116.160 38.590 116.205 ;
        RECT 40.400 116.160 40.690 116.205 ;
        RECT 41.970 116.160 42.260 116.205 ;
        RECT 38.300 116.020 42.260 116.160 ;
        RECT 49.370 116.200 49.660 116.245 ;
        RECT 51.470 116.200 51.760 116.245 ;
        RECT 53.040 116.200 53.330 116.245 ;
        RECT 38.300 115.975 38.590 116.020 ;
        RECT 40.400 115.975 40.690 116.020 ;
        RECT 41.970 115.975 42.260 116.020 ;
        RECT 38.695 115.820 38.985 115.865 ;
        RECT 39.885 115.820 40.175 115.865 ;
        RECT 42.405 115.820 42.695 115.865 ;
        RECT 31.345 114.965 38.185 115.695 ;
        RECT 38.695 115.680 42.695 115.820 ;
        RECT 38.695 115.635 38.985 115.680 ;
        RECT 39.885 115.635 40.175 115.680 ;
        RECT 42.405 115.635 42.695 115.680 ;
        RECT 46.050 115.750 46.430 116.110 ;
        RECT 49.370 116.060 53.330 116.200 ;
        RECT 49.370 116.015 49.660 116.060 ;
        RECT 51.470 116.015 51.760 116.060 ;
        RECT 53.040 116.015 53.330 116.060 ;
        RECT 49.765 115.860 50.055 115.905 ;
        RECT 50.955 115.860 51.245 115.905 ;
        RECT 53.475 115.860 53.765 115.905 ;
        RECT 46.050 115.735 47.810 115.750 ;
        RECT 46.050 115.590 49.255 115.735 ;
        RECT 49.765 115.720 53.765 115.860 ;
        RECT 49.765 115.675 50.055 115.720 ;
        RECT 50.955 115.675 51.245 115.720 ;
        RECT 53.475 115.675 53.765 115.720 ;
        RECT 57.120 115.650 57.500 116.150 ;
        RECT 60.370 116.110 60.660 116.155 ;
        RECT 62.470 116.110 62.760 116.155 ;
        RECT 64.040 116.110 64.330 116.155 ;
        RECT 60.370 115.970 64.330 116.110 ;
        RECT 71.440 116.150 71.730 116.195 ;
        RECT 73.540 116.150 73.830 116.195 ;
        RECT 75.110 116.150 75.400 116.195 ;
        RECT 60.370 115.925 60.660 115.970 ;
        RECT 62.470 115.925 62.760 115.970 ;
        RECT 64.040 115.925 64.330 115.970 ;
        RECT 60.765 115.770 61.055 115.815 ;
        RECT 61.955 115.770 62.245 115.815 ;
        RECT 64.475 115.770 64.765 115.815 ;
        RECT 57.120 115.645 59.180 115.650 ;
        RECT 57.120 115.630 60.255 115.645 ;
        RECT 46.060 115.580 49.255 115.590 ;
        RECT 46.060 115.290 46.310 115.580 ;
        RECT 31.345 92.425 32.075 114.965 ;
        RECT 39.100 114.935 46.330 115.290 ;
        RECT 47.290 115.005 49.255 115.580 ;
        RECT 57.130 115.470 60.255 115.630 ;
        RECT 60.765 115.630 64.765 115.770 ;
        RECT 60.765 115.585 61.055 115.630 ;
        RECT 61.955 115.585 62.245 115.630 ;
        RECT 64.475 115.585 64.765 115.630 ;
        RECT 68.120 115.700 68.500 116.060 ;
        RECT 71.440 116.010 75.400 116.150 ;
        RECT 82.970 116.190 83.260 116.235 ;
        RECT 85.070 116.190 85.360 116.235 ;
        RECT 86.640 116.190 86.930 116.235 ;
        RECT 71.440 115.965 71.730 116.010 ;
        RECT 73.540 115.965 73.830 116.010 ;
        RECT 75.110 115.965 75.400 116.010 ;
        RECT 71.835 115.810 72.125 115.855 ;
        RECT 73.025 115.810 73.315 115.855 ;
        RECT 75.545 115.810 75.835 115.855 ;
        RECT 68.120 115.685 69.880 115.700 ;
        RECT 68.120 115.540 71.325 115.685 ;
        RECT 71.835 115.670 75.835 115.810 ;
        RECT 71.835 115.625 72.125 115.670 ;
        RECT 73.025 115.625 73.315 115.670 ;
        RECT 75.545 115.625 75.835 115.670 ;
        RECT 79.190 115.730 79.570 116.100 ;
        RECT 82.970 116.050 86.930 116.190 ;
        RECT 82.970 116.005 83.260 116.050 ;
        RECT 85.070 116.005 85.360 116.050 ;
        RECT 86.640 116.005 86.930 116.050 ;
        RECT 83.365 115.850 83.655 115.895 ;
        RECT 84.555 115.850 84.845 115.895 ;
        RECT 87.075 115.850 87.365 115.895 ;
        RECT 90.720 115.870 91.100 116.140 ;
        RECT 93.615 115.870 94.335 121.710 ;
        RECT 79.190 115.725 81.860 115.730 ;
        RECT 79.190 115.580 82.855 115.725 ;
        RECT 83.365 115.710 87.365 115.850 ;
        RECT 83.365 115.665 83.655 115.710 ;
        RECT 84.555 115.665 84.845 115.710 ;
        RECT 87.075 115.665 87.365 115.710 ;
        RECT 57.130 115.330 57.380 115.470 ;
        RECT 50.170 114.975 57.400 115.330 ;
        RECT 58.510 114.915 60.255 115.470 ;
        RECT 68.130 115.530 71.325 115.540 ;
        RECT 68.130 115.240 68.380 115.530 ;
        RECT 61.170 114.885 68.400 115.240 ;
        RECT 69.360 114.955 71.325 115.530 ;
        RECT 79.200 115.380 82.855 115.580 ;
        RECT 79.200 115.280 79.470 115.380 ;
        RECT 72.240 114.925 79.470 115.280 ;
        RECT 81.550 114.995 82.855 115.380 ;
        RECT 90.700 115.320 94.335 115.870 ;
        RECT 83.770 115.150 94.335 115.320 ;
        RECT 83.770 114.965 91.000 115.150 ;
        RECT 37.730 113.980 46.930 114.460 ;
        RECT 48.800 114.020 58.000 114.500 ;
        RECT 59.800 113.930 69.000 114.410 ;
        RECT 70.870 113.970 80.070 114.450 ;
        RECT 82.400 114.010 91.600 114.490 ;
        RECT 31.345 91.695 130.315 92.425 ;
        RECT 47.150 88.730 48.910 89.210 ;
        RECT 77.405 87.990 79.215 88.470 ;
        RECT 81.335 88.180 83.105 88.660 ;
        RECT 85.665 88.190 87.475 88.670 ;
        RECT 89.555 88.490 91.315 88.620 ;
        RECT 95.135 88.530 96.925 88.630 ;
        RECT 89.545 88.160 91.315 88.490 ;
        RECT 95.125 88.200 96.925 88.530 ;
        RECT 89.555 88.140 91.315 88.160 ;
        RECT 95.135 88.150 96.925 88.200 ;
        RECT 99.465 88.160 101.295 88.640 ;
        RECT 103.315 88.110 105.135 88.590 ;
        RECT 106.825 88.100 108.665 88.580 ;
        RECT 110.745 88.110 112.575 88.590 ;
        RECT 115.035 88.060 116.865 88.540 ;
        RECT 33.015 87.485 47.695 87.935 ;
        RECT 47.865 87.485 68.665 87.935 ;
        RECT 47.150 86.430 48.910 86.490 ;
        RECT 47.150 86.100 48.980 86.430 ;
        RECT 47.150 86.010 48.910 86.100 ;
        RECT 45.225 85.270 57.410 85.275 ;
        RECT 45.180 85.205 57.410 85.270 ;
        RECT 43.935 84.885 57.410 85.205 ;
        RECT 43.935 84.820 47.485 84.885 ;
        RECT 43.935 84.815 45.000 84.820 ;
        RECT 45.800 84.815 47.485 84.820 ;
        RECT 21.880 83.080 25.560 83.170 ;
        RECT 21.820 82.750 25.560 83.080 ;
        RECT 21.880 82.690 25.560 82.750 ;
        RECT 22.730 81.190 23.030 82.690 ;
        RECT 29.730 82.020 30.740 82.190 ;
        RECT 25.160 81.690 31.295 82.020 ;
        RECT 29.730 81.560 30.740 81.690 ;
        RECT 23.180 81.260 23.730 81.540 ;
        RECT 23.350 80.450 23.505 81.260 ;
        RECT 21.880 80.380 25.560 80.450 ;
        RECT 21.800 80.050 25.560 80.380 ;
        RECT 21.880 79.970 25.560 80.050 ;
        RECT 22.380 78.970 25.130 79.450 ;
        RECT 22.870 77.570 23.250 77.930 ;
        RECT 23.880 77.850 24.150 78.970 ;
        RECT 30.965 78.165 31.295 81.690 ;
        RECT 33.040 78.780 36.720 78.900 ;
        RECT 32.740 78.450 36.720 78.780 ;
        RECT 33.040 78.420 36.720 78.450 ;
        RECT 22.920 76.730 23.190 77.570 ;
        RECT 23.830 77.540 24.170 77.850 ;
        RECT 30.965 77.835 35.235 78.165 ;
        RECT 33.955 77.820 34.285 77.835 ;
        RECT 24.790 77.180 25.220 77.550 ;
        RECT 25.970 77.290 34.280 77.580 ;
        RECT 25.970 77.260 34.285 77.290 ;
        RECT 23.830 76.730 24.170 76.740 ;
        RECT 22.380 76.250 25.130 76.730 ;
        RECT 21.930 74.870 25.610 75.350 ;
        RECT 22.780 73.370 23.080 74.870 ;
        RECT 25.970 74.710 26.290 77.260 ;
        RECT 32.890 76.710 33.410 77.120 ;
        RECT 33.955 76.950 34.285 77.260 ;
        RECT 34.450 76.570 34.740 76.650 ;
        RECT 28.750 76.370 31.510 76.400 ;
        RECT 28.740 76.040 31.510 76.370 ;
        RECT 31.740 76.350 34.740 76.570 ;
        RECT 28.750 75.920 31.510 76.040 ;
        RECT 31.750 75.780 32.150 76.350 ;
        RECT 34.450 76.320 34.740 76.350 ;
        RECT 34.905 76.330 35.235 77.835 ;
        RECT 35.890 77.200 36.170 77.220 ;
        RECT 35.890 76.950 38.095 77.200 ;
        RECT 35.890 76.930 36.170 76.950 ;
        RECT 36.735 76.940 36.985 76.950 ;
        RECT 33.040 76.110 36.720 76.180 ;
        RECT 32.730 75.780 36.720 76.110 ;
        RECT 25.200 74.390 26.290 74.710 ;
        RECT 26.450 75.400 30.100 75.660 ;
        RECT 30.520 75.490 32.150 75.780 ;
        RECT 33.040 75.700 36.720 75.780 ;
        RECT 23.230 73.440 23.780 73.720 ;
        RECT 23.400 72.630 23.555 73.440 ;
        RECT 21.930 72.150 25.610 72.630 ;
        RECT 22.430 71.150 25.180 71.630 ;
        RECT 22.920 69.750 23.300 70.120 ;
        RECT 23.940 70.030 24.170 71.150 ;
        RECT 22.960 68.910 23.230 69.750 ;
        RECT 23.880 69.720 24.220 70.030 ;
        RECT 24.830 69.100 25.690 69.570 ;
        RECT 22.430 68.430 25.180 68.910 ;
        RECT 21.890 66.530 25.570 67.010 ;
        RECT 26.450 66.830 26.710 75.400 ;
        RECT 29.840 74.780 30.100 75.400 ;
        RECT 28.850 74.755 29.530 74.760 ;
        RECT 27.810 74.390 29.530 74.755 ;
        RECT 29.700 74.450 30.100 74.780 ;
        RECT 27.810 74.365 29.225 74.390 ;
        RECT 27.810 69.855 28.200 74.365 ;
        RECT 28.750 73.580 31.510 73.680 ;
        RECT 28.740 73.250 31.510 73.580 ;
        RECT 28.750 73.200 31.510 73.250 ;
        RECT 36.735 73.365 36.985 73.370 ;
        RECT 37.845 73.365 38.095 76.950 ;
        RECT 36.735 73.115 38.095 73.365 ;
        RECT 28.660 71.090 32.340 71.570 ;
        RECT 36.735 70.885 36.985 73.115 ;
        RECT 38.610 71.010 41.830 71.490 ;
        RECT 36.735 70.860 36.990 70.885 ;
        RECT 36.735 70.625 40.370 70.860 ;
        RECT 36.950 70.620 40.370 70.625 ;
        RECT 43.935 70.480 44.325 84.815 ;
        RECT 46.210 82.710 49.890 83.190 ;
        RECT 47.060 81.210 47.360 82.710 ;
        RECT 54.060 82.040 55.070 82.210 ;
        RECT 49.490 81.710 55.625 82.040 ;
        RECT 54.060 81.580 55.070 81.710 ;
        RECT 47.510 81.280 48.060 81.560 ;
        RECT 47.680 80.470 47.835 81.280 ;
        RECT 46.210 80.440 49.890 80.470 ;
        RECT 46.160 80.110 49.890 80.440 ;
        RECT 46.210 79.990 49.890 80.110 ;
        RECT 46.710 78.990 49.460 79.470 ;
        RECT 47.200 77.590 47.580 77.950 ;
        RECT 48.210 77.870 48.480 78.990 ;
        RECT 55.295 78.185 55.625 81.710 ;
        RECT 57.370 78.860 61.050 78.920 ;
        RECT 57.050 78.530 61.050 78.860 ;
        RECT 57.370 78.440 61.050 78.530 ;
        RECT 47.250 76.750 47.520 77.590 ;
        RECT 48.160 77.560 48.500 77.870 ;
        RECT 55.295 77.855 59.565 78.185 ;
        RECT 58.285 77.840 58.615 77.855 ;
        RECT 49.120 77.200 49.550 77.570 ;
        RECT 50.300 77.310 58.610 77.600 ;
        RECT 50.300 77.280 58.615 77.310 ;
        RECT 48.160 76.750 48.500 76.760 ;
        RECT 46.710 76.270 49.460 76.750 ;
        RECT 46.260 74.890 49.940 75.370 ;
        RECT 47.110 73.390 47.410 74.890 ;
        RECT 50.300 74.730 50.620 77.280 ;
        RECT 57.220 76.730 57.740 77.140 ;
        RECT 58.285 76.970 58.615 77.280 ;
        RECT 58.780 76.590 59.070 76.670 ;
        RECT 53.080 75.940 55.840 76.420 ;
        RECT 56.070 76.370 59.070 76.590 ;
        RECT 56.080 75.800 56.480 76.370 ;
        RECT 58.780 76.340 59.070 76.370 ;
        RECT 59.235 76.350 59.565 77.855 ;
        RECT 60.220 77.220 60.500 77.240 ;
        RECT 60.220 76.970 62.425 77.220 ;
        RECT 60.220 76.950 60.500 76.970 ;
        RECT 61.065 76.950 61.315 76.970 ;
        RECT 57.370 76.150 61.050 76.200 ;
        RECT 57.020 75.820 61.050 76.150 ;
        RECT 49.530 74.410 50.620 74.730 ;
        RECT 50.780 75.420 54.430 75.680 ;
        RECT 54.850 75.510 56.480 75.800 ;
        RECT 57.370 75.720 61.050 75.820 ;
        RECT 47.560 73.460 48.110 73.740 ;
        RECT 47.730 72.650 47.885 73.460 ;
        RECT 46.260 72.170 49.940 72.650 ;
        RECT 46.750 71.170 49.510 71.650 ;
        RECT 37.230 70.150 40.570 70.450 ;
        RECT 29.115 69.855 29.505 70.145 ;
        RECT 37.230 70.090 37.600 70.150 ;
        RECT 27.810 69.465 29.505 69.855 ;
        RECT 22.740 65.030 23.040 66.530 ;
        RECT 26.450 66.480 26.880 66.830 ;
        RECT 26.450 66.140 26.710 66.480 ;
        RECT 25.180 65.880 26.710 66.140 ;
        RECT 27.810 65.425 28.200 69.465 ;
        RECT 30.010 68.990 30.360 69.680 ;
        RECT 30.500 69.000 30.840 69.930 ;
        RECT 31.010 69.020 31.370 69.940 ;
        RECT 31.900 68.990 33.330 69.360 ;
        RECT 33.970 69.220 36.710 69.700 ;
        RECT 37.230 69.650 37.590 70.090 ;
        RECT 38.180 69.870 38.710 69.880 ;
        RECT 32.925 68.925 33.330 68.990 ;
        RECT 37.230 68.930 37.580 69.650 ;
        RECT 38.180 69.280 39.030 69.870 ;
        RECT 39.180 69.790 39.880 69.960 ;
        RECT 40.210 69.860 40.570 70.150 ;
        RECT 40.910 70.090 44.325 70.480 ;
        RECT 43.010 69.950 43.190 70.090 ;
        RECT 39.180 69.450 39.870 69.790 ;
        RECT 40.100 69.520 40.570 69.860 ;
        RECT 47.250 69.770 47.630 70.140 ;
        RECT 48.270 70.050 48.500 71.170 ;
        RECT 47.290 68.930 47.560 69.770 ;
        RECT 48.210 69.740 48.550 70.050 ;
        RECT 49.160 69.120 50.020 69.590 ;
        RECT 28.660 68.370 32.340 68.850 ;
        RECT 32.925 68.555 35.315 68.925 ;
        RECT 35.600 68.570 37.580 68.930 ;
        RECT 32.720 67.515 34.465 67.885 ;
        RECT 29.280 66.880 32.040 67.360 ;
        RECT 30.600 66.340 31.090 66.720 ;
        RECT 32.720 66.490 33.090 67.515 ;
        RECT 34.945 67.445 35.315 68.555 ;
        RECT 38.200 68.290 41.830 68.770 ;
        RECT 46.750 68.450 49.510 68.930 ;
        RECT 38.200 68.280 38.670 68.290 ;
        RECT 33.970 66.500 36.710 66.980 ;
        RECT 46.220 66.550 49.900 67.030 ;
        RECT 50.780 66.850 51.040 75.420 ;
        RECT 54.170 74.800 54.430 75.420 ;
        RECT 53.180 74.775 53.860 74.780 ;
        RECT 52.140 74.410 53.860 74.775 ;
        RECT 54.030 74.470 54.430 74.800 ;
        RECT 52.140 74.385 53.555 74.410 ;
        RECT 52.140 69.875 52.530 74.385 ;
        RECT 62.175 73.705 62.425 76.970 ;
        RECT 61.705 73.700 62.425 73.705 ;
        RECT 53.080 73.220 55.840 73.700 ;
        RECT 61.045 73.455 62.425 73.700 ;
        RECT 68.215 73.485 68.665 87.485 ;
        RECT 81.995 87.330 82.305 87.390 ;
        RECT 76.800 87.180 78.415 87.290 ;
        RECT 74.800 87.035 75.130 87.180 ;
        RECT 75.610 87.035 78.415 87.180 ;
        RECT 74.800 81.830 74.945 87.035 ;
        RECT 76.800 86.840 78.415 87.035 ;
        RECT 78.565 87.055 79.510 87.240 ;
        RECT 79.715 87.180 82.305 87.330 ;
        RECT 79.715 87.055 79.865 87.180 ;
        RECT 80.935 87.170 81.085 87.180 ;
        RECT 78.565 86.905 79.865 87.055 ;
        RECT 81.995 87.050 82.305 87.180 ;
        RECT 82.465 87.040 86.675 87.490 ;
        RECT 86.825 87.070 90.515 87.440 ;
        RECT 90.665 87.370 91.005 87.450 ;
        RECT 90.665 87.360 95.895 87.370 ;
        RECT 90.665 87.090 96.125 87.360 ;
        RECT 90.665 87.030 91.005 87.090 ;
        RECT 95.815 87.020 96.125 87.090 ;
        RECT 96.285 87.010 100.495 87.460 ;
        RECT 104.485 87.415 104.815 87.420 ;
        RECT 100.645 87.040 104.335 87.410 ;
        RECT 104.485 87.340 105.535 87.415 ;
        RECT 104.485 87.310 107.125 87.340 ;
        RECT 104.485 87.110 107.405 87.310 ;
        RECT 104.485 87.000 104.815 87.110 ;
        RECT 106.525 87.100 107.405 87.110 ;
        RECT 107.095 86.970 107.405 87.100 ;
        RECT 107.565 86.960 111.775 87.410 ;
        RECT 115.765 87.365 116.095 87.370 ;
        RECT 111.925 86.990 115.615 87.360 ;
        RECT 115.765 87.215 117.160 87.365 ;
        RECT 115.765 86.950 116.095 87.215 ;
        RECT 78.565 86.870 79.510 86.905 ;
        RECT 77.405 85.270 79.215 85.750 ;
        RECT 81.335 85.460 83.105 85.940 ;
        RECT 85.665 85.470 87.475 85.950 ;
        RECT 89.555 85.800 91.315 85.900 ;
        RECT 89.525 85.470 91.315 85.800 ;
        RECT 89.555 85.420 91.315 85.470 ;
        RECT 95.135 85.430 96.925 85.910 ;
        RECT 99.465 85.440 101.295 85.920 ;
        RECT 103.315 85.390 105.135 85.870 ;
        RECT 106.825 85.380 108.665 85.860 ;
        RECT 110.745 85.390 112.575 85.870 ;
        RECT 115.035 85.340 116.865 85.820 ;
        RECT 117.010 84.685 117.160 87.215 ;
        RECT 117.010 84.530 117.395 84.685 ;
        RECT 117.015 84.385 117.395 84.530 ;
        RECT 81.230 83.230 83.060 83.710 ;
        RECT 85.520 83.180 87.350 83.660 ;
        RECT 89.430 83.190 91.270 83.670 ;
        RECT 92.960 83.180 94.780 83.660 ;
        RECT 96.800 83.130 98.630 83.610 ;
        RECT 101.170 83.140 102.960 83.620 ;
        RECT 106.780 83.580 108.540 83.630 ;
        RECT 106.780 83.250 108.570 83.580 ;
        RECT 106.780 83.150 108.540 83.250 ;
        RECT 110.620 83.100 112.430 83.580 ;
        RECT 114.990 83.110 116.760 83.590 ;
        RECT 82.000 81.835 82.330 82.100 ;
        RECT 81.120 81.830 82.330 81.835 ;
        RECT 74.800 81.685 75.130 81.830 ;
        RECT 75.610 81.685 82.330 81.830 ;
        RECT 82.480 81.690 86.170 82.060 ;
        RECT 82.000 81.680 82.330 81.685 ;
        RECT 86.320 81.640 90.530 82.090 ;
        RECT 90.690 81.950 91.000 82.080 ;
        RECT 90.690 81.940 91.570 81.950 ;
        RECT 93.280 81.940 93.610 82.050 ;
        RECT 90.690 81.740 93.610 81.940 ;
        RECT 90.970 81.710 93.610 81.740 ;
        RECT 92.560 81.635 93.610 81.710 ;
        RECT 93.760 81.640 97.450 82.010 ;
        RECT 93.280 81.630 93.610 81.635 ;
        RECT 97.600 81.590 101.810 82.040 ;
        RECT 101.970 81.960 102.280 82.030 ;
        RECT 107.090 81.960 107.430 82.020 ;
        RECT 101.970 81.690 107.430 81.960 ;
        RECT 102.200 81.680 107.430 81.690 ;
        RECT 107.090 81.600 107.430 81.680 ;
        RECT 107.580 81.610 111.270 81.980 ;
        RECT 111.420 81.560 115.630 82.010 ;
        RECT 115.790 81.870 116.100 82.000 ;
        RECT 117.245 81.870 117.395 84.385 ;
        RECT 115.790 81.720 117.395 81.870 ;
        RECT 115.790 81.660 116.100 81.720 ;
        RECT 81.230 80.510 83.060 80.990 ;
        RECT 85.520 80.460 87.350 80.940 ;
        RECT 89.430 80.470 91.270 80.950 ;
        RECT 92.960 80.460 94.780 80.940 ;
        RECT 96.800 80.410 98.630 80.890 ;
        RECT 101.170 80.850 102.960 80.900 ;
        RECT 106.780 80.890 108.540 80.910 ;
        RECT 101.170 80.520 102.970 80.850 ;
        RECT 106.780 80.560 108.550 80.890 ;
        RECT 101.170 80.420 102.960 80.520 ;
        RECT 106.780 80.430 108.540 80.560 ;
        RECT 110.620 80.380 112.430 80.860 ;
        RECT 114.990 80.390 116.760 80.870 ;
        RECT 116.865 79.575 117.015 79.590 ;
        RECT 117.245 79.575 117.395 81.720 ;
        RECT 116.865 79.425 117.395 79.575 ;
        RECT 116.865 78.035 117.015 79.425 ;
        RECT 116.860 78.030 117.015 78.035 ;
        RECT 114.875 77.885 117.015 78.030 ;
        RECT 114.875 73.745 115.025 77.885 ;
        RECT 117.420 73.920 127.540 74.400 ;
        RECT 114.875 73.595 117.090 73.745 ;
        RECT 52.990 71.110 56.670 71.590 ;
        RECT 61.065 70.905 61.315 73.455 ;
        RECT 68.215 73.035 113.985 73.485 ;
        RECT 116.940 73.375 117.090 73.595 ;
        RECT 116.940 73.370 118.500 73.375 ;
        RECT 116.940 73.225 118.655 73.370 ;
        RECT 118.505 73.070 118.655 73.225 ;
        RECT 62.940 71.030 66.160 71.510 ;
        RECT 68.215 70.910 68.665 73.035 ;
        RECT 113.090 72.995 113.985 73.035 ;
        RECT 113.090 72.545 117.905 72.995 ;
        RECT 113.090 72.540 113.680 72.545 ;
        RECT 118.220 72.450 118.660 73.070 ;
        RECT 120.690 72.890 120.990 73.630 ;
        RECT 121.685 73.380 121.975 73.425 ;
        RECT 124.915 73.380 125.205 73.425 ;
        RECT 121.685 73.240 125.205 73.380 ;
        RECT 129.585 73.290 130.315 91.695 ;
        RECT 121.685 73.195 121.975 73.240 ;
        RECT 124.915 73.195 125.205 73.240 ;
        RECT 119.810 72.700 120.100 72.745 ;
        RECT 121.650 72.700 121.940 72.745 ;
        RECT 119.810 72.560 121.940 72.700 ;
        RECT 119.810 72.515 120.100 72.560 ;
        RECT 121.650 72.515 121.940 72.560 ;
        RECT 122.220 72.510 122.550 73.100 ;
        RECT 122.750 72.510 123.020 73.100 ;
        RECT 123.420 72.590 123.850 73.090 ;
        RECT 123.995 72.700 124.285 72.745 ;
        RECT 125.835 72.700 126.125 72.745 ;
        RECT 123.995 72.560 126.125 72.700 ;
        RECT 126.740 72.580 130.315 73.290 ;
        RECT 129.585 72.570 130.315 72.580 ;
        RECT 123.995 72.515 124.285 72.560 ;
        RECT 125.835 72.515 126.125 72.560 ;
        RECT 118.890 72.360 119.180 72.405 ;
        RECT 124.410 72.360 124.700 72.405 ;
        RECT 125.330 72.360 125.620 72.405 ;
        RECT 118.890 72.220 125.620 72.360 ;
        RECT 118.890 72.175 119.180 72.220 ;
        RECT 124.410 72.175 124.700 72.220 ;
        RECT 125.330 72.175 125.620 72.220 ;
        RECT 117.420 71.200 127.540 71.680 ;
        RECT 61.065 70.880 61.320 70.905 ;
        RECT 61.065 70.645 64.700 70.880 ;
        RECT 61.280 70.640 64.700 70.645 ;
        RECT 67.350 70.660 68.665 70.910 ;
        RECT 67.350 70.500 68.660 70.660 ;
        RECT 61.560 70.170 64.900 70.470 ;
        RECT 53.445 69.875 53.835 70.165 ;
        RECT 61.560 70.110 61.930 70.170 ;
        RECT 52.140 69.485 53.835 69.875 ;
        RECT 31.660 66.120 33.090 66.490 ;
        RECT 23.190 65.100 23.740 65.380 ;
        RECT 23.360 64.290 23.515 65.100 ;
        RECT 27.810 65.035 30.405 65.425 ;
        RECT 21.890 63.810 25.570 64.290 ;
        RECT 22.390 62.810 25.140 63.290 ;
        RECT 22.880 61.410 23.260 61.820 ;
        RECT 23.880 61.690 24.130 62.810 ;
        RECT 22.950 60.570 23.210 61.410 ;
        RECT 23.840 61.380 24.180 61.690 ;
        RECT 24.800 61.530 25.550 62.020 ;
        RECT 27.810 60.605 28.200 65.035 ;
        RECT 30.880 64.850 31.290 65.770 ;
        RECT 47.070 65.050 47.370 66.550 ;
        RECT 50.780 66.500 51.210 66.850 ;
        RECT 50.780 66.160 51.040 66.500 ;
        RECT 49.510 65.900 51.040 66.160 ;
        RECT 52.140 65.445 52.530 69.485 ;
        RECT 54.340 69.010 54.690 69.700 ;
        RECT 54.830 69.020 55.170 69.950 ;
        RECT 55.340 69.040 55.700 69.960 ;
        RECT 56.230 69.010 57.660 69.380 ;
        RECT 58.300 69.240 61.050 69.720 ;
        RECT 61.560 69.670 61.920 70.110 ;
        RECT 62.510 69.890 63.040 69.900 ;
        RECT 57.255 68.945 57.660 69.010 ;
        RECT 61.560 68.950 61.910 69.670 ;
        RECT 62.510 69.300 63.360 69.890 ;
        RECT 63.510 69.810 64.210 69.980 ;
        RECT 64.540 69.880 64.900 70.170 ;
        RECT 65.240 70.110 68.660 70.500 ;
        RECT 67.340 69.980 68.660 70.110 ;
        RECT 67.340 69.970 67.520 69.980 ;
        RECT 63.510 69.470 64.200 69.810 ;
        RECT 64.430 69.540 64.900 69.880 ;
        RECT 52.990 68.390 56.670 68.870 ;
        RECT 57.255 68.575 59.645 68.945 ;
        RECT 59.930 68.590 61.910 68.950 ;
        RECT 57.050 67.535 58.795 67.905 ;
        RECT 53.610 66.900 56.370 67.380 ;
        RECT 54.930 66.360 55.420 66.740 ;
        RECT 57.050 66.510 57.420 67.535 ;
        RECT 59.275 67.465 59.645 68.575 ;
        RECT 62.530 68.310 66.160 68.790 ;
        RECT 62.530 68.300 63.000 68.310 ;
        RECT 58.300 66.970 61.050 67.000 ;
        RECT 58.300 66.640 61.100 66.970 ;
        RECT 58.300 66.520 61.050 66.640 ;
        RECT 55.990 66.140 57.420 66.510 ;
        RECT 47.520 65.120 48.070 65.400 ;
        RECT 29.280 64.160 32.040 64.640 ;
        RECT 47.690 64.310 47.845 65.120 ;
        RECT 52.140 65.055 54.735 65.445 ;
        RECT 46.220 63.830 49.900 64.310 ;
        RECT 46.710 62.830 49.470 63.310 ;
        RECT 29.260 61.780 32.020 62.260 ;
        RECT 47.210 61.430 47.590 61.840 ;
        RECT 48.210 61.710 48.460 62.830 ;
        RECT 31.670 60.750 32.010 61.090 ;
        RECT 22.390 60.090 25.140 60.570 ;
        RECT 27.810 60.215 30.475 60.605 ;
        RECT 30.710 60.300 31.060 60.630 ;
        RECT 47.280 60.590 47.540 61.430 ;
        RECT 48.170 61.400 48.510 61.710 ;
        RECT 49.130 61.550 49.880 62.040 ;
        RECT 52.140 60.625 52.530 65.055 ;
        RECT 55.210 64.870 55.620 65.790 ;
        RECT 53.610 64.180 56.370 64.660 ;
        RECT 53.590 62.160 56.350 62.280 ;
        RECT 53.530 61.830 56.350 62.160 ;
        RECT 53.590 61.800 56.350 61.830 ;
        RECT 56.000 60.770 56.340 61.110 ;
        RECT 21.940 58.710 25.620 59.190 ;
        RECT 22.790 57.210 23.090 58.710 ;
        RECT 27.810 58.350 28.200 60.215 ;
        RECT 46.710 60.110 49.470 60.590 ;
        RECT 52.140 60.235 54.805 60.625 ;
        RECT 55.040 60.320 55.390 60.650 ;
        RECT 29.260 59.440 32.020 59.540 ;
        RECT 29.220 59.110 32.020 59.440 ;
        RECT 29.260 59.060 32.020 59.110 ;
        RECT 46.270 58.730 49.950 59.210 ;
        RECT 25.210 57.960 28.200 58.350 ;
        RECT 23.240 57.280 23.790 57.560 ;
        RECT 23.410 56.470 23.565 57.280 ;
        RECT 47.120 57.230 47.420 58.730 ;
        RECT 52.140 58.370 52.530 60.235 ;
        RECT 53.590 59.490 56.350 59.560 ;
        RECT 53.570 59.160 56.350 59.490 ;
        RECT 53.590 59.080 56.350 59.160 ;
        RECT 49.540 57.980 52.530 58.370 ;
        RECT 47.570 57.300 48.120 57.580 ;
        RECT 47.740 56.490 47.895 57.300 ;
        RECT 21.940 55.990 25.620 56.470 ;
        RECT 46.270 56.010 49.950 56.490 ;
        RECT 22.430 54.990 25.190 55.470 ;
        RECT 46.760 55.010 49.520 55.490 ;
        RECT 22.930 53.590 23.310 53.930 ;
        RECT 23.880 53.650 24.240 54.990 ;
        RECT 23.030 52.750 23.280 53.590 ;
        RECT 23.890 53.540 24.230 53.650 ;
        RECT 24.850 53.260 26.010 53.810 ;
        RECT 47.260 53.610 47.640 53.950 ;
        RECT 48.210 53.670 48.570 55.010 ;
        RECT 47.360 52.770 47.610 53.610 ;
        RECT 48.220 53.560 48.560 53.670 ;
        RECT 49.180 53.280 50.340 53.830 ;
        RECT 48.220 52.770 48.560 52.790 ;
        RECT 23.890 52.750 24.230 52.770 ;
        RECT 22.430 52.270 25.190 52.750 ;
        RECT 46.760 52.290 49.520 52.770 ;
        RECT 30.560 33.140 32.350 33.240 ;
        RECT 30.560 32.810 32.420 33.140 ;
        RECT 30.560 32.760 32.350 32.810 ;
        RECT 30.670 31.660 31.140 31.990 ;
        RECT 31.310 31.690 31.640 31.990 ;
        RECT 30.560 30.040 32.350 30.520 ;
        RECT 49.640 29.600 57.450 30.080 ;
        RECT 51.070 28.720 51.360 28.765 ;
        RECT 51.500 28.720 51.640 29.600 ;
        RECT 59.940 29.540 67.760 30.020 ;
        RECT 69.730 29.980 77.550 30.060 ;
        RECT 79.710 30.040 87.520 30.090 ;
        RECT 69.720 29.650 77.550 29.980 ;
        RECT 79.690 29.710 87.520 30.040 ;
        RECT 69.730 29.580 77.550 29.650 ;
        RECT 79.710 29.610 87.520 29.710 ;
        RECT 51.990 29.060 52.280 29.105 ;
        RECT 55.690 29.060 55.980 29.105 ;
        RECT 51.990 28.920 55.980 29.060 ;
        RECT 51.990 28.875 52.280 28.920 ;
        RECT 55.690 28.875 55.980 28.920 ;
        RECT 52.910 28.720 53.200 28.765 ;
        RECT 54.770 28.720 55.060 28.765 ;
        RECT 56.150 28.720 56.440 28.765 ;
        RECT 51.070 28.580 56.440 28.720 ;
        RECT 51.070 28.535 51.360 28.580 ;
        RECT 52.910 28.535 53.200 28.580 ;
        RECT 54.770 28.535 55.060 28.580 ;
        RECT 56.150 28.535 56.440 28.580 ;
        RECT 61.380 28.660 61.670 28.705 ;
        RECT 61.810 28.660 61.950 29.540 ;
        RECT 62.300 29.000 62.590 29.045 ;
        RECT 66.000 29.000 66.290 29.045 ;
        RECT 62.300 28.860 66.290 29.000 ;
        RECT 62.300 28.815 62.590 28.860 ;
        RECT 66.000 28.815 66.290 28.860 ;
        RECT 63.220 28.660 63.510 28.705 ;
        RECT 65.080 28.660 65.370 28.705 ;
        RECT 66.460 28.660 66.750 28.705 ;
        RECT 61.380 28.520 66.750 28.660 ;
        RECT 61.380 28.475 61.670 28.520 ;
        RECT 63.220 28.475 63.510 28.520 ;
        RECT 65.080 28.475 65.370 28.520 ;
        RECT 66.460 28.475 66.750 28.520 ;
        RECT 71.170 28.700 71.460 28.745 ;
        RECT 71.600 28.700 71.740 29.580 ;
        RECT 72.090 29.040 72.380 29.085 ;
        RECT 75.790 29.040 76.080 29.085 ;
        RECT 72.090 28.900 76.080 29.040 ;
        RECT 72.090 28.855 72.380 28.900 ;
        RECT 75.790 28.855 76.080 28.900 ;
        RECT 73.010 28.700 73.300 28.745 ;
        RECT 74.870 28.700 75.160 28.745 ;
        RECT 76.250 28.700 76.540 28.745 ;
        RECT 71.170 28.560 76.540 28.700 ;
        RECT 71.170 28.515 71.460 28.560 ;
        RECT 73.010 28.515 73.300 28.560 ;
        RECT 74.870 28.515 75.160 28.560 ;
        RECT 76.250 28.515 76.540 28.560 ;
        RECT 81.140 28.730 81.430 28.775 ;
        RECT 81.570 28.730 81.710 29.610 ;
        RECT 82.060 29.070 82.350 29.115 ;
        RECT 85.760 29.070 86.050 29.115 ;
        RECT 82.060 28.930 86.050 29.070 ;
        RECT 82.060 28.885 82.350 28.930 ;
        RECT 85.760 28.885 86.050 28.930 ;
        RECT 82.980 28.730 83.270 28.775 ;
        RECT 84.840 28.730 85.130 28.775 ;
        RECT 86.220 28.730 86.510 28.775 ;
        RECT 81.140 28.590 86.510 28.730 ;
        RECT 81.140 28.545 81.430 28.590 ;
        RECT 82.980 28.545 83.270 28.590 ;
        RECT 84.840 28.545 85.130 28.590 ;
        RECT 86.220 28.545 86.510 28.590 ;
        RECT 51.530 28.380 51.820 28.425 ;
        RECT 53.830 28.380 54.120 28.425 ;
        RECT 55.690 28.380 55.980 28.425 ;
        RECT 51.530 28.240 55.980 28.380 ;
        RECT 51.530 28.195 51.820 28.240 ;
        RECT 53.830 28.195 54.120 28.240 ;
        RECT 8.730 27.950 16.540 27.980 ;
        RECT 8.680 27.620 16.540 27.950 ;
        RECT 8.730 27.500 16.540 27.620 ;
        RECT 10.160 26.620 10.450 26.665 ;
        RECT 10.590 26.620 10.730 27.500 ;
        RECT 19.400 27.460 27.210 27.940 ;
        RECT 29.150 27.460 36.970 27.940 ;
        RECT 39.160 27.490 46.980 27.970 ;
        RECT 52.020 27.810 52.350 28.100 ;
        RECT 11.080 26.960 11.370 27.005 ;
        RECT 14.780 26.960 15.070 27.005 ;
        RECT 11.080 26.820 15.070 26.960 ;
        RECT 11.080 26.775 11.370 26.820 ;
        RECT 14.780 26.775 15.070 26.820 ;
        RECT 12.000 26.620 12.290 26.665 ;
        RECT 13.860 26.620 14.150 26.665 ;
        RECT 15.240 26.620 15.530 26.665 ;
        RECT 10.160 26.480 15.530 26.620 ;
        RECT 10.160 26.435 10.450 26.480 ;
        RECT 12.000 26.435 12.290 26.480 ;
        RECT 13.860 26.435 14.150 26.480 ;
        RECT 15.240 26.435 15.530 26.480 ;
        RECT 20.830 26.580 21.120 26.625 ;
        RECT 21.260 26.580 21.400 27.460 ;
        RECT 21.750 26.920 22.040 26.965 ;
        RECT 25.450 26.920 25.740 26.965 ;
        RECT 21.750 26.780 25.740 26.920 ;
        RECT 21.750 26.735 22.040 26.780 ;
        RECT 25.450 26.735 25.740 26.780 ;
        RECT 22.670 26.580 22.960 26.625 ;
        RECT 24.530 26.580 24.820 26.625 ;
        RECT 25.910 26.580 26.200 26.625 ;
        RECT 20.830 26.440 26.200 26.580 ;
        RECT 20.830 26.395 21.120 26.440 ;
        RECT 22.670 26.395 22.960 26.440 ;
        RECT 24.530 26.395 24.820 26.440 ;
        RECT 25.910 26.395 26.200 26.440 ;
        RECT 30.590 26.580 30.880 26.625 ;
        RECT 31.020 26.580 31.160 27.460 ;
        RECT 31.510 26.920 31.800 26.965 ;
        RECT 35.210 26.920 35.500 26.965 ;
        RECT 31.510 26.780 35.500 26.920 ;
        RECT 31.510 26.735 31.800 26.780 ;
        RECT 35.210 26.735 35.500 26.780 ;
        RECT 32.430 26.580 32.720 26.625 ;
        RECT 34.290 26.580 34.580 26.625 ;
        RECT 35.670 26.580 35.960 26.625 ;
        RECT 30.590 26.440 35.960 26.580 ;
        RECT 30.590 26.395 30.880 26.440 ;
        RECT 32.430 26.395 32.720 26.440 ;
        RECT 34.290 26.395 34.580 26.440 ;
        RECT 35.670 26.395 35.960 26.440 ;
        RECT 40.600 26.610 40.890 26.655 ;
        RECT 41.030 26.610 41.170 27.490 ;
        RECT 54.300 27.360 54.440 28.240 ;
        RECT 55.690 28.195 55.980 28.240 ;
        RECT 61.840 28.320 62.130 28.365 ;
        RECT 64.140 28.320 64.430 28.365 ;
        RECT 66.000 28.320 66.290 28.365 ;
        RECT 61.840 28.180 66.290 28.320 ;
        RECT 57.060 28.020 57.360 28.150 ;
        RECT 61.840 28.135 62.130 28.180 ;
        RECT 64.140 28.135 64.430 28.180 ;
        RECT 57.060 27.980 59.090 28.020 ;
        RECT 62.320 27.980 62.620 28.030 ;
        RECT 57.060 27.830 62.620 27.980 ;
        RECT 57.060 27.770 57.360 27.830 ;
        RECT 59.020 27.810 62.620 27.830 ;
        RECT 59.480 27.790 62.620 27.810 ;
        RECT 62.320 27.720 62.620 27.790 ;
        RECT 41.520 26.950 41.810 26.995 ;
        RECT 45.220 26.950 45.510 26.995 ;
        RECT 41.520 26.810 45.510 26.950 ;
        RECT 49.640 26.880 57.450 27.360 ;
        RECT 64.610 27.300 64.750 28.180 ;
        RECT 66.000 28.135 66.290 28.180 ;
        RECT 71.630 28.360 71.920 28.405 ;
        RECT 73.930 28.360 74.220 28.405 ;
        RECT 75.790 28.360 76.080 28.405 ;
        RECT 71.630 28.220 76.080 28.360 ;
        RECT 71.630 28.175 71.920 28.220 ;
        RECT 73.930 28.175 74.220 28.220 ;
        RECT 67.410 27.970 67.670 28.060 ;
        RECT 72.110 28.020 72.410 28.070 ;
        RECT 67.825 27.970 72.410 28.020 ;
        RECT 67.400 27.830 72.410 27.970 ;
        RECT 67.400 27.780 67.940 27.830 ;
        RECT 67.410 27.730 67.670 27.780 ;
        RECT 72.110 27.760 72.410 27.830 ;
        RECT 74.400 27.340 74.540 28.220 ;
        RECT 75.790 28.175 76.080 28.220 ;
        RECT 81.600 28.390 81.890 28.435 ;
        RECT 83.900 28.390 84.190 28.435 ;
        RECT 85.760 28.390 86.050 28.435 ;
        RECT 81.600 28.250 86.050 28.390 ;
        RECT 81.600 28.205 81.890 28.250 ;
        RECT 83.900 28.205 84.190 28.250 ;
        RECT 77.200 28.010 77.460 28.100 ;
        RECT 82.080 28.050 82.380 28.100 ;
        RECT 79.240 28.030 82.380 28.050 ;
        RECT 77.620 28.010 82.380 28.030 ;
        RECT 77.190 27.860 82.380 28.010 ;
        RECT 77.190 27.820 79.420 27.860 ;
        RECT 77.200 27.770 77.460 27.820 ;
        RECT 82.080 27.790 82.380 27.860 ;
        RECT 84.370 27.370 84.510 28.250 ;
        RECT 85.760 28.205 86.050 28.250 ;
        RECT 87.170 28.040 87.430 28.130 ;
        RECT 87.160 27.980 87.700 28.040 ;
        RECT 87.160 27.850 89.110 27.980 ;
        RECT 87.170 27.820 89.110 27.850 ;
        RECT 87.170 27.800 87.570 27.820 ;
        RECT 59.940 26.820 67.760 27.300 ;
        RECT 69.730 26.860 77.550 27.340 ;
        RECT 79.710 26.890 87.520 27.370 ;
        RECT 41.520 26.765 41.810 26.810 ;
        RECT 45.220 26.765 45.510 26.810 ;
        RECT 42.440 26.610 42.730 26.655 ;
        RECT 44.300 26.610 44.590 26.655 ;
        RECT 45.680 26.610 45.970 26.655 ;
        RECT 40.600 26.470 45.970 26.610 ;
        RECT 40.600 26.425 40.890 26.470 ;
        RECT 42.440 26.425 42.730 26.470 ;
        RECT 44.300 26.425 44.590 26.470 ;
        RECT 45.680 26.425 45.970 26.470 ;
        RECT 88.950 26.510 89.110 27.820 ;
        RECT 91.510 27.200 96.110 27.220 ;
        RECT 91.510 26.870 96.130 27.200 ;
        RECT 91.510 26.740 96.110 26.870 ;
        RECT 88.950 26.350 93.660 26.510 ;
        RECT 10.620 26.280 10.910 26.325 ;
        RECT 12.920 26.280 13.210 26.325 ;
        RECT 14.780 26.280 15.070 26.325 ;
        RECT 10.620 26.140 15.070 26.280 ;
        RECT 10.620 26.095 10.910 26.140 ;
        RECT 12.920 26.095 13.210 26.140 ;
        RECT 11.110 25.710 11.440 26.000 ;
        RECT 13.390 25.260 13.530 26.140 ;
        RECT 14.780 26.095 15.070 26.140 ;
        RECT 21.290 26.240 21.580 26.285 ;
        RECT 23.590 26.240 23.880 26.285 ;
        RECT 25.450 26.240 25.740 26.285 ;
        RECT 21.290 26.100 25.740 26.240 ;
        RECT 21.290 26.055 21.580 26.100 ;
        RECT 23.590 26.055 23.880 26.100 ;
        RECT 16.150 25.920 16.450 26.050 ;
        RECT 16.150 25.900 19.185 25.920 ;
        RECT 21.770 25.900 22.070 25.950 ;
        RECT 16.150 25.730 22.070 25.900 ;
        RECT 16.150 25.670 16.450 25.730 ;
        RECT 18.180 25.710 22.070 25.730 ;
        RECT 21.770 25.640 22.070 25.710 ;
        RECT 8.730 24.780 16.540 25.260 ;
        RECT 24.060 25.220 24.200 26.100 ;
        RECT 25.450 26.055 25.740 26.100 ;
        RECT 31.050 26.240 31.340 26.285 ;
        RECT 33.350 26.240 33.640 26.285 ;
        RECT 35.210 26.240 35.500 26.285 ;
        RECT 31.050 26.100 35.500 26.240 ;
        RECT 31.050 26.055 31.340 26.100 ;
        RECT 33.350 26.055 33.640 26.100 ;
        RECT 26.860 25.890 27.120 25.980 ;
        RECT 31.530 25.900 31.830 25.950 ;
        RECT 28.060 25.890 31.830 25.900 ;
        RECT 26.850 25.710 31.830 25.890 ;
        RECT 26.850 25.700 28.295 25.710 ;
        RECT 26.860 25.650 27.120 25.700 ;
        RECT 31.530 25.640 31.830 25.710 ;
        RECT 33.820 25.220 33.960 26.100 ;
        RECT 35.210 26.055 35.500 26.100 ;
        RECT 41.060 26.270 41.350 26.315 ;
        RECT 43.360 26.270 43.650 26.315 ;
        RECT 45.220 26.270 45.510 26.315 ;
        RECT 41.060 26.130 45.510 26.270 ;
        RECT 41.060 26.085 41.350 26.130 ;
        RECT 43.360 26.085 43.650 26.130 ;
        RECT 36.620 25.890 36.880 25.980 ;
        RECT 41.540 25.930 41.840 25.980 ;
        RECT 37.750 25.890 41.840 25.930 ;
        RECT 36.610 25.740 41.840 25.890 ;
        RECT 36.610 25.700 38.055 25.740 ;
        RECT 36.620 25.650 36.880 25.700 ;
        RECT 41.540 25.670 41.840 25.740 ;
        RECT 43.830 25.250 43.970 26.130 ;
        RECT 45.220 26.085 45.510 26.130 ;
        RECT 49.530 26.050 87.620 26.210 ;
        RECT 46.630 25.920 46.890 26.010 ;
        RECT 49.530 25.920 49.690 26.050 ;
        RECT 46.620 25.730 49.690 25.920 ;
        RECT 46.630 25.680 46.890 25.730 ;
        RECT 48.810 25.720 49.690 25.730 ;
        RECT 87.460 25.730 87.620 26.050 ;
        RECT 50.230 25.690 58.050 25.710 ;
        RECT 50.230 25.360 58.070 25.690 ;
        RECT 87.460 25.570 90.890 25.730 ;
        RECT 92.990 25.670 93.240 26.210 ;
        RECT 90.730 25.510 90.890 25.570 ;
        RECT 92.130 25.540 92.400 25.600 ;
        RECT 91.250 25.510 92.860 25.540 ;
        RECT 19.400 24.740 27.210 25.220 ;
        RECT 29.150 24.740 36.970 25.220 ;
        RECT 39.160 24.770 46.980 25.250 ;
        RECT 50.230 25.230 58.050 25.360 ;
        RECT 51.210 24.350 51.500 24.395 ;
        RECT 51.640 24.350 51.780 25.230 ;
        RECT 61.140 25.010 68.940 25.490 ;
        RECT 52.130 24.690 52.420 24.735 ;
        RECT 55.830 24.690 56.120 24.735 ;
        RECT 52.130 24.550 56.120 24.690 ;
        RECT 52.130 24.505 52.420 24.550 ;
        RECT 55.830 24.505 56.120 24.550 ;
        RECT 53.050 24.350 53.340 24.395 ;
        RECT 54.910 24.350 55.200 24.395 ;
        RECT 56.290 24.350 56.580 24.395 ;
        RECT 51.210 24.210 56.580 24.350 ;
        RECT 51.210 24.165 51.500 24.210 ;
        RECT 53.050 24.165 53.340 24.210 ;
        RECT 54.910 24.165 55.200 24.210 ;
        RECT 56.290 24.165 56.580 24.210 ;
        RECT 62.560 24.130 62.850 24.175 ;
        RECT 62.990 24.130 63.130 25.010 ;
        RECT 71.140 24.980 78.950 25.460 ;
        RECT 63.480 24.470 63.770 24.515 ;
        RECT 67.180 24.470 67.470 24.515 ;
        RECT 63.480 24.330 67.470 24.470 ;
        RECT 63.480 24.285 63.770 24.330 ;
        RECT 67.180 24.285 67.470 24.330 ;
        RECT 64.400 24.130 64.690 24.175 ;
        RECT 66.260 24.130 66.550 24.175 ;
        RECT 67.640 24.130 67.930 24.175 ;
        RECT 51.670 24.010 51.960 24.055 ;
        RECT 53.970 24.010 54.260 24.055 ;
        RECT 55.830 24.010 56.120 24.055 ;
        RECT 51.670 23.870 56.120 24.010 ;
        RECT 62.560 23.990 67.930 24.130 ;
        RECT 62.560 23.945 62.850 23.990 ;
        RECT 64.400 23.945 64.690 23.990 ;
        RECT 66.260 23.945 66.550 23.990 ;
        RECT 67.640 23.945 67.930 23.990 ;
        RECT 72.570 24.100 72.860 24.145 ;
        RECT 73.000 24.100 73.140 24.980 ;
        RECT 81.260 24.890 89.060 25.370 ;
        RECT 90.730 25.350 92.860 25.510 ;
        RECT 92.130 25.270 92.400 25.350 ;
        RECT 93.040 25.120 93.200 25.670 ;
        RECT 93.390 25.570 93.660 26.350 ;
        RECT 93.390 25.550 93.580 25.570 ;
        RECT 91.250 25.115 93.200 25.120 ;
        RECT 90.845 24.960 93.200 25.115 ;
        RECT 90.845 24.925 91.385 24.960 ;
        RECT 73.490 24.440 73.780 24.485 ;
        RECT 77.190 24.440 77.480 24.485 ;
        RECT 73.490 24.300 77.480 24.440 ;
        RECT 73.490 24.255 73.780 24.300 ;
        RECT 77.190 24.255 77.480 24.300 ;
        RECT 74.410 24.100 74.700 24.145 ;
        RECT 76.270 24.100 76.560 24.145 ;
        RECT 77.650 24.100 77.940 24.145 ;
        RECT 72.570 23.960 77.940 24.100 ;
        RECT 72.570 23.915 72.860 23.960 ;
        RECT 74.410 23.915 74.700 23.960 ;
        RECT 76.270 23.915 76.560 23.960 ;
        RECT 77.650 23.915 77.940 23.960 ;
        RECT 82.680 24.010 82.970 24.055 ;
        RECT 83.110 24.010 83.250 24.890 ;
        RECT 83.600 24.350 83.890 24.395 ;
        RECT 87.300 24.350 87.590 24.395 ;
        RECT 83.600 24.210 87.590 24.350 ;
        RECT 83.600 24.165 83.890 24.210 ;
        RECT 87.300 24.165 87.590 24.210 ;
        RECT 84.520 24.010 84.810 24.055 ;
        RECT 86.380 24.010 86.670 24.055 ;
        RECT 87.760 24.010 88.050 24.055 ;
        RECT 51.670 23.825 51.960 23.870 ;
        RECT 53.970 23.825 54.260 23.870 ;
        RECT 52.160 23.440 52.490 23.730 ;
        RECT 54.440 22.990 54.580 23.870 ;
        RECT 55.830 23.825 56.120 23.870 ;
        RECT 82.680 23.870 88.050 24.010 ;
        RECT 63.020 23.790 63.310 23.835 ;
        RECT 65.320 23.790 65.610 23.835 ;
        RECT 67.180 23.790 67.470 23.835 ;
        RECT 82.680 23.825 82.970 23.870 ;
        RECT 84.520 23.825 84.810 23.870 ;
        RECT 86.380 23.825 86.670 23.870 ;
        RECT 87.760 23.825 88.050 23.870 ;
        RECT 57.200 23.650 57.500 23.780 ;
        RECT 63.020 23.650 67.470 23.790 ;
        RECT 57.200 23.560 59.090 23.650 ;
        RECT 63.020 23.605 63.310 23.650 ;
        RECT 65.320 23.605 65.610 23.650 ;
        RECT 57.200 23.460 60.510 23.560 ;
        RECT 57.200 23.400 57.500 23.460 ;
        RECT 58.870 23.450 60.510 23.460 ;
        RECT 63.500 23.450 63.800 23.500 ;
        RECT 58.870 23.260 63.800 23.450 ;
        RECT 63.500 23.190 63.800 23.260 ;
        RECT 50.230 22.950 58.050 22.990 ;
        RECT 50.230 22.620 58.060 22.950 ;
        RECT 65.790 22.770 65.930 23.650 ;
        RECT 67.180 23.605 67.470 23.650 ;
        RECT 73.030 23.760 73.320 23.805 ;
        RECT 75.330 23.760 75.620 23.805 ;
        RECT 77.190 23.760 77.480 23.805 ;
        RECT 73.030 23.620 77.480 23.760 ;
        RECT 73.030 23.575 73.320 23.620 ;
        RECT 75.330 23.575 75.620 23.620 ;
        RECT 68.590 23.440 68.850 23.530 ;
        RECT 68.580 23.420 70.525 23.440 ;
        RECT 73.510 23.420 73.810 23.470 ;
        RECT 68.580 23.250 73.810 23.420 ;
        RECT 68.590 23.200 68.850 23.250 ;
        RECT 70.410 23.230 73.810 23.250 ;
        RECT 73.510 23.160 73.810 23.230 ;
        RECT 50.230 22.510 58.050 22.620 ;
        RECT 61.140 22.290 68.940 22.770 ;
        RECT 75.800 22.740 75.940 23.620 ;
        RECT 77.190 23.575 77.480 23.620 ;
        RECT 83.140 23.670 83.430 23.715 ;
        RECT 85.440 23.670 85.730 23.715 ;
        RECT 87.300 23.670 87.590 23.715 ;
        RECT 83.140 23.530 87.590 23.670 ;
        RECT 78.600 23.410 78.860 23.500 ;
        RECT 83.140 23.485 83.430 23.530 ;
        RECT 85.440 23.485 85.730 23.530 ;
        RECT 78.590 23.330 79.350 23.410 ;
        RECT 83.620 23.330 83.920 23.380 ;
        RECT 78.590 23.220 83.920 23.330 ;
        RECT 78.600 23.170 78.860 23.220 ;
        RECT 79.225 23.140 83.920 23.220 ;
        RECT 83.620 23.070 83.920 23.140 ;
        RECT 71.140 22.260 78.950 22.740 ;
        RECT 85.910 22.650 86.050 23.530 ;
        RECT 87.300 23.485 87.590 23.530 ;
        RECT 88.710 23.320 88.970 23.410 ;
        RECT 90.845 23.320 91.035 24.925 ;
        RECT 95.230 24.720 95.560 25.490 ;
        RECT 91.510 24.470 96.110 24.500 ;
        RECT 91.510 24.140 96.130 24.470 ;
        RECT 91.510 24.020 96.110 24.140 ;
        RECT 88.700 23.130 91.035 23.320 ;
        RECT 88.710 23.080 88.970 23.130 ;
        RECT 81.260 22.170 89.060 22.650 ;
        RECT 29.970 16.460 31.790 16.940 ;
        RECT 30.520 15.360 30.990 15.690 ;
        RECT 31.160 15.390 31.490 15.690 ;
        RECT 29.970 13.740 31.790 14.220 ;
        RECT 38.665 11.690 39.495 11.700 ;
        RECT 48.500 11.690 49.415 11.700 ;
        RECT 58.420 11.690 59.135 11.700 ;
        RECT 68.065 11.690 69.145 11.700 ;
        RECT 78.530 11.690 79.675 11.700 ;
        RECT 8.580 11.660 16.390 11.680 ;
        RECT 18.940 11.660 19.805 11.670 ;
        RECT 28.735 11.660 29.375 11.670 ;
        RECT 8.475 11.505 16.390 11.660 ;
        RECT 8.580 11.200 16.390 11.505 ;
        RECT 10.010 10.320 10.300 10.365 ;
        RECT 10.440 10.320 10.580 11.200 ;
        RECT 18.930 11.180 26.740 11.660 ;
        RECT 28.710 11.180 36.500 11.660 ;
        RECT 38.665 11.545 46.510 11.690 ;
        RECT 38.700 11.210 46.510 11.545 ;
        RECT 48.480 11.210 56.270 11.690 ;
        RECT 58.420 11.210 66.230 11.690 ;
        RECT 68.065 11.545 75.990 11.690 ;
        RECT 68.190 11.210 75.990 11.545 ;
        RECT 78.500 11.210 86.310 11.690 ;
        RECT 10.930 10.660 11.220 10.705 ;
        RECT 14.630 10.660 14.920 10.705 ;
        RECT 10.930 10.520 14.920 10.660 ;
        RECT 10.930 10.475 11.220 10.520 ;
        RECT 14.630 10.475 14.920 10.520 ;
        RECT 11.850 10.320 12.140 10.365 ;
        RECT 13.710 10.320 14.000 10.365 ;
        RECT 15.090 10.320 15.380 10.365 ;
        RECT 10.010 10.180 15.380 10.320 ;
        RECT 10.010 10.135 10.300 10.180 ;
        RECT 11.850 10.135 12.140 10.180 ;
        RECT 13.710 10.135 14.000 10.180 ;
        RECT 15.090 10.135 15.380 10.180 ;
        RECT 20.360 10.300 20.650 10.345 ;
        RECT 20.790 10.300 20.930 11.180 ;
        RECT 21.280 10.640 21.570 10.685 ;
        RECT 24.980 10.640 25.270 10.685 ;
        RECT 21.280 10.500 25.270 10.640 ;
        RECT 21.280 10.455 21.570 10.500 ;
        RECT 24.980 10.455 25.270 10.500 ;
        RECT 22.200 10.300 22.490 10.345 ;
        RECT 24.060 10.300 24.350 10.345 ;
        RECT 25.440 10.300 25.730 10.345 ;
        RECT 20.360 10.160 25.730 10.300 ;
        RECT 20.360 10.115 20.650 10.160 ;
        RECT 22.200 10.115 22.490 10.160 ;
        RECT 24.060 10.115 24.350 10.160 ;
        RECT 25.440 10.115 25.730 10.160 ;
        RECT 30.120 10.300 30.410 10.345 ;
        RECT 30.550 10.300 30.690 11.180 ;
        RECT 31.040 10.640 31.330 10.685 ;
        RECT 34.740 10.640 35.030 10.685 ;
        RECT 31.040 10.500 35.030 10.640 ;
        RECT 31.040 10.455 31.330 10.500 ;
        RECT 34.740 10.455 35.030 10.500 ;
        RECT 31.960 10.300 32.250 10.345 ;
        RECT 33.820 10.300 34.110 10.345 ;
        RECT 35.200 10.300 35.490 10.345 ;
        RECT 30.120 10.160 35.490 10.300 ;
        RECT 30.120 10.115 30.410 10.160 ;
        RECT 31.960 10.115 32.250 10.160 ;
        RECT 33.820 10.115 34.110 10.160 ;
        RECT 35.200 10.115 35.490 10.160 ;
        RECT 40.130 10.330 40.420 10.375 ;
        RECT 40.560 10.330 40.700 11.210 ;
        RECT 41.050 10.670 41.340 10.715 ;
        RECT 44.750 10.670 45.040 10.715 ;
        RECT 41.050 10.530 45.040 10.670 ;
        RECT 41.050 10.485 41.340 10.530 ;
        RECT 44.750 10.485 45.040 10.530 ;
        RECT 41.970 10.330 42.260 10.375 ;
        RECT 43.830 10.330 44.120 10.375 ;
        RECT 45.210 10.330 45.500 10.375 ;
        RECT 40.130 10.190 45.500 10.330 ;
        RECT 40.130 10.145 40.420 10.190 ;
        RECT 41.970 10.145 42.260 10.190 ;
        RECT 43.830 10.145 44.120 10.190 ;
        RECT 45.210 10.145 45.500 10.190 ;
        RECT 49.890 10.330 50.180 10.375 ;
        RECT 50.320 10.330 50.460 11.210 ;
        RECT 50.810 10.670 51.100 10.715 ;
        RECT 54.510 10.670 54.800 10.715 ;
        RECT 50.810 10.530 54.800 10.670 ;
        RECT 50.810 10.485 51.100 10.530 ;
        RECT 54.510 10.485 54.800 10.530 ;
        RECT 51.730 10.330 52.020 10.375 ;
        RECT 53.590 10.330 53.880 10.375 ;
        RECT 54.970 10.330 55.260 10.375 ;
        RECT 49.890 10.190 55.260 10.330 ;
        RECT 49.890 10.145 50.180 10.190 ;
        RECT 51.730 10.145 52.020 10.190 ;
        RECT 53.590 10.145 53.880 10.190 ;
        RECT 54.970 10.145 55.260 10.190 ;
        RECT 59.850 10.330 60.140 10.375 ;
        RECT 60.280 10.330 60.420 11.210 ;
        RECT 60.770 10.670 61.060 10.715 ;
        RECT 64.470 10.670 64.760 10.715 ;
        RECT 60.770 10.530 64.760 10.670 ;
        RECT 60.770 10.485 61.060 10.530 ;
        RECT 64.470 10.485 64.760 10.530 ;
        RECT 61.690 10.330 61.980 10.375 ;
        RECT 63.550 10.330 63.840 10.375 ;
        RECT 64.930 10.330 65.220 10.375 ;
        RECT 59.850 10.190 65.220 10.330 ;
        RECT 59.850 10.145 60.140 10.190 ;
        RECT 61.690 10.145 61.980 10.190 ;
        RECT 63.550 10.145 63.840 10.190 ;
        RECT 64.930 10.145 65.220 10.190 ;
        RECT 69.610 10.330 69.900 10.375 ;
        RECT 70.040 10.330 70.180 11.210 ;
        RECT 70.530 10.670 70.820 10.715 ;
        RECT 74.230 10.670 74.520 10.715 ;
        RECT 70.530 10.530 74.520 10.670 ;
        RECT 70.530 10.485 70.820 10.530 ;
        RECT 74.230 10.485 74.520 10.530 ;
        RECT 71.450 10.330 71.740 10.375 ;
        RECT 73.310 10.330 73.600 10.375 ;
        RECT 74.690 10.330 74.980 10.375 ;
        RECT 69.610 10.190 74.980 10.330 ;
        RECT 69.610 10.145 69.900 10.190 ;
        RECT 71.450 10.145 71.740 10.190 ;
        RECT 73.310 10.145 73.600 10.190 ;
        RECT 74.690 10.145 74.980 10.190 ;
        RECT 79.930 10.330 80.220 10.375 ;
        RECT 80.360 10.330 80.500 11.210 ;
        RECT 80.850 10.670 81.140 10.715 ;
        RECT 84.550 10.670 84.840 10.715 ;
        RECT 80.850 10.530 84.840 10.670 ;
        RECT 80.850 10.485 81.140 10.530 ;
        RECT 84.550 10.485 84.840 10.530 ;
        RECT 81.770 10.330 82.060 10.375 ;
        RECT 83.630 10.330 83.920 10.375 ;
        RECT 85.010 10.330 85.300 10.375 ;
        RECT 79.930 10.190 85.300 10.330 ;
        RECT 79.930 10.145 80.220 10.190 ;
        RECT 81.770 10.145 82.060 10.190 ;
        RECT 83.630 10.145 83.920 10.190 ;
        RECT 85.010 10.145 85.300 10.190 ;
        RECT 10.470 9.980 10.760 10.025 ;
        RECT 12.770 9.980 13.060 10.025 ;
        RECT 14.630 9.980 14.920 10.025 ;
        RECT 10.470 9.840 14.920 9.980 ;
        RECT 10.470 9.795 10.760 9.840 ;
        RECT 12.770 9.795 13.060 9.840 ;
        RECT 10.960 9.410 11.290 9.700 ;
        RECT 13.240 8.960 13.380 9.840 ;
        RECT 14.630 9.795 14.920 9.840 ;
        RECT 20.820 9.960 21.110 10.005 ;
        RECT 23.120 9.960 23.410 10.005 ;
        RECT 24.980 9.960 25.270 10.005 ;
        RECT 20.820 9.820 25.270 9.960 ;
        RECT 20.820 9.775 21.110 9.820 ;
        RECT 23.120 9.775 23.410 9.820 ;
        RECT 16.000 9.620 16.300 9.750 ;
        RECT 21.300 9.620 21.600 9.670 ;
        RECT 16.000 9.430 21.600 9.620 ;
        RECT 16.000 9.370 16.300 9.430 ;
        RECT 21.300 9.360 21.600 9.430 ;
        RECT 8.580 8.480 16.390 8.960 ;
        RECT 23.590 8.940 23.730 9.820 ;
        RECT 24.980 9.775 25.270 9.820 ;
        RECT 30.580 9.960 30.870 10.005 ;
        RECT 32.880 9.960 33.170 10.005 ;
        RECT 34.740 9.960 35.030 10.005 ;
        RECT 30.580 9.820 35.030 9.960 ;
        RECT 30.580 9.775 30.870 9.820 ;
        RECT 32.880 9.775 33.170 9.820 ;
        RECT 26.390 9.610 26.650 9.700 ;
        RECT 31.060 9.620 31.360 9.670 ;
        RECT 27.590 9.610 31.360 9.620 ;
        RECT 26.380 9.430 31.360 9.610 ;
        RECT 26.380 9.420 27.825 9.430 ;
        RECT 26.390 9.370 26.650 9.420 ;
        RECT 31.060 9.360 31.360 9.430 ;
        RECT 33.350 8.940 33.490 9.820 ;
        RECT 34.740 9.775 35.030 9.820 ;
        RECT 40.590 9.990 40.880 10.035 ;
        RECT 42.890 9.990 43.180 10.035 ;
        RECT 44.750 9.990 45.040 10.035 ;
        RECT 40.590 9.850 45.040 9.990 ;
        RECT 40.590 9.805 40.880 9.850 ;
        RECT 42.890 9.805 43.180 9.850 ;
        RECT 36.150 9.610 36.410 9.700 ;
        RECT 41.070 9.650 41.370 9.700 ;
        RECT 37.280 9.610 41.370 9.650 ;
        RECT 36.140 9.460 41.370 9.610 ;
        RECT 36.140 9.420 37.585 9.460 ;
        RECT 36.150 9.370 36.410 9.420 ;
        RECT 41.070 9.390 41.370 9.460 ;
        RECT 43.360 8.970 43.500 9.850 ;
        RECT 44.750 9.805 45.040 9.850 ;
        RECT 50.350 9.990 50.640 10.035 ;
        RECT 52.650 9.990 52.940 10.035 ;
        RECT 54.510 9.990 54.800 10.035 ;
        RECT 50.350 9.850 54.800 9.990 ;
        RECT 50.350 9.805 50.640 9.850 ;
        RECT 52.650 9.805 52.940 9.850 ;
        RECT 46.160 9.640 46.420 9.730 ;
        RECT 50.830 9.650 51.130 9.700 ;
        RECT 47.360 9.640 51.130 9.650 ;
        RECT 46.150 9.460 51.130 9.640 ;
        RECT 46.150 9.450 47.595 9.460 ;
        RECT 46.160 9.400 46.420 9.450 ;
        RECT 50.830 9.390 51.130 9.460 ;
        RECT 53.120 8.970 53.260 9.850 ;
        RECT 54.510 9.805 54.800 9.850 ;
        RECT 60.310 9.990 60.600 10.035 ;
        RECT 62.610 9.990 62.900 10.035 ;
        RECT 64.470 9.990 64.760 10.035 ;
        RECT 60.310 9.850 64.760 9.990 ;
        RECT 60.310 9.805 60.600 9.850 ;
        RECT 62.610 9.805 62.900 9.850 ;
        RECT 55.920 9.640 56.180 9.730 ;
        RECT 60.790 9.650 61.090 9.700 ;
        RECT 56.585 9.640 61.090 9.650 ;
        RECT 55.910 9.460 61.090 9.640 ;
        RECT 55.910 9.450 56.910 9.460 ;
        RECT 55.920 9.400 56.180 9.450 ;
        RECT 60.790 9.390 61.090 9.460 ;
        RECT 63.080 8.970 63.220 9.850 ;
        RECT 64.470 9.805 64.760 9.850 ;
        RECT 70.070 9.990 70.360 10.035 ;
        RECT 72.370 9.990 72.660 10.035 ;
        RECT 74.230 9.990 74.520 10.035 ;
        RECT 70.070 9.850 74.520 9.990 ;
        RECT 70.070 9.805 70.360 9.850 ;
        RECT 72.370 9.805 72.660 9.850 ;
        RECT 65.880 9.640 66.140 9.730 ;
        RECT 70.550 9.650 70.850 9.700 ;
        RECT 67.080 9.640 70.850 9.650 ;
        RECT 65.870 9.460 70.850 9.640 ;
        RECT 65.870 9.450 67.315 9.460 ;
        RECT 65.880 9.400 66.140 9.450 ;
        RECT 70.550 9.390 70.850 9.460 ;
        RECT 72.840 8.970 72.980 9.850 ;
        RECT 74.230 9.805 74.520 9.850 ;
        RECT 80.390 9.990 80.680 10.035 ;
        RECT 82.690 9.990 82.980 10.035 ;
        RECT 84.550 9.990 84.840 10.035 ;
        RECT 80.390 9.850 84.840 9.990 ;
        RECT 80.390 9.805 80.680 9.850 ;
        RECT 82.690 9.805 82.980 9.850 ;
        RECT 75.640 9.640 75.900 9.730 ;
        RECT 80.870 9.650 81.170 9.700 ;
        RECT 77.690 9.640 81.170 9.650 ;
        RECT 75.630 9.460 81.170 9.640 ;
        RECT 75.630 9.450 77.875 9.460 ;
        RECT 75.640 9.400 75.900 9.450 ;
        RECT 80.870 9.390 81.170 9.460 ;
        RECT 83.160 8.970 83.300 9.850 ;
        RECT 84.550 9.805 84.840 9.850 ;
        RECT 85.960 9.640 86.220 9.730 ;
        RECT 86.810 9.640 87.440 9.910 ;
        RECT 85.950 9.450 87.440 9.640 ;
        RECT 85.960 9.400 86.220 9.450 ;
        RECT 86.810 9.140 87.440 9.450 ;
        RECT 18.930 8.625 26.740 8.940 ;
        RECT 28.710 8.625 36.500 8.940 ;
        RECT 8.595 8.460 9.245 8.480 ;
        RECT 18.915 8.470 26.740 8.625 ;
        RECT 28.690 8.470 36.500 8.625 ;
        RECT 38.700 8.490 46.510 8.970 ;
        RECT 48.480 8.490 56.270 8.970 ;
        RECT 58.420 8.490 66.230 8.970 ;
        RECT 68.190 8.490 75.990 8.970 ;
        RECT 78.500 8.655 86.310 8.970 ;
        RECT 78.405 8.500 86.310 8.655 ;
        RECT 78.500 8.490 86.310 8.500 ;
        RECT 18.930 8.460 26.740 8.470 ;
        RECT 28.710 8.460 36.500 8.470 ;
      LAYER met2 ;
        RECT 92.950 219.140 95.640 220.840 ;
        RECT 92.770 212.880 93.220 215.010 ;
        RECT 95.590 212.650 96.040 214.780 ;
        RECT 92.650 203.460 93.100 205.590 ;
        RECT 95.450 203.350 95.900 205.480 ;
        RECT 92.740 195.430 93.190 197.560 ;
        RECT 95.460 195.290 95.910 197.420 ;
        RECT 92.790 189.360 93.240 191.490 ;
        RECT 95.530 189.470 95.980 191.600 ;
        RECT 92.840 184.070 93.290 186.200 ;
        RECT 95.570 184.020 96.020 186.150 ;
        RECT 92.870 180.890 93.350 181.360 ;
        RECT 95.600 180.900 96.090 181.600 ;
        RECT 91.700 171.100 92.560 173.240 ;
        RECT 94.800 171.020 95.580 173.130 ;
        RECT 91.740 159.570 92.600 161.710 ;
        RECT 94.840 159.490 95.620 161.600 ;
        RECT 91.780 148.500 92.640 150.640 ;
        RECT 94.880 148.420 95.660 150.530 ;
        RECT 91.690 137.500 92.550 139.640 ;
        RECT 94.790 137.420 95.570 139.530 ;
        RECT 91.730 126.430 92.590 128.570 ;
        RECT 94.830 126.350 95.610 128.460 ;
        RECT 41.900 116.710 44.040 117.570 ;
        RECT 52.970 116.750 55.110 117.610 ;
        RECT 63.970 116.660 66.110 117.520 ;
        RECT 75.040 116.700 77.180 117.560 ;
        RECT 86.570 116.740 88.710 117.600 ;
        RECT 41.820 113.690 43.930 114.470 ;
        RECT 52.890 113.730 55.000 114.510 ;
        RECT 63.890 113.640 66.000 114.420 ;
        RECT 74.960 113.680 77.070 114.460 ;
        RECT 86.490 113.720 88.600 114.500 ;
        RECT 47.150 88.730 48.530 89.220 ;
        RECT 78.045 88.000 79.105 88.460 ;
        RECT 81.955 88.200 83.015 88.660 ;
        RECT 86.305 88.200 87.365 88.660 ;
        RECT 90.255 88.160 91.315 88.620 ;
        RECT 95.775 88.170 96.835 88.630 ;
        RECT 100.125 88.170 101.185 88.630 ;
        RECT 104.075 88.130 105.135 88.590 ;
        RECT 107.055 88.120 108.115 88.580 ;
        RECT 111.405 88.120 112.465 88.580 ;
        RECT 115.355 88.080 116.415 88.540 ;
        RECT 32.315 87.935 32.725 87.940 ;
        RECT 32.315 87.930 33.795 87.935 ;
        RECT 32.315 87.525 33.800 87.930 ;
        RECT 22.360 82.680 23.660 83.180 ;
        RECT 29.730 81.560 30.740 82.190 ;
        RECT 24.430 79.970 25.530 80.450 ;
        RECT 22.810 78.960 24.690 79.400 ;
        RECT 24.790 77.360 25.330 77.550 ;
        RECT 24.790 77.180 27.290 77.360 ;
        RECT 24.180 76.270 25.140 76.750 ;
        RECT 22.380 74.890 23.750 75.350 ;
        RECT 24.730 72.170 25.590 72.620 ;
        RECT 22.880 71.160 24.350 71.600 ;
        RECT 27.110 70.490 27.290 77.180 ;
        RECT 28.740 73.200 29.540 73.680 ;
        RECT 30.050 72.550 30.390 81.560 ;
        RECT 32.315 77.120 32.725 87.525 ;
        RECT 33.020 87.490 33.800 87.525 ;
        RECT 47.160 86.010 48.530 86.510 ;
        RECT 57.005 85.270 57.415 85.275 ;
        RECT 78.095 85.270 79.155 85.730 ;
        RECT 81.895 85.470 82.955 85.930 ;
        RECT 86.355 85.470 87.415 85.930 ;
        RECT 90.205 85.440 91.265 85.900 ;
        RECT 95.715 85.440 96.775 85.900 ;
        RECT 100.175 85.440 101.235 85.900 ;
        RECT 104.025 85.410 105.085 85.870 ;
        RECT 106.995 85.390 108.055 85.850 ;
        RECT 111.455 85.390 112.515 85.850 ;
        RECT 115.305 85.360 116.365 85.820 ;
        RECT 57.000 85.165 57.530 85.270 ;
        RECT 57.000 84.060 57.535 85.165 ;
        RECT 56.645 83.650 57.535 84.060 ;
        RECT 46.690 82.700 47.990 83.200 ;
        RECT 54.060 81.580 55.070 82.210 ;
        RECT 48.760 79.990 49.860 80.470 ;
        RECT 47.140 78.980 49.020 79.420 ;
        RECT 33.040 78.420 34.470 78.900 ;
        RECT 49.120 77.380 49.660 77.570 ;
        RECT 49.120 77.200 51.620 77.380 ;
        RECT 32.315 76.710 33.410 77.120 ;
        RECT 30.540 75.920 31.270 76.400 ;
        RECT 48.510 76.290 49.470 76.770 ;
        RECT 35.230 75.700 36.260 76.190 ;
        RECT 46.710 74.910 48.080 75.370 ;
        RECT 30.050 72.210 30.840 72.550 ;
        RECT 27.110 70.310 30.160 70.490 ;
        RECT 29.980 69.680 30.160 70.310 ;
        RECT 24.840 69.400 25.690 69.560 ;
        RECT 29.980 69.400 30.360 69.680 ;
        RECT 24.840 69.160 28.570 69.400 ;
        RECT 29.970 69.160 30.360 69.400 ;
        RECT 24.840 69.090 25.690 69.160 ;
        RECT 24.100 68.420 25.200 68.900 ;
        RECT 28.320 67.960 28.560 69.160 ;
        RECT 30.010 68.970 30.360 69.160 ;
        RECT 30.500 68.960 30.840 72.210 ;
        RECT 38.175 72.435 42.655 72.905 ;
        RECT 31.610 71.090 32.350 71.580 ;
        RECT 31.005 69.005 31.375 69.925 ;
        RECT 38.175 69.870 38.645 72.435 ;
        RECT 39.200 71.020 40.360 71.480 ;
        RECT 33.970 69.210 34.730 69.690 ;
        RECT 38.175 69.285 39.030 69.870 ;
        RECT 39.190 69.450 39.880 69.960 ;
        RECT 38.620 69.280 39.030 69.285 ;
        RECT 29.120 68.360 29.870 68.850 ;
        RECT 31.005 68.635 31.715 69.005 ;
        RECT 28.320 67.720 30.870 67.960 ;
        RECT 22.340 66.550 23.690 66.980 ;
        RECT 29.750 66.890 30.420 67.350 ;
        RECT 30.630 66.860 30.870 67.720 ;
        RECT 26.800 66.830 28.830 66.840 ;
        RECT 26.450 66.480 28.830 66.830 ;
        RECT 28.470 65.850 28.830 66.480 ;
        RECT 30.600 66.340 31.090 66.860 ;
        RECT 31.345 65.860 31.715 68.635 ;
        RECT 38.210 68.290 38.720 68.770 ;
        RECT 39.290 68.280 39.630 69.450 ;
        RECT 39.190 68.270 39.630 68.280 ;
        RECT 38.890 67.930 39.630 68.270 ;
        RECT 35.480 66.500 36.240 66.980 ;
        RECT 30.700 65.850 31.715 65.860 ;
        RECT 28.470 65.490 31.715 65.850 ;
        RECT 30.930 64.720 31.290 65.490 ;
        RECT 24.610 63.830 25.560 64.270 ;
        RECT 29.740 64.170 30.500 64.640 ;
        RECT 22.870 62.800 23.900 63.270 ;
        RECT 24.800 61.690 25.550 62.020 ;
        RECT 31.150 61.780 32.010 62.260 ;
        RECT 24.800 61.530 30.950 61.690 ;
        RECT 30.790 60.630 30.950 61.530 ;
        RECT 38.890 61.090 39.230 67.930 ;
        RECT 31.670 60.750 39.230 61.090 ;
        RECT 24.290 60.110 25.120 60.580 ;
        RECT 30.710 60.300 31.060 60.630 ;
        RECT 22.550 58.730 23.450 59.170 ;
        RECT 29.720 59.060 30.500 59.540 ;
        RECT 24.690 56.020 25.590 56.460 ;
        RECT 22.900 54.980 23.880 55.460 ;
        RECT 42.185 53.810 42.655 72.435 ;
        RECT 49.060 72.190 49.920 72.640 ;
        RECT 47.210 71.180 48.680 71.620 ;
        RECT 51.440 70.510 51.620 77.200 ;
        RECT 53.070 73.220 53.870 73.700 ;
        RECT 54.380 72.570 54.720 81.580 ;
        RECT 56.645 77.140 57.055 83.650 ;
        RECT 81.730 83.230 82.790 83.690 ;
        RECT 85.580 83.200 86.640 83.660 ;
        RECT 90.040 83.200 91.100 83.660 ;
        RECT 93.010 83.180 94.070 83.640 ;
        RECT 96.860 83.150 97.920 83.610 ;
        RECT 101.320 83.150 102.380 83.610 ;
        RECT 106.830 83.150 107.890 83.610 ;
        RECT 110.680 83.120 111.740 83.580 ;
        RECT 115.140 83.120 116.200 83.580 ;
        RECT 81.680 80.510 82.740 80.970 ;
        RECT 85.630 80.470 86.690 80.930 ;
        RECT 89.980 80.470 91.040 80.930 ;
        RECT 92.960 80.460 94.020 80.920 ;
        RECT 96.910 80.420 97.970 80.880 ;
        RECT 101.260 80.420 102.320 80.880 ;
        RECT 106.780 80.430 107.840 80.890 ;
        RECT 110.730 80.390 111.790 80.850 ;
        RECT 115.080 80.390 116.140 80.850 ;
        RECT 57.370 78.440 58.800 78.920 ;
        RECT 56.645 76.730 57.740 77.140 ;
        RECT 54.870 75.940 55.600 76.420 ;
        RECT 59.560 75.720 60.590 76.210 ;
        RECT 121.560 73.940 122.710 74.400 ;
        RECT 131.945 74.215 137.320 74.605 ;
        RECT 131.945 73.700 132.335 74.215 ;
        RECT 131.945 73.630 132.330 73.700 ;
        RECT 120.690 73.290 132.330 73.630 ;
        RECT 54.380 72.230 55.170 72.570 ;
        RECT 51.440 70.330 54.490 70.510 ;
        RECT 54.310 69.700 54.490 70.330 ;
        RECT 49.170 69.420 50.020 69.580 ;
        RECT 54.310 69.420 54.690 69.700 ;
        RECT 49.170 69.180 52.900 69.420 ;
        RECT 54.300 69.180 54.690 69.420 ;
        RECT 49.170 69.110 50.020 69.180 ;
        RECT 48.430 68.440 49.530 68.920 ;
        RECT 52.650 67.980 52.890 69.180 ;
        RECT 54.340 68.990 54.690 69.180 ;
        RECT 54.830 68.980 55.170 72.230 ;
        RECT 62.505 72.455 66.985 72.925 ;
        RECT 120.690 72.890 120.990 73.290 ;
        RECT 131.945 73.285 132.330 73.290 ;
        RECT 134.740 73.630 135.860 73.970 ;
        RECT 134.740 73.290 135.880 73.630 ;
        RECT 55.940 71.110 56.680 71.600 ;
        RECT 55.335 69.025 55.705 69.945 ;
        RECT 62.505 69.890 62.975 72.455 ;
        RECT 63.530 71.040 64.690 71.500 ;
        RECT 58.300 69.230 59.060 69.710 ;
        RECT 62.505 69.305 63.360 69.890 ;
        RECT 63.520 69.470 64.210 69.980 ;
        RECT 62.950 69.300 63.360 69.305 ;
        RECT 53.450 68.380 54.200 68.870 ;
        RECT 55.335 68.655 56.045 69.025 ;
        RECT 52.650 67.740 55.200 67.980 ;
        RECT 46.670 66.570 48.020 67.000 ;
        RECT 54.080 66.910 54.750 67.370 ;
        RECT 54.960 66.880 55.200 67.740 ;
        RECT 51.130 66.850 53.160 66.860 ;
        RECT 50.780 66.500 53.160 66.850 ;
        RECT 52.800 65.870 53.160 66.500 ;
        RECT 54.930 66.360 55.420 66.880 ;
        RECT 55.675 65.880 56.045 68.655 ;
        RECT 62.540 68.310 63.050 68.790 ;
        RECT 63.620 68.300 63.960 69.470 ;
        RECT 63.520 68.290 63.960 68.300 ;
        RECT 63.220 67.950 63.960 68.290 ;
        RECT 59.810 66.520 60.570 67.000 ;
        RECT 55.030 65.870 56.045 65.880 ;
        RECT 52.800 65.510 56.045 65.870 ;
        RECT 55.260 64.740 55.620 65.510 ;
        RECT 48.940 63.850 49.890 64.290 ;
        RECT 54.070 64.190 54.830 64.660 ;
        RECT 47.200 62.820 48.230 63.290 ;
        RECT 49.130 61.710 49.880 62.040 ;
        RECT 55.480 61.800 56.340 62.280 ;
        RECT 49.130 61.550 55.280 61.710 ;
        RECT 55.120 60.650 55.280 61.550 ;
        RECT 63.220 61.110 63.560 67.950 ;
        RECT 56.000 60.770 63.560 61.110 ;
        RECT 48.620 60.130 49.450 60.600 ;
        RECT 55.040 60.320 55.390 60.650 ;
        RECT 46.880 58.750 47.780 59.190 ;
        RECT 54.050 59.080 54.830 59.560 ;
        RECT 49.020 56.040 49.920 56.480 ;
        RECT 47.230 55.000 48.210 55.480 ;
        RECT 66.515 53.830 66.985 72.455 ;
        RECT 119.250 71.200 121.060 71.670 ;
        RECT 122.240 70.560 122.520 73.100 ;
        RECT 122.240 70.280 122.510 70.560 ;
        RECT 24.850 53.340 42.655 53.810 ;
        RECT 49.180 53.360 66.985 53.830 ;
        RECT 116.290 70.000 122.510 70.280 ;
        RECT 24.850 53.260 26.010 53.340 ;
        RECT 49.180 53.280 50.340 53.360 ;
        RECT 24.280 52.290 25.180 52.730 ;
        RECT 48.610 52.310 49.510 52.750 ;
        RECT 30.560 32.790 31.940 33.240 ;
        RECT 27.925 31.990 28.255 32.020 ;
        RECT 11.110 31.660 31.140 31.990 ;
        RECT 31.310 31.970 65.780 31.990 ;
        RECT 116.290 31.970 116.570 70.000 ;
        RECT 122.730 66.450 123.030 73.110 ;
        RECT 123.425 72.705 124.350 73.095 ;
        RECT 134.740 73.020 135.860 73.290 ;
        RECT 123.425 72.495 123.815 72.705 ;
        RECT 123.960 72.570 124.350 72.705 ;
        RECT 134.965 72.570 135.355 73.020 ;
        RECT 123.960 72.180 135.355 72.570 ;
        RECT 136.930 72.570 137.320 74.215 ;
        RECT 136.930 72.550 138.020 72.570 ;
        RECT 136.930 72.180 138.650 72.550 ;
        RECT 137.560 71.680 138.650 72.180 ;
        RECT 31.310 31.700 116.570 31.970 ;
        RECT 31.310 31.690 80.250 31.700 ;
        RECT 85.750 31.690 116.570 31.700 ;
        RECT 121.260 66.150 123.040 66.450 ;
        RECT 93.965 31.680 94.240 31.690 ;
        RECT 11.110 25.710 11.450 31.660 ;
        RECT 30.550 30.090 31.370 30.520 ;
        RECT 12.550 27.510 13.450 27.980 ;
        RECT 23.140 27.460 24.040 27.930 ;
        RECT 32.900 27.460 33.800 27.930 ;
        RECT 42.910 27.490 43.810 27.960 ;
        RECT 52.020 27.810 52.360 30.090 ;
        RECT 53.540 29.610 54.440 30.080 ;
        RECT 63.690 29.540 64.590 30.010 ;
        RECT 73.480 29.580 74.380 30.050 ;
        RECT 83.450 29.610 84.350 30.080 ;
        RECT 55.710 26.890 56.620 27.370 ;
        RECT 63.690 26.820 64.590 27.290 ;
        RECT 73.480 26.860 74.380 27.330 ;
        RECT 83.450 26.890 84.350 27.360 ;
        RECT 93.290 26.740 94.190 27.220 ;
        RECT 95.965 25.875 96.240 31.690 ;
        RECT 12.600 24.780 13.500 25.250 ;
        RECT 23.140 24.740 24.040 25.210 ;
        RECT 32.900 24.740 33.800 25.210 ;
        RECT 42.910 24.770 43.810 25.240 ;
        RECT 50.640 25.230 51.540 25.710 ;
        RECT 95.980 25.490 96.220 25.875 ;
        RECT 64.870 25.010 65.770 25.480 ;
        RECT 74.880 24.980 75.780 25.450 ;
        RECT 84.990 24.890 85.890 25.360 ;
        RECT 95.240 25.250 96.220 25.490 ;
        RECT 95.240 24.710 95.560 25.250 ;
        RECT 52.160 22.510 52.500 24.010 ;
        RECT 93.310 23.990 94.210 24.470 ;
        RECT 53.670 22.490 54.570 22.970 ;
        RECT 64.870 22.290 65.770 22.760 ;
        RECT 74.880 22.260 75.780 22.730 ;
        RECT 84.990 22.170 85.890 22.640 ;
        RECT 30.410 16.460 31.770 16.930 ;
        RECT 121.260 15.690 121.560 66.150 ;
        RECT 10.960 15.360 30.990 15.690 ;
        RECT 31.160 15.390 121.560 15.690 ;
        RECT 10.960 9.410 11.300 15.360 ;
        RECT 30.400 13.760 31.500 14.210 ;
        RECT 12.700 11.210 13.600 11.680 ;
        RECT 22.670 11.180 23.570 11.650 ;
        RECT 32.430 11.180 33.330 11.650 ;
        RECT 42.440 11.210 43.340 11.680 ;
        RECT 52.200 11.210 53.100 11.680 ;
        RECT 62.160 11.210 63.060 11.680 ;
        RECT 71.920 11.210 72.820 11.680 ;
        RECT 82.240 11.210 83.140 11.680 ;
        RECT 86.950 9.910 87.250 15.390 ;
        RECT 86.810 9.140 87.440 9.910 ;
        RECT 12.690 8.500 13.590 8.970 ;
        RECT 22.670 8.460 23.570 8.930 ;
        RECT 32.430 8.460 33.330 8.930 ;
        RECT 42.440 8.490 43.340 8.960 ;
        RECT 52.200 8.490 53.100 8.960 ;
        RECT 62.160 8.490 63.060 8.960 ;
        RECT 71.920 8.490 72.820 8.960 ;
        RECT 82.240 8.490 83.140 8.960 ;
      LAYER met3 ;
        RECT 92.950 219.140 95.640 220.840 ;
        RECT 88.260 215.010 90.380 217.030 ;
        RECT 88.260 212.890 93.360 215.010 ;
        RECT 97.240 214.780 99.400 218.110 ;
        RECT 88.260 205.550 90.380 212.890 ;
        RECT 95.510 212.620 99.400 214.780 ;
        RECT 92.650 205.550 93.100 205.590 ;
        RECT 88.260 203.430 93.180 205.550 ;
        RECT 97.240 205.510 99.400 212.620 ;
        RECT 95.580 205.480 99.400 205.510 ;
        RECT 88.260 197.540 90.380 203.430 ;
        RECT 95.450 203.350 99.400 205.480 ;
        RECT 88.260 195.420 93.180 197.540 ;
        RECT 97.240 197.430 99.400 203.350 ;
        RECT 95.580 197.420 99.400 197.430 ;
        RECT 88.260 191.430 90.380 195.420 ;
        RECT 95.460 195.290 99.400 197.420 ;
        RECT 95.580 195.270 99.400 195.290 ;
        RECT 97.240 191.550 99.400 195.270 ;
        RECT 92.790 191.430 93.240 191.490 ;
        RECT 88.260 189.310 93.290 191.430 ;
        RECT 95.470 189.390 99.400 191.550 ;
        RECT 88.260 186.140 90.380 189.310 ;
        RECT 88.260 184.020 93.280 186.140 ;
        RECT 97.240 186.110 99.400 189.390 ;
        RECT 88.260 182.230 90.380 184.020 ;
        RECT 95.580 183.950 99.400 186.110 ;
        RECT 97.240 182.240 99.400 183.950 ;
        RECT 88.260 180.110 93.370 182.230 ;
        RECT 88.260 173.220 90.380 180.110 ;
        RECT 95.600 180.080 99.400 182.240 ;
        RECT 88.260 171.100 92.560 173.220 ;
        RECT 97.240 173.140 99.400 180.080 ;
        RECT 88.260 169.560 89.440 171.100 ;
        RECT 94.800 171.020 99.400 173.140 ;
        RECT 88.260 161.690 90.380 169.560 ;
        RECT 88.260 159.570 92.600 161.690 ;
        RECT 97.240 161.610 99.400 171.020 ;
        RECT 88.260 158.490 89.440 159.570 ;
        RECT 94.840 159.490 99.400 161.610 ;
        RECT 88.260 150.620 90.380 158.490 ;
        RECT 88.260 148.500 92.640 150.620 ;
        RECT 97.240 150.540 99.400 159.490 ;
        RECT 88.260 147.490 89.440 148.500 ;
        RECT 94.880 148.420 99.400 150.540 ;
        RECT 88.260 139.620 90.380 147.490 ;
        RECT 88.260 137.500 92.550 139.620 ;
        RECT 97.240 139.540 99.400 148.420 ;
        RECT 88.260 136.420 89.440 137.500 ;
        RECT 94.790 137.420 99.400 139.540 ;
        RECT 88.260 128.550 90.380 136.420 ;
        RECT 88.260 126.430 92.590 128.550 ;
        RECT 97.240 128.470 99.400 137.420 ;
        RECT 88.260 124.890 89.440 126.430 ;
        RECT 94.830 126.350 99.400 128.470 ;
        RECT 88.260 121.980 90.380 124.890 ;
        RECT 1.140 119.860 90.380 121.980 ;
        RECT 41.900 116.710 44.020 119.860 ;
        RECT 52.970 116.750 55.090 119.860 ;
        RECT 63.970 116.660 66.090 119.860 ;
        RECT 75.040 116.700 77.160 119.860 ;
        RECT 86.570 116.740 88.690 119.860 ;
        RECT 41.820 111.220 43.940 114.470 ;
        RECT 52.890 111.220 55.010 114.510 ;
        RECT 63.890 111.220 66.010 114.420 ;
        RECT 74.960 111.220 77.080 114.460 ;
        RECT 86.490 111.260 88.610 114.500 ;
        RECT 97.240 111.260 99.400 126.350 ;
        RECT 81.550 111.220 99.400 111.260 ;
        RECT 4.490 109.100 99.400 111.220 ;
        RECT 4.070 88.610 119.355 89.680 ;
        RECT 76.800 88.230 79.520 88.610 ;
        RECT 80.420 88.590 119.355 88.610 ;
        RECT 78.030 88.005 79.100 88.230 ;
        RECT 81.960 88.175 83.030 88.590 ;
        RECT 86.290 88.205 87.360 88.590 ;
        RECT 90.260 88.135 91.330 88.590 ;
        RECT 95.780 88.145 96.850 88.590 ;
        RECT 100.110 88.175 101.180 88.590 ;
        RECT 104.080 88.105 105.150 88.590 ;
        RECT 107.060 88.095 108.130 88.590 ;
        RECT 111.390 88.125 112.460 88.590 ;
        RECT 115.360 88.055 116.430 88.590 ;
        RECT 1.000 85.190 66.530 86.650 ;
        RECT 78.055 85.190 79.195 85.720 ;
        RECT 81.865 85.370 83.005 85.940 ;
        RECT 86.315 85.370 87.455 85.920 ;
        RECT 90.155 85.370 91.295 85.870 ;
        RECT 95.685 85.370 96.825 85.910 ;
        RECT 100.135 85.370 101.275 85.890 ;
        RECT 103.975 85.370 105.115 85.840 ;
        RECT 106.965 85.370 108.105 85.860 ;
        RECT 111.415 85.370 112.555 85.840 ;
        RECT 115.255 85.370 116.395 85.790 ;
        RECT 80.670 85.190 116.940 85.370 ;
        RECT 1.000 84.050 116.940 85.190 ;
        RECT 1.000 84.040 66.530 84.050 ;
        RECT 20.180 83.140 21.400 84.040 ;
        RECT 20.180 82.680 24.220 83.140 ;
        RECT 20.180 79.420 21.400 82.680 ;
        RECT 24.400 79.970 27.920 80.410 ;
        RECT 26.710 79.560 27.920 79.970 ;
        RECT 20.180 78.960 24.690 79.420 ;
        RECT 20.180 75.330 21.400 78.960 ;
        RECT 26.700 76.720 27.920 79.560 ;
        RECT 24.170 76.280 27.920 76.720 ;
        RECT 31.600 78.900 32.510 84.040 ;
        RECT 31.600 78.420 34.480 78.900 ;
        RECT 31.600 76.390 32.510 78.420 ;
        RECT 20.180 74.870 24.500 75.330 ;
        RECT 20.180 71.620 21.400 74.870 ;
        RECT 26.700 73.690 27.920 76.280 ;
        RECT 30.440 75.900 32.510 76.390 ;
        RECT 26.700 73.210 30.130 73.690 ;
        RECT 26.700 72.610 27.920 73.210 ;
        RECT 24.710 72.170 27.920 72.610 ;
        RECT 20.180 71.160 24.400 71.620 ;
        RECT 20.180 67.020 21.400 71.160 ;
        RECT 26.700 68.880 27.920 72.170 ;
        RECT 31.600 72.165 32.510 75.900 ;
        RECT 35.250 75.700 37.760 76.180 ;
        RECT 31.605 72.150 32.510 72.165 ;
        RECT 31.605 71.670 33.420 72.150 ;
        RECT 31.605 71.640 32.510 71.670 ;
        RECT 31.600 71.065 32.510 71.640 ;
        RECT 32.945 69.690 33.420 71.670 ;
        RECT 32.920 69.230 34.740 69.690 ;
        RECT 24.110 68.860 27.920 68.880 ;
        RECT 24.110 68.440 30.430 68.860 ;
        RECT 26.700 68.380 30.430 68.440 ;
        RECT 20.180 66.560 24.420 67.020 ;
        RECT 20.180 63.290 21.400 66.560 ;
        RECT 26.700 64.640 27.920 68.380 ;
        RECT 32.945 67.350 33.420 69.230 ;
        RECT 29.740 66.890 33.420 67.350 ;
        RECT 36.740 68.760 37.760 75.700 ;
        RECT 39.190 70.940 40.360 84.040 ;
        RECT 44.510 83.960 46.210 84.040 ;
        RECT 55.930 83.960 57.320 84.040 ;
        RECT 63.520 83.960 65.170 84.040 ;
        RECT 44.510 83.160 45.730 83.960 ;
        RECT 44.510 82.700 48.550 83.160 ;
        RECT 44.510 79.440 45.730 82.700 ;
        RECT 48.730 79.990 52.250 80.430 ;
        RECT 51.040 79.580 52.250 79.990 ;
        RECT 44.510 78.980 49.020 79.440 ;
        RECT 44.510 75.350 45.730 78.980 ;
        RECT 51.030 76.740 52.250 79.580 ;
        RECT 48.500 76.300 52.250 76.740 ;
        RECT 55.930 78.920 56.840 83.960 ;
        RECT 55.930 78.440 58.810 78.920 ;
        RECT 55.930 76.410 56.840 78.440 ;
        RECT 44.510 74.890 48.830 75.350 ;
        RECT 44.510 71.640 45.730 74.890 ;
        RECT 51.030 73.710 52.250 76.300 ;
        RECT 54.770 75.920 56.840 76.410 ;
        RECT 51.030 73.230 54.460 73.710 ;
        RECT 51.030 72.630 52.250 73.230 ;
        RECT 49.040 72.190 52.250 72.630 ;
        RECT 44.510 71.180 48.730 71.640 ;
        RECT 36.740 68.280 38.730 68.760 ;
        RECT 36.740 66.970 37.760 68.280 ;
        RECT 26.700 64.270 30.490 64.640 ;
        RECT 24.630 64.160 30.490 64.270 ;
        RECT 24.630 63.830 27.920 64.160 ;
        RECT 20.180 62.830 24.760 63.290 ;
        RECT 20.180 59.200 21.400 62.830 ;
        RECT 26.700 60.550 27.920 63.830 ;
        RECT 32.945 62.270 33.420 66.890 ;
        RECT 35.460 66.490 37.760 66.970 ;
        RECT 30.965 61.795 33.420 62.270 ;
        RECT 24.250 60.110 27.920 60.550 ;
        RECT 26.700 59.530 27.920 60.110 ;
        RECT 20.180 58.740 24.190 59.200 ;
        RECT 26.700 59.050 30.500 59.530 ;
        RECT 20.180 55.450 21.400 58.740 ;
        RECT 26.700 56.470 27.920 59.050 ;
        RECT 24.680 56.000 27.920 56.470 ;
        RECT 20.180 54.990 24.520 55.450 ;
        RECT 20.180 54.980 21.400 54.990 ;
        RECT 26.700 52.770 27.920 56.000 ;
        RECT 24.260 52.240 27.920 52.770 ;
        RECT 26.700 49.410 27.920 52.240 ;
        RECT 36.740 49.410 37.760 66.490 ;
        RECT 44.510 67.040 45.730 71.180 ;
        RECT 51.030 68.900 52.250 72.190 ;
        RECT 55.930 72.185 56.840 75.920 ;
        RECT 59.580 75.720 62.090 76.200 ;
        RECT 55.935 72.170 56.840 72.185 ;
        RECT 55.935 71.690 57.750 72.170 ;
        RECT 55.935 71.660 56.840 71.690 ;
        RECT 55.930 71.085 56.840 71.660 ;
        RECT 57.275 69.710 57.750 71.690 ;
        RECT 57.250 69.250 59.070 69.710 ;
        RECT 48.440 68.880 52.250 68.900 ;
        RECT 48.440 68.460 54.760 68.880 ;
        RECT 51.030 68.400 54.760 68.460 ;
        RECT 44.510 66.580 48.750 67.040 ;
        RECT 44.510 63.310 45.730 66.580 ;
        RECT 51.030 64.660 52.250 68.400 ;
        RECT 57.275 67.370 57.750 69.250 ;
        RECT 54.070 66.910 57.750 67.370 ;
        RECT 61.070 68.780 62.090 75.720 ;
        RECT 63.520 70.960 64.690 83.960 ;
        RECT 75.990 77.030 77.130 84.050 ;
        RECT 80.670 83.970 116.940 84.050 ;
        RECT 81.700 83.260 82.840 83.970 ;
        RECT 85.540 83.210 86.680 83.970 ;
        RECT 89.990 83.190 91.130 83.970 ;
        RECT 92.980 83.210 94.120 83.970 ;
        RECT 96.820 83.160 97.960 83.970 ;
        RECT 101.270 83.140 102.410 83.970 ;
        RECT 106.800 83.180 107.940 83.970 ;
        RECT 110.640 83.130 111.780 83.970 ;
        RECT 115.090 83.110 116.230 83.970 ;
        RECT 81.665 80.135 82.735 80.995 ;
        RECT 85.635 80.135 86.705 80.925 ;
        RECT 89.965 80.135 91.035 80.955 ;
        RECT 80.985 80.090 91.500 80.135 ;
        RECT 80.985 80.085 92.550 80.090 ;
        RECT 92.945 80.085 94.015 80.945 ;
        RECT 96.915 80.085 97.985 80.875 ;
        RECT 101.245 80.085 102.315 80.905 ;
        RECT 106.765 80.085 107.835 80.915 ;
        RECT 80.985 80.055 107.835 80.085 ;
        RECT 110.735 80.055 111.805 80.845 ;
        RECT 115.065 80.135 116.135 80.875 ;
        RECT 118.285 80.135 119.355 88.590 ;
        RECT 113.135 80.055 119.355 80.135 ;
        RECT 80.985 80.050 108.550 80.055 ;
        RECT 108.950 80.050 109.830 80.055 ;
        RECT 80.985 80.030 109.830 80.050 ;
        RECT 110.470 80.030 119.355 80.055 ;
        RECT 80.985 79.480 119.355 80.030 ;
        RECT 80.985 79.065 119.370 79.480 ;
        RECT 91.460 79.015 119.370 79.065 ;
        RECT 102.985 78.985 119.370 79.015 ;
        RECT 116.350 78.970 119.370 78.985 ;
        RECT 75.990 75.890 122.680 77.030 ;
        RECT 121.550 75.750 122.680 75.890 ;
        RECT 121.550 73.950 122.690 75.750 ;
        RECT 134.780 73.020 135.870 73.940 ;
        RECT 137.560 71.680 138.650 72.550 ;
        RECT 119.260 70.640 121.060 71.670 ;
        RECT 119.260 69.730 121.020 70.640 ;
        RECT 61.070 68.300 63.060 68.780 ;
        RECT 75.550 68.630 121.020 69.730 ;
        RECT 61.070 66.990 62.090 68.300 ;
        RECT 51.030 64.290 54.820 64.660 ;
        RECT 48.960 64.180 54.820 64.290 ;
        RECT 48.960 63.850 52.250 64.180 ;
        RECT 44.510 62.850 49.090 63.310 ;
        RECT 44.510 59.220 45.730 62.850 ;
        RECT 51.030 60.570 52.250 63.850 ;
        RECT 57.275 62.290 57.750 66.910 ;
        RECT 59.790 66.510 62.090 66.990 ;
        RECT 55.295 61.815 57.750 62.290 ;
        RECT 48.580 60.130 52.250 60.570 ;
        RECT 51.030 59.550 52.250 60.130 ;
        RECT 44.510 58.760 48.520 59.220 ;
        RECT 51.030 59.070 54.830 59.550 ;
        RECT 44.510 55.470 45.730 58.760 ;
        RECT 51.030 56.490 52.250 59.070 ;
        RECT 49.010 56.020 52.250 56.490 ;
        RECT 44.510 55.010 48.850 55.470 ;
        RECT 44.510 55.000 45.730 55.010 ;
        RECT 51.030 52.790 52.250 56.020 ;
        RECT 48.590 52.260 52.250 52.790 ;
        RECT 51.030 49.720 52.250 52.260 ;
        RECT 61.070 49.720 62.090 66.510 ;
        RECT 75.550 67.930 121.040 68.630 ;
        RECT 51.030 49.610 52.700 49.720 ;
        RECT 61.070 49.610 62.540 49.720 ;
        RECT 66.290 49.610 68.130 49.630 ;
        RECT 41.960 49.450 73.480 49.610 ;
        RECT 75.550 49.450 77.350 67.930 ;
        RECT 41.960 49.430 77.350 49.450 ;
        RECT 41.560 49.410 77.350 49.430 ;
        RECT 4.000 47.650 77.350 49.410 ;
        RECT 4.000 46.880 66.265 47.650 ;
        RECT 30.540 32.780 33.230 33.680 ;
        RECT 1.860 29.770 31.370 30.540 ;
        RECT 32.330 29.070 33.230 32.780 ;
        RECT 48.260 30.250 94.190 31.110 ;
        RECT 48.260 30.210 59.090 30.250 ;
        RECT 48.260 29.070 49.160 30.210 ;
        RECT 4.010 28.170 49.220 29.070 ;
        RECT 12.560 27.530 13.460 28.170 ;
        RECT 21.890 28.100 22.790 28.170 ;
        RECT 23.140 27.870 24.040 28.170 ;
        RECT 30.520 28.100 31.420 28.170 ;
        RECT 32.860 28.010 33.830 28.170 ;
        RECT 40.050 28.100 40.950 28.170 ;
        RECT 32.860 27.870 33.810 28.010 ;
        RECT 23.140 27.460 24.050 27.870 ;
        RECT 32.850 27.460 33.810 27.870 ;
        RECT 42.920 27.870 43.810 28.170 ;
        RECT 42.920 27.490 43.820 27.870 ;
        RECT 23.140 27.390 24.040 27.460 ;
        RECT 32.850 27.440 33.750 27.460 ;
        RECT 12.600 24.250 13.500 25.240 ;
        RECT 21.900 24.250 22.800 24.290 ;
        RECT 23.140 24.250 24.040 25.240 ;
        RECT 32.900 24.740 33.800 25.240 ;
        RECT 30.460 24.250 31.360 24.290 ;
        RECT 32.870 24.250 33.800 24.740 ;
        RECT 40.010 24.260 40.910 24.290 ;
        RECT 42.910 24.260 43.810 25.270 ;
        RECT 50.640 25.230 51.540 30.210 ;
        RECT 53.540 29.620 54.440 30.210 ;
        RECT 63.680 29.610 64.610 30.250 ;
        RECT 63.700 29.540 64.600 29.610 ;
        RECT 54.860 26.500 64.680 27.400 ;
        RECT 38.370 24.250 49.175 24.260 ;
        RECT 0.990 23.350 49.175 24.250 ;
        RECT 48.260 22.480 49.160 23.350 ;
        RECT 48.260 21.880 49.170 22.480 ;
        RECT 53.660 21.880 54.560 22.990 ;
        RECT 57.880 21.880 58.780 26.500 ;
        RECT 68.130 25.870 68.990 30.250 ;
        RECT 73.480 29.760 74.410 30.250 ;
        RECT 83.450 29.790 84.380 30.250 ;
        RECT 87.550 30.210 94.190 30.250 ;
        RECT 73.490 29.580 74.390 29.760 ;
        RECT 83.460 29.610 84.360 29.790 ;
        RECT 73.440 26.540 84.450 27.400 ;
        RECT 64.880 25.620 75.770 25.870 ;
        RECT 64.880 25.360 75.780 25.620 ;
        RECT 64.880 25.010 75.790 25.360 ;
        RECT 74.890 24.980 75.790 25.010 ;
        RECT 48.260 21.840 59.090 21.880 ;
        RECT 64.870 21.840 65.770 22.790 ;
        RECT 74.880 21.840 75.780 22.760 ;
        RECT 79.390 21.840 80.250 26.540 ;
        RECT 88.240 25.840 89.140 30.210 ;
        RECT 93.290 26.770 94.190 30.210 ;
        RECT 85.010 25.530 89.140 25.840 ;
        RECT 85.000 24.940 89.140 25.530 ;
        RECT 85.000 24.890 85.900 24.940 ;
        RECT 48.260 21.760 80.250 21.840 ;
        RECT 84.990 21.840 85.890 22.670 ;
        RECT 93.310 21.880 94.210 24.440 ;
        RECT 87.550 21.840 94.200 21.880 ;
        RECT 84.990 21.760 94.200 21.840 ;
        RECT 48.260 21.640 94.200 21.760 ;
        RECT 48.280 20.980 94.200 21.640 ;
        RECT 30.410 16.140 33.280 17.040 ;
        RECT 1.470 13.320 31.490 14.290 ;
        RECT 32.380 12.770 33.280 16.140 ;
        RECT 3.970 11.900 83.165 12.770 ;
        RECT 3.970 11.870 17.130 11.900 ;
        RECT 18.130 11.870 27.380 11.900 ;
        RECT 28.380 11.880 83.165 11.900 ;
        RECT 12.700 11.220 13.600 11.870 ;
        RECT 22.680 11.180 23.580 11.870 ;
        RECT 32.380 11.180 33.340 11.880 ;
        RECT 42.450 11.210 43.350 11.880 ;
        RECT 52.150 11.210 53.110 11.880 ;
        RECT 62.170 11.210 63.070 11.880 ;
        RECT 71.870 11.210 72.830 11.880 ;
        RECT 82.190 11.210 83.150 11.880 ;
        RECT 52.150 11.190 53.050 11.210 ;
        RECT 71.870 11.190 72.770 11.210 ;
        RECT 82.190 11.190 83.090 11.210 ;
        RECT 32.380 11.160 33.280 11.180 ;
        RECT 12.710 7.950 13.610 8.950 ;
        RECT 22.670 7.950 23.570 8.960 ;
        RECT 32.430 8.460 33.330 8.960 ;
        RECT 32.400 7.950 33.330 8.460 ;
        RECT 42.440 7.980 43.340 8.990 ;
        RECT 52.200 8.490 53.100 8.990 ;
        RECT 52.170 7.980 53.100 8.490 ;
        RECT 62.160 7.980 63.060 8.990 ;
        RECT 71.920 8.490 72.820 8.990 ;
        RECT 82.240 8.580 83.140 8.990 ;
        RECT 71.890 7.980 72.820 8.490 ;
        RECT 82.210 8.430 83.140 8.580 ;
        RECT 82.210 8.280 83.130 8.430 ;
        RECT 37.900 7.960 47.150 7.980 ;
        RECT 48.150 7.960 57.010 7.980 ;
        RECT 57.620 7.960 66.870 7.980 ;
        RECT 67.870 7.960 76.730 7.980 ;
        RECT 37.280 7.950 76.730 7.960 ;
        RECT 1.050 7.930 17.130 7.950 ;
        RECT 18.130 7.930 27.380 7.950 ;
        RECT 28.380 7.940 78.150 7.950 ;
        RECT 82.230 7.940 83.130 8.280 ;
        RECT 28.380 7.930 83.130 7.940 ;
        RECT 1.050 7.050 83.130 7.930 ;
      LAYER met4 ;
        RECT 94.150 220.840 94.450 224.760 ;
        RECT 92.950 219.150 95.650 220.840 ;
        RECT 135.550 73.940 135.850 224.760 ;
        RECT 134.780 73.020 135.870 73.940 ;
        RECT 138.310 72.550 138.610 224.760 ;
        RECT 137.560 71.680 138.650 72.550 ;
  END
END tt_um_ohmy90_adders
END LIBRARY

