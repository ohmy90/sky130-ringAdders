* NGSPICE file created from tt_um_ohmy90_flat_adders.ext - technology: sky130A

.subckt tt_um_ohmy90_flat_adders clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7] VDPWR VGND
X0 sky130_fd_sc_hd__dfxbp_1_3.CLK a_13161_23139# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X1 VDPWR VGND a_12281_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X2 VDPWR a_9703_16093# a_11501_15239# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X3 a_24234_14385# ui_in[0] a_24152_14385# VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.10855 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X4 VGND a_9381_11547# a_9715_11297# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X5 VGND a_18671_29731# a_18671_30311# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=3880,195
X6 a_14729_22875# sky130_fd_sc_hd__dfxbp_1_3.Q_N VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X7 a_16793_4785# a_15711_4547# a_17210_4895# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X8 VDPWR VGND a_16539_5473# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X9 a_16679_4895# VDPWR a_16583_4895# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X10 a_4711_15373# VGND a_4625_15373# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X11 a_5174_5409# VDPWR a_4423_5299# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X12 a_18625_4938# a_17733_4529# a_18553_4938# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=7728,268
X13 sky130_fd_sc_hd__inv_6_0.A sky130_fd_sc_hd__inv_4_0.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X14 VGND VGND a_9369_16343# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X15 VDPWR VGND a_2313_1791# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X16 sky130_fd_sc_hd__dfxbp_1_9.CLK a_18671_29731# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X17 a_12533_5715# a_11411_5471# a_12950_5825# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X18 a_14545_5467# a_14491_5723# a_14152_5441# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X19 a_1950_5025# a_2217_5025# a_2175_5051# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X20 a_12419_5825# VDPWR a_12323_5825# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X21 VDPWR a_12194_5433# a_12142_5459# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X22 a_16033_2159# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X23 a_18667_34470# a_18667_33636# a_18667_33834# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.07121 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X24 sky130_fd_sc_hd__dfxbp_1_6.Q_N a_18671_30311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3880,195 d=6760,364
X25 a_17236_5839# VDPWR a_16485_5729# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X26 a_4513_14775# VDPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X27 a_6129_12927# a_4913_13781# a_6057_12927# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=1764,126
X28 VGND VGND a_16297_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X29 sky130_fd_sc_hd__inv_4_0.A sky130_fd_sc_hd__inv_2_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X30 sky130_fd_sc_hd__dfxbp_1_8.Q_N a_18667_34839# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=6160,267 d=10400,504
X31 a_18697_29647# a_18671_29108# a_18671_29942# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X32 a_9715_11297# a_9381_11547# a_9631_11547# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X33 a_7113_13395# a_6862_13645# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4010,197 d=6760,364
X34 a_12323_5459# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X35 VGND a_19235_17155# a_18113_17153# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X36 a_11255_13773# a_10717_13773# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X37 VDPWR VGND a_7032_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X38 a_11501_15239# a_8193_13753# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X39 a_4383_2153# a_4329_2043# a_3990_1761# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X40 uo_out[0] sky130_fd_sc_hd__inv_16_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X41 a_14281_5833# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X42 VGND sky130_fd_sc_hd__inv_6_0.A sky130_fd_sc_hd__inv_8_0.A VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X43 VDPWR VGND a_4587_13107# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X44 a_9631_11297# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X45 a_8169_1793# VDPWR a_8073_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X46 a_14771_4803# a_13709_4553# a_15188_4547# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X47 a_22274_16171# a_21506_16181# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X48 a_2175_5417# VDPWR a_2079_5417# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X49 a_6089_11935# a_4849_11293# a_6003_11935# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X50 VDPWR VDPWR a_14596_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X51 VGND a_11888_1767# a_11836_1793# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X52 a_10289_2159# a_10235_2049# a_9896_1767# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X53 a_12697_14007# a_9781_10553# a_12615_14007# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2772,150
X54 VDPWR VGND a_4597_11543# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X55 a_7221_1787# a_6281_2043# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X56 sky130_fd_sc_hd__inv_8_0.A sky130_fd_sc_hd__inv_6_0.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X57 a_18671_29438# a_18671_29203# a_18697_29053# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.07505 ps=0.76615 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X58 a_18663_27120# a_18663_27252# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14038 pd=1.37821 as=0.15033 ps=1.4282 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X59 VDPWR VDPWR a_9491_15377# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X60 VDPWR VDPWR a_6792_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X61 VDPWR VDPWR a_14825_4547# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X62 a_12644_2159# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X63 VDPWR VDPWR a_16660_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X64 VDPWR VDPWR a_16847_4529# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X65 a_9629_14779# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X66 a_10525_5837# a_10471_5727# a_10132_5445# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X67 a_18693_24621# sky130_fd_sc_hd__dfxbp_1_5.Q_N VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08755 pd=0.89385 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X68 VDPWR VGND a_14233_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X69 a_5942_1761# a_5269_1787# a_6167_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X70 VGND a_18671_29731# a_19063_29704# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.07108 ps=0.80231 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X71 a_6238_6077# a_18625_4938# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=6334,279 d=10400,504
X72 a_18693_31479# a_18667_31449# a_18667_31684# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X73 VDPWR VDPWR a_10289_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X74 VGND a_1920_1765# a_1868_1791# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X75 a_8038_5023# a_7315_5043# a_8263_5049# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X76 VDPWR sky130_fd_sc_hd__inv_12_0.A sky130_fd_sc_hd__inv_16_0.A VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=20600,606
X77 sky130_fd_sc_hd__inv_12_0.A sky130_fd_sc_hd__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X78 a_18693_31299# sky130_fd_sc_hd__dfxbp_1_9.Q_N VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X79 VDPWR a_18671_29731# a_18697_29647# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X80 a_19059_25272# a_18667_24771# a_18667_25510# VGND sky130_fd_pr__special_nfet_01v8 ad=0.06092 pd=0.68769 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X81 VDPWR a_9556_17271# a_6629_15387# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X82 a_7126_5409# VDPWR a_6375_5299# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X83 VDPWR VDPWR a_4753_16339# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X84 VGND VGND a_5174_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X85 a_12769_4809# a_11439_4597# a_13186_4553# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X86 VGND sky130_fd_sc_hd__inv_2_0.A sky130_fd_sc_hd__inv_4_0.A VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X87 VDPWR a_18667_31552# a_18693_31479# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X88 a_17096_23241# a_16657_22875# a_17011_22875# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.07505 ps=0.76615 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X89 VDPWR VDPWR a_4746_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X90 VDPWR VDPWR a_8431_5049# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X91 VDPWR a_14982_22987# a_14909_23241# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X92 a_4903_15345# a_4625_15373# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X93 VDPWR sky130_fd_sc_hd__inv_16_0.A uo_out[0] VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X94 VGND sky130_fd_sc_hd__dfxbp_1_7.Q a_18671_29203# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X95 VGND a_15407_23143# a_15365_22875# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.07108 ps=0.80231 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X96 VDPWR VDPWR a_4763_14775# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X97 VDPWR VDPWR a_12823_4553# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X98 a_13520_4919# VDPWR a_12769_4809# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X99 a_18693_25215# a_18667_24676# a_18667_25510# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X100 a_4913_13781# a_4635_13809# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X101 VGND a_15693_17123# a_15641_17149# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X102 VGND VDPWR a_17210_4895# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X103 a_10160_4571# VDPWR a_10385_4963# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X104 a_4084_5017# a_3229_5051# a_4309_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X105 VGND VGND a_14930_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X106 a_8645_23241# a_7863_22875# a_8561_23241# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X107 a_17011_22875# sky130_fd_sc_hd__dfxbp_1_4.Q_N VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08755 pd=0.89385 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X108 a_16847_4895# a_15711_4547# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X109 VGND sky130_fd_sc_hd__inv_12_0.A sky130_fd_sc_hd__inv_16_0.A VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X110 a_4723_10577# VGND a_4637_10577# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X111 a_15431_5467# a_14491_5723# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X112 a_4587_13107# VDPWR a_4505_13107# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X113 VGND VGND a_9381_11547# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X114 a_16146_5447# a_15431_5467# a_16371_5839# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X115 a_14377_5467# VDPWR a_14281_5467# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X116 a_2079_5051# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X117 a_16902_5839# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X118 a_9223_1793# a_8283_2049# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X119 VGND VDPWR a_16539_5839# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X120 VDPWR a_17345_17163# a_16471_17161# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X121 a_4597_11543# VDPWR a_4515_11543# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X122 sky130_fd_sc_hd__inv_16_0.A sky130_fd_sc_hd__inv_12_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X123 a_9491_15377# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X124 a_6944_13645# a_6329_12927# a_6862_13645# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X125 a_10132_5445# VGND a_10357_5471# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X126 VGND a_13840_1767# a_13788_1793# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X127 a_8700_1793# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X128 a_4635_13809# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X129 a_2706_5417# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X130 VDPWR VGND a_2343_5051# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X131 VGND a_4513_14775# a_4847_14525# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X132 a_10986_2159# VDPWR a_10235_2049# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X133 a_4215_2153# VDPWR a_4119_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X134 sky130_fd_sc_hd__dfxbp_1_7.Q a_18663_27545# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X135 a_10550_22991# a_10382_23245# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.12659 pd=1.2736 as=0.12379 ps=1.28732 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X136 a_17096_23241# a_16823_22875# a_17011_22875# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X137 VGND a_11979_13399# a_12615_14007# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2268,138 d=4075,198
X138 VGND VGND a_12978_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X139 VGND a_17689_23143# a_18120_23197# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=3880,195
X140 a_9779_13785# a_9501_13813# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X141 a_10888_5471# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X142 a_18625_4938# a_17425_5473# a_18625_5265# VGND sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=3990,179
X143 VGND a_4503_16339# a_4837_16089# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X144 a_8337_1793# a_7221_1787# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X145 VGND VGND a_7126_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X146 VDPWR VDPWR a_10525_5471# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X147 a_14825_4547# a_13709_4553# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X148 VDPWR sky130_fd_sc_hd__inv_16_0.A uo_out[0] VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X149 a_18663_26922# a_18663_27017# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X150 VGND a_18667_25299# a_19059_25272# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.07108 ps=0.80231 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X151 a_8377_5305# a_7315_5043# a_8794_5415# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X152 VDPWR VDPWR a_9503_10581# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X153 VDPWR a_8038_5023# a_7986_5049# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X154 sky130_fd_sc_hd__inv_16_0.A sky130_fd_sc_hd__inv_12_0.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X155 a_11888_1767# a_11175_1793# a_12113_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X156 VGND sky130_fd_sc_hd__inv_16_0.A uo_out[0] VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X157 VGND a_9556_17271# a_23511_14335# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X158 VGND a_3990_1761# a_3938_1787# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X159 a_9371_13111# VDPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X160 VDPWR VDPWR a_6698_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X161 a_18689_26867# sky130_fd_sc_hd__dfxbp_1_7.Q_N VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08755 pd=0.89385 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X162 a_6805_15235# a_4847_14525# a_6717_15235# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X163 a_9705_12861# VDPWR a_9621_12861# VGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X164 VGND VGND a_13520_4919# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X165 VDPWR a_8729_23143# a_9160_23197# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.12828 pd=1.21873 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=6160,267
X166 sky130_fd_sc_hd__dfxbp_1_2.CLK a_10975_23147# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X167 VGND a_15239_23241# a_15407_23143# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X168 VDPWR VGND a_10289_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X169 a_8167_5049# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X170 a_1920_1765# a_2187_1765# a_2145_2157# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X171 a_5269_1787# a_4329_2043# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X172 sky130_fd_sc_hd__dfxbp_1_0.Q_N a_9160_23197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3880,195 d=6760,364
X173 a_15323_23241# a_14541_22875# a_15239_23241# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X174 VDPWR VDPWR a_13186_4553# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X175 a_10297_22879# sky130_fd_sc_hd__dfxbp_1_1.Q_N VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X176 a_16486_16197# a_15641_17149# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X177 a_23677_14701# ui_in[0] a_23761_14335# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.36 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=4316,272
X178 a_4905_12113# a_4627_12141# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X179 a_12823_4553# a_11439_4597# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X180 VGND a_18663_27756# a_18663_27545# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X181 a_4915_10549# a_4637_10577# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X182 VGND a_18663_27545# a_18663_28125# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=3880,195
X183 a_6087_14735# a_5809_14763# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X184 a_12793_14007# a_11147_11911# a_12697_14007# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X185 VGND VDPWR a_2313_2157# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X186 a_17521_23241# a_16823_22875# a_17264_22987# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.07121 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X187 VGND a_14152_5441# a_14100_5467# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X188 VDPWR VGND a_17236_5473# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X189 a_14940_22875# a_14541_22875# a_14814_23241# VGND sky130_fd_pr__special_nfet_01v8 ad=0.06425 pd=0.70615 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X190 a_7749_14003# a_7173_15235# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X191 VGND a_9317_5049# a_18371_4938# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=5796,222
X192 a_19059_31950# a_18667_31449# a_18667_32188# VGND sky130_fd_pr__special_nfet_01v8 ad=0.06092 pd=0.68769 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X193 a_4213_5409# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X194 a_10121_1793# VDPWR a_10025_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X195 a_4383_1787# a_3199_1791# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X196 a_10289_4963# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X197 VDPWR VGND a_3010_1791# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X198 a_14432_4521# a_13709_4553# a_14657_4913# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X199 a_12615_14007# a_12039_15239# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X200 a_12227_2049# a_11175_1793# a_12644_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X201 VDPWR a_7944_1767# a_7892_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X202 a_19059_24851# a_18667_24676# a_18667_25006# VGND sky130_fd_pr__special_nfet_01v8 ad=0.06425 pd=0.70615 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X203 uo_out[0] sky130_fd_sc_hd__inv_16_0.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X204 VGND a_18667_34259# a_18667_34839# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=3880,195
X205 a_4763_14525# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X206 a_16275_5839# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X207 a_17425_5473# a_16485_5729# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X208 a_18667_33834# a_18667_33966# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.12659 pd=1.2736 as=0.12379 ps=1.28732 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X209 a_18667_24676# a_18667_24771# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.12828 ps=1.21873 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X210 a_24962_14701# ui_in[1] a_24234_14385# VGND sky130_fd_pr__nfet_01v8 ad=0.15102 pd=1.285 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=6041,257
X211 VGND VGND a_16994_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X212 VDPWR a_10132_5445# a_10080_5471# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X213 VGND VGND a_16539_5839# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X214 a_15188_4913# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X215 a_18693_31893# a_18667_31354# a_18667_32188# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X216 a_18667_25510# a_18667_24771# a_18667_24874# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.07862 ps=0.77179 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X217 VGND VDPWR a_12587_5825# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X218 a_2259_2047# a_2187_1765# a_2676_1791# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X219 a_4746_2153# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X220 VGND VGND a_10553_4963# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X221 VGND sky130_fd_sc_hd__dfxbp_1_9.CLK a_18667_31449# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X222 VGND a_16471_17161# a_15693_17123# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X223 a_9503_10581# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X224 a_9781_10553# a_9503_10581# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X225 a_8337_2159# a_8283_2049# a_7944_1767# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X226 a_18667_24874# a_18667_25006# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14038 pd=1.37821 as=0.15033 ps=1.4282 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X227 VDPWR a_17689_23143# a_17605_23241# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X228 a_1950_5025# a_2217_5025# a_2175_5417# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X229 a_14179_2049# a_13167_1793# a_14596_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X230 a_10261_5471# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X231 a_10652_2159# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X232 a_18667_31354# a_18667_31449# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X233 a_8561_23241# a_7863_22875# a_8304_22987# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.07121 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X234 VGND a_10807_23245# a_10975_23147# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X235 a_15904_1767# a_15119_1793# a_16129_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X236 sky130_fd_sc_hd__dfxbp_1_5.Q_N a_18667_25879# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3880,195 d=6760,364
X237 a_12865_14007# a_12039_15239# a_12793_14007# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X238 VDPWR a_13161_23139# a_13592_23193# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.12828 pd=1.21873 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=6160,267
X239 VDPWR VGND a_9461_14779# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X240 a_7749_14003# a_4915_10549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4368,272 d=2772,150
X241 a_14541_22875# a_14375_22875# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X242 VDPWR VGND a_10525_5471# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X243 VDPWR sky130_fd_sc_hd__inv_12_0.A sky130_fd_sc_hd__inv_16_0.A VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X244 VDPWR sky130_fd_sc_hd__inv_6_0.A sky130_fd_sc_hd__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10800,508
X245 VGND VDPWR a_14233_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X246 a_18667_31684# a_18667_31449# a_18693_31299# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.07505 ps=0.76615 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X247 sky130_fd_sc_hd__dfxbp_1_7.CLK a_18667_25299# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X248 a_14982_22987# a_14814_23241# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.12659 pd=1.2736 as=0.12379 ps=1.28732 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X249 VDPWR a_22365_17147# a_21491_17145# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X250 VDPWR a_9317_5049# a_18839_4938# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=6334,279
X251 a_3040_5051# VDPWR a_2289_5307# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X252 a_5895_14763# a_4849_11293# a_5809_14763# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X253 a_8431_5415# a_7315_5043# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X254 a_18697_29233# a_18671_29203# a_18671_29438# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X255 VGND VDPWR a_4711_15373# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X256 VDPWR a_18667_25299# a_18667_25879# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.12828 pd=1.21873 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=6160,267
X257 VDPWR sky130_fd_sc_hd__dfxbp_1_5.CLK a_18667_24771# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.12828 pd=1.21873 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X258 VDPWR a_10550_22991# a_10477_23245# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X259 a_10508_22879# a_10109_22879# a_10382_23245# VGND sky130_fd_pr__special_nfet_01v8 ad=0.06425 pd=0.70615 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X260 a_14541_22875# a_14375_22875# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.12828 ps=1.21873 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X261 a_18697_29053# sky130_fd_sc_hd__dfxbp_1_6.Q_N VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X262 VGND a_6281_11907# a_7749_14003# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2772,150 d=2268,138
X263 a_10499_4853# VDPWR a_10916_4597# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X264 a_18671_29438# a_18671_29108# a_18697_29053# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X265 a_18693_24801# a_18667_24771# a_18667_25006# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X266 a_6335_1787# a_5269_1787# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X267 VDPWR sky130_fd_sc_hd__inv_8_0.A sky130_fd_sc_hd__inv_12_0.A VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X268 a_18667_32188# a_18667_31449# a_18667_31552# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.07862 ps=0.77179 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X269 a_18693_24621# sky130_fd_sc_hd__dfxbp_1_5.Q_N VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X270 VDPWR a_9896_1767# a_9844_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X271 a_18667_25006# a_18667_24676# a_18693_24621# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X272 VGND VDPWR a_6792_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X273 VGND VDPWR a_2676_2157# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X274 VGND VGND a_4513_14775# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X275 a_10717_13773# a_9703_16093# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X276 a_11810_13649# a_11195_12931# a_11728_13649# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X277 VGND VGND a_12281_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X278 a_16847_4529# a_16793_4785# a_16454_4503# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X279 a_16243_2049# a_15119_1793# a_16660_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X280 a_8304_22987# a_8136_23241# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14038 pd=1.37821 as=0.15033 ps=1.4282 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X281 a_10025_1793# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X282 VGND VGND a_2313_2157# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X283 a_8193_13753# a_7749_14003# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5930,268 d=10800,508
X284 a_14152_5441# a_13473_5459# a_14377_5467# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X285 sky130_fd_sc_hd__inv_16_0.A sky130_fd_sc_hd__inv_12_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X286 sky130_fd_sc_hd__inv_8_0.A sky130_fd_sc_hd__inv_6_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X287 sky130_fd_sc_hd__dfxbp_1_0.CLK a_24962_14701# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X288 a_4755_13107# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X289 a_12769_4809# a_11439_4597# a_13186_4919# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X290 VDPWR sky130_fd_sc_hd__inv_16_0.A uo_out[0] VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X291 VGND VDPWR a_9587_13813# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X292 a_9128_5049# VDPWR a_8377_5305# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X293 sky130_fd_sc_hd__inv_16_0.A sky130_fd_sc_hd__inv_12_0.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X294 VGND a_10975_23147# a_10933_22879# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.07108 ps=0.80231 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X295 a_5933_13769# a_4849_11293# a_5851_13769# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
X296 a_7032_2153# VDPWR a_6281_2043# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X297 VGND sky130_fd_sc_hd__inv_16_0.A uo_out[0] VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X298 a_12568_23237# a_12295_22871# a_12483_22871# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X299 VGND a_7113_13395# a_7749_14003# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2268,138 d=4075,198
X300 VGND a_9371_13111# a_9705_12861# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X301 a_10869_11939# a_9715_11297# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X302 VDPWR VDPWR a_12644_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X303 a_4765_11543# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X304 VGND VGND a_16847_4895# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X305 a_10109_22879# a_9943_22879# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X306 a_12993_23237# a_12295_22871# a_12736_22983# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.07121 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X307 a_13119_22871# a_12129_22871# a_12993_23237# VGND sky130_fd_pr__special_nfet_01v8 ad=0.06092 pd=0.68769 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X308 a_21506_16181# a_20384_16179# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X309 a_14561_4913# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X310 VGND VDPWR a_12823_4919# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X311 VGND sky130_fd_sc_hd__dfxbp_1_3.CLK a_14375_22875# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X312 VDPWR VDPWR a_4840_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X313 a_19063_29704# a_18671_29203# a_18671_29942# VGND sky130_fd_pr__special_nfet_01v8 ad=0.06092 pd=0.68769 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X314 VGND VGND a_12587_5825# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X315 a_3990_1761# a_3199_1791# a_4215_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X316 sky130_fd_sc_hd__dfxbp_1_2.CLK a_10975_23147# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X317 a_4503_16339# VDPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X318 VGND VGND a_14825_4913# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X319 VDPWR VDPWR a_16902_5473# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X320 a_8169_2159# VDPWR a_8073_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X321 VDPWR VGND a_3040_5051# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X322 VDPWR sky130_fd_sc_hd__inv_16_0.A uo_out[0] VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X323 a_10109_22879# a_9943_22879# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.12828 ps=1.21873 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X324 VDPWR sky130_fd_sc_hd__dfxbp_1_2.CLK a_12129_22871# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.12828 pd=1.21873 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X325 VGND a_18667_34470# a_18667_34259# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X326 sky130_fd_sc_hd__dfxbp_1_7.Q_N a_18663_28125# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=6160,267 d=10400,504
X327 VDPWR sky130_fd_sc_hd__dfxbp_1_3.CLK a_14375_22875# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.12828 pd=1.21873 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X328 VDPWR a_11255_13773# a_11810_13649# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5830,267
X329 a_2079_5417# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X330 a_3229_5051# a_2289_5307# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X331 VGND VDPWR a_14596_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X332 VDPWR sky130_fd_sc_hd__inv_8_0.A sky130_fd_sc_hd__inv_12_0.A VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X333 VDPWR a_18667_34259# a_18693_34175# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X334 VGND a_18667_33834# a_19059_33811# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.07495 ps=0.82385 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X335 VGND a_6238_6077# a_2217_5025# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X336 VGND sky130_fd_sc_hd__inv_8_0.A sky130_fd_sc_hd__inv_12_0.A VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X337 VGND VDPWR a_4383_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X338 VGND a_18667_31977# a_19059_31950# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.07108 ps=0.80231 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X339 a_17647_22875# a_16657_22875# a_17521_23241# VGND sky130_fd_pr__special_nfet_01v8 ad=0.06092 pd=0.68769 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X340 VGND VDPWR a_16660_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X341 a_11250_4963# VDPWR a_10499_4853# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X342 a_10132_5445# VGND a_10357_5837# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X343 a_2289_5307# a_2217_5025# a_2706_5051# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X344 a_23761_14335# a_23731_14309# a_23677_14335# VGND sky130_fd_pr__nfet_01v8 ad=0.09322 pd=1.07 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3409,185
X345 a_6389_13769# a_5851_13769# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X346 VGND VGND a_14233_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X347 a_17222_22875# a_16823_22875# a_17096_23241# VGND sky130_fd_pr__special_nfet_01v8 ad=0.06425 pd=0.70615 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X348 uo_out[0] sky130_fd_sc_hd__inv_16_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X349 VDPWR a_4903_15345# a_5851_13769# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X350 VGND VGND a_2343_5417# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X351 uo_out[0] sky130_fd_sc_hd__inv_16_0.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X352 VGND sky130_fd_sc_hd__inv_12_0.A sky130_fd_sc_hd__inv_16_0.A VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X353 VGND VDPWR a_10289_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X354 uo_out[0] sky130_fd_sc_hd__inv_16_0.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X355 VDPWR VDPWR a_2343_5051# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X356 a_9451_16343# VDPWR a_9369_16343# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X357 a_10888_5837# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X358 a_12736_22983# a_12568_23237# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14038 pd=1.37821 as=0.15033 ps=1.4282 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X359 a_9379_14779# VDPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X360 VGND VDPWR a_4723_10577# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X361 VGND VDPWR a_10525_5837# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X362 VDPWR VGND a_10986_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X363 sky130_fd_sc_hd__dfxbp_1_4.Q_N a_18120_23197# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=6160,267 d=10400,504
X364 VDPWR VDPWR a_9619_16343# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X365 a_4625_15373# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X366 a_10675_14767# a_9715_11297# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X367 a_9713_14529# VDPWR a_9629_14529# VGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X368 a_11222_5471# VDPWR a_10471_5727# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X369 a_19510_16177# a_18742_16187# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X370 a_9587_13813# VGND a_9501_13813# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X371 VGND VDPWR a_14908_5833# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X372 a_10553_4597# VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X373 VDPWR sky130_fd_sc_hd__inv_4_0.A sky130_fd_sc_hd__inv_6_0.A VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X374 VDPWR a_18667_25510# a_18667_25299# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X375 a_14491_5723# a_13473_5459# a_14908_5833# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X376 VDPWR VGND a_9128_5049# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X377 a_9769_15349# a_9491_15377# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X378 VDPWR a_11979_13399# a_12865_14007# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=5930,268
X379 a_11175_1793# a_10235_2049# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X380 a_16793_4785# a_15711_4547# a_17210_4529# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X381 a_17733_4529# a_16793_4785# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X382 VGND a_10160_4571# a_10108_4597# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X383 a_24774_14701# ui_in[1] VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X384 a_16679_4529# VDPWR a_16583_4529# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X385 a_14657_4547# VDPWR a_14561_4547# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X386 uo_out[0] sky130_fd_sc_hd__inv_16_0.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X387 sky130_fd_sc_hd__inv_12_0.A sky130_fd_sc_hd__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X388 a_8687_22875# a_7697_22875# a_8561_23241# VGND sky130_fd_pr__special_nfet_01v8 ad=0.06092 pd=0.68769 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X389 a_9896_1767# a_9223_1793# a_10121_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X390 sky130_fd_sc_hd__inv_6_0.A sky130_fd_sc_hd__inv_4_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X391 a_18742_16187# a_18128_16189# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X392 sky130_fd_sc_hd__inv_12_0.A sky130_fd_sc_hd__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X393 VDPWR a_10807_23245# a_10975_23147# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X394 VDPWR a_15407_23143# a_15838_23197# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.12828 pd=1.21873 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=6160,267
X395 VDPWR VDPWR a_4635_13809# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X396 a_9317_5049# a_8377_5305# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X397 a_8431_5415# a_8377_5305# a_8038_5023# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X398 a_14909_23241# a_14375_22875# a_14814_23241# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X399 a_6281_2043# a_5269_1787# a_6698_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X400 sky130_fd_sc_hd__dfxbp_1_3.Q_N a_15838_23197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3880,195 d=6760,364
X401 a_6375_5299# a_5363_5043# a_6792_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X402 VGND VDPWR a_13186_4919# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X403 a_9705_12861# a_9371_13111# a_9621_13111# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X404 a_13167_1793# a_12227_2049# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X405 a_12823_4919# a_11439_4597# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X406 VGND sky130_fd_sc_hd__inv_16_0.A uo_out[0] VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X407 VDPWR a_9556_17271# a_23511_14701# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X408 a_11979_13399# a_11728_13649# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5830,267 d=13600,536
X409 a_6335_1787# a_6281_2043# a_5942_1761# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X410 VDPWR a_6208_2817# a_2187_1765# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X411 a_13709_4553# a_12769_4809# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X412 a_23133_17137# a_22274_16171# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X413 a_23761_14335# a_24774_14701# a_24962_14701# VGND sky130_fd_pr__nfet_01v8 ad=0.09322 pd=1.07 as=0.15102 ps=1.285 w=0.42 l=0.15
**devattr s=6041,257 d=4368,272
X414 a_6057_12927# a_4849_11293# a_5975_12927# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X415 a_8700_2159# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X416 VGND VDPWR a_6335_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X417 a_17011_22875# sky130_fd_sc_hd__dfxbp_1_4.Q_N VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X418 VGND VGND a_17236_5839# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X419 a_3199_1791# a_2259_2047# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X420 VGND VGND a_11250_4963# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X421 a_23677_14335# a_23133_17137# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X422 VDPWR VGND a_14545_5467# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X423 VGND VGND a_9371_13111# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X424 VDPWR a_9771_12117# a_10869_11939# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X425 a_4119_2153# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X426 a_12655_4553# VDPWR a_12559_4553# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X427 VDPWR sky130_fd_sc_hd__inv_12_0.A sky130_fd_sc_hd__inv_16_0.A VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X428 VGND a_6389_13769# a_6862_13645# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4010,197
X429 a_18625_5265# a_18371_4938# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=5796,222 d=2772,150
X430 a_12281_1793# a_11175_1793# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X431 a_8337_2159# a_7221_1787# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X432 sky130_fd_sc_hd__dfxbp_1_9.Q_N a_18667_32557# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3880,195 d=6760,364
X433 a_18667_25510# a_18667_24676# a_18667_24874# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.07121 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X434 sky130_fd_sc_hd__dfxbp_1_4.CLK a_15407_23143# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X435 a_17544_4895# VDPWR a_16793_4785# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X436 a_4477_5043# a_3229_5051# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X437 a_9619_16343# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X438 a_9629_14529# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X439 sky130_fd_sc_hd__dfxbp_1_9.Q a_18667_31977# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X440 a_12483_22871# sky130_fd_sc_hd__dfxbp_1_2.Q_N VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X441 VDPWR VGND a_11222_5471# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X442 a_2313_1791# a_2187_1765# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X443 a_8051_22875# sky130_fd_sc_hd__dfxbp_1_0.Q_N VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08755 pd=0.89385 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X444 a_5975_12927# a_4913_13781# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0805 pd=0.94333 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2646,147
X445 a_13284_5825# VDPWR a_12533_5715# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X446 VGND VGND a_4383_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X447 a_10916_4963# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X448 VGND sky130_fd_sc_hd__inv_4_0.A sky130_fd_sc_hd__inv_6_0.A VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X449 VDPWR VDPWR a_2706_5051# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X450 a_15522_4913# VDPWR a_14771_4803# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X451 VGND VDPWR a_10553_4963# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X452 VDPWR a_18667_31977# a_18667_32557# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.12828 pd=1.21873 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=6160,267
X453 VGND a_4837_16089# a_6911_15235# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X454 VGND VGND a_10289_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X455 a_11195_12931# a_10841_12931# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5689,267 d=10400,504
X456 a_10261_5837# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X457 a_11411_5471# a_10471_5727# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X458 a_18671_29942# a_18671_29203# a_18671_29306# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.07862 ps=0.77179 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X459 a_9463_11547# VDPWR a_9381_11547# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X460 VDPWR a_18667_33834# a_18693_33761# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X461 a_18667_31684# a_18667_31354# a_18693_31299# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X462 VGND VGND a_10525_5837# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X463 a_4847_14525# VDPWR a_4763_14525# VGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X464 VDPWR VDPWR a_9631_11547# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X465 a_9034_1793# VDPWR a_8283_2049# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X466 VGND a_14432_4521# a_14380_4547# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X467 a_18671_29306# a_18671_29438# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14038 pd=1.37821 as=0.15033 ps=1.4282 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X468 a_15119_1793# a_14179_2049# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X469 VGND a_16454_4503# a_16402_4529# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X470 sky130_fd_sc_hd__inv_16_0.A sky130_fd_sc_hd__inv_12_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X471 a_3040_5417# VDPWR a_2289_5307# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X472 VDPWR VDPWR a_12950_5459# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X473 sky130_fd_sc_hd__inv_8_0.A sky130_fd_sc_hd__inv_6_0.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=9880,412 d=3510,184
X474 a_18667_32188# a_18667_31354# a_18667_31552# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.07121 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X475 a_14545_5833# a_13473_5459# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X476 a_6208_2817# a_16243_2049# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X477 VDPWR VDPWR a_17210_4529# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X478 VDPWR VDPWR a_15188_4547# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X479 a_4713_12141# VGND a_4627_12141# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X480 a_12587_5459# a_11411_5471# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X481 a_10121_2159# VDPWR a_10025_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X482 a_16847_4529# a_15711_4547# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X483 VDPWR a_20109_17157# a_19235_17155# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X484 VGND a_6036_5017# a_5984_5043# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X485 a_6792_5043# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X486 VGND VGND a_3010_2157# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X487 VDPWR a_18667_32188# a_18667_31977# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X488 a_18663_27252# a_18663_27017# a_18689_26867# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.07505 ps=0.76615 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X489 a_12227_2049# a_11175_1793# a_12644_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X490 a_6717_15235# a_6629_15387# a_6635_15235# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
X491 a_8263_5415# VDPWR a_8167_5415# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X492 VDPWR VDPWR a_10652_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X493 a_4837_16089# a_4503_16339# a_4753_16339# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X494 a_14233_1793# a_13167_1793# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X495 VGND a_10550_22991# a_10508_22879# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.07495 ps=0.82385 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X496 a_6071_2153# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X497 a_6429_5043# a_5363_5043# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X498 VGND VGND a_17544_4895# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X499 VDPWR VDPWR a_8794_5049# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X500 a_10891_23245# a_10109_22879# a_10807_23245# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X501 a_16297_1793# a_15119_1793# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X502 a_6167_1787# VDPWR a_6071_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X503 a_2259_2047# a_2187_1765# a_2676_2157# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X504 VGND a_12430_4527# a_12378_4553# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X505 VGND a_9379_14779# a_9713_14529# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X506 a_10553_4597# a_10499_4853# a_10160_4571# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X507 VDPWR sky130_fd_sc_hd__inv_8_0.A sky130_fd_sc_hd__inv_12_0.A VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X508 a_4753_16089# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X509 VDPWR a_4849_11293# a_5975_12927# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0805 ps=0.94333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X510 VGND VGND a_6335_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X511 a_19063_29283# a_18671_29108# a_18671_29438# VGND sky130_fd_pr__special_nfet_01v8 ad=0.06425 pd=0.70615 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X512 VGND a_4839_12857# a_5895_14763# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X513 a_12483_22871# sky130_fd_sc_hd__dfxbp_1_2.Q_N VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08755 pd=0.89385 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X514 VGND VGND a_13284_5825# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X515 sky130_fd_sc_hd__inv_4_0.A sky130_fd_sc_hd__inv_2_0.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X516 VGND VGND a_15522_4913# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X517 VDPWR VGND a_8431_5049# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X518 a_12039_15239# a_11501_15239# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X519 a_16454_4503# a_15711_4547# a_16679_4895# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X520 uo_out[0] sky130_fd_sc_hd__inv_16_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X521 sky130_fd_sc_hd__dfxbp_1_6.Q_N a_18671_30311# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=6160,267 d=10400,504
X522 a_18128_16189# a_17254_16187# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X523 a_9771_12117# a_9493_12145# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X524 a_17210_4895# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X525 uo_out[0] sky130_fd_sc_hd__inv_16_0.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X526 VDPWR VDPWR a_9493_12145# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X527 VGND VDPWR a_4840_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X528 VGND VDPWR a_10916_4963# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X529 a_12194_5433# a_11411_5471# a_12419_5825# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X530 a_15242_5467# VDPWR a_14491_5723# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X531 a_9556_17271# a_12615_14007# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4075,198 d=7020,368
X532 a_12950_5825# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X533 VGND a_9556_17271# a_6629_15387# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X534 VGND VDPWR a_16902_5839# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X535 a_16823_22875# a_16657_22875# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X536 VGND VGND a_3040_5417# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X537 VGND a_4505_13107# a_4839_12857# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X538 a_10953_14739# a_10675_14767# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X539 VDPWR VDPWR a_4755_13107# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X540 a_4477_5043# a_4423_5299# a_4084_5017# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X541 a_16823_22875# a_16657_22875# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.12828 ps=1.21873 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X542 a_4905_12113# a_4627_12141# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X543 a_2289_5307# a_2217_5025# a_2706_5417# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X544 a_7944_1767# a_7221_1787# a_8169_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X545 a_5080_2153# VDPWR a_4329_2043# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X546 VGND sky130_fd_sc_hd__inv_12_0.A sky130_fd_sc_hd__inv_16_0.A VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=13390,466
X547 VGND a_18663_27545# a_19055_27518# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.07108 ps=0.80231 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X548 a_8136_23241# a_7697_22875# a_8051_22875# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.07505 ps=0.76615 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X549 VDPWR a_6238_6077# a_24407_14651# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.09013 ps=0.995 w=0.42 l=0.15
**devattr s=3605,199 d=2268,138
X550 VDPWR VDPWR a_4765_11543# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X551 a_18671_29108# a_18671_29203# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.12828 ps=1.21873 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X552 VDPWR VDPWR a_10888_5471# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X553 VDPWR a_15904_1767# a_15852_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X554 a_16539_5473# a_16485_5729# a_16146_5447# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X555 a_10471_5727# VGND a_10888_5471# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X556 a_16243_2049# a_15119_1793# a_16660_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X557 a_10807_23245# a_9943_22879# a_10550_22991# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.07862 ps=0.77179 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X558 VDPWR VDPWR a_8337_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X559 VDPWR a_18663_27545# a_18689_27461# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X560 a_10477_23245# a_9943_22879# a_10382_23245# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X561 a_13969_1793# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X562 a_10025_2159# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X563 sky130_fd_sc_hd__dfxbp_1_1.Q_N a_11406_23201# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3880,195 d=6760,364
X564 VGND VGND a_4503_16339# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X565 VGND VDPWR a_2343_5417# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X566 a_8794_5415# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X567 a_7221_1787# a_6281_2043# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X568 VGND sky130_fd_sc_hd__inv_16_0.A uo_out[0] VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X569 sky130_fd_sc_hd__dfxbp_1_4.CLK a_15407_23143# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X570 VGND a_17264_22987# a_17222_22875# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.07495 ps=0.82385 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X571 a_9621_13111# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X572 a_11222_5837# VDPWR a_10471_5727# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X573 VGND sky130_fd_sc_hd__dfxbp_1_7.CLK a_18663_27017# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X574 a_12295_22871# a_12129_22871# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.12828 ps=1.21873 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X575 VGND a_17345_17163# a_16471_17161# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X576 VGND VDPWR a_12644_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X577 a_6698_1787# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X578 a_20384_16179# a_19510_16177# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X579 a_6238_6077# a_18625_4938# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4514,209 d=6760,364
X580 sky130_fd_sc_hd__dfxbp_1_2.Q_N a_13592_23193# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=6160,267 d=10400,504
X581 a_9493_12145# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X582 a_17254_16187# a_16486_16197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X583 VGND VDPWR a_9577_15377# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X584 a_6862_13645# a_6329_12927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X585 a_12587_5459# a_12533_5715# a_12194_5433# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X586 a_10385_4597# VDPWR a_10289_4597# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X587 a_14825_4547# a_14771_4803# a_14432_4521# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X588 VDPWR VGND a_15242_5467# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X589 VGND a_14982_22987# a_14940_22875# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.07495 ps=0.82385 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X590 sky130_fd_sc_hd__inv_16_0.A sky130_fd_sc_hd__inv_12_0.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X591 VDPWR a_18671_29942# a_18671_29731# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X592 a_5851_13769# a_4849_11293# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X593 a_4721_13809# VGND a_4635_13809# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X594 a_6375_5299# a_5363_5043# a_6792_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X595 a_14545_5833# a_14491_5723# a_14152_5441# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X596 VDPWR a_15693_17123# a_15641_17149# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X597 VDPWR VGND a_9451_16343# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X598 VDPWR a_4847_14525# a_6635_15235# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X599 VGND VGND a_9379_14779# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X600 a_18667_33636# a_18667_33731# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X601 sky130_fd_sc_hd__dfxbp_1_7.CLK a_18667_25299# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X602 a_8136_23241# a_7863_22875# a_8051_22875# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X603 VGND a_8729_23143# a_9160_23197# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=3880,195
X604 VDPWR a_9705_12861# a_10675_14767# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X605 a_16583_4895# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X606 a_18663_26922# a_18663_27017# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.12828 ps=1.21873 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X607 VDPWR VDPWR a_4625_15373# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X608 a_6429_5043# a_6375_5299# a_6036_5017# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X609 a_15431_5467# a_14491_5723# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X610 a_16297_1793# a_16243_2049# a_15904_1767# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X611 VGND a_18113_17153# a_17345_17163# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X612 a_14233_1793# a_14179_2049# a_13840_1767# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X613 a_18667_33966# a_18667_33731# a_18693_33581# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.07505 ps=0.76615 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X614 VGND VGND a_5080_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X615 a_18693_33581# sky130_fd_sc_hd__dfxbp_1_8.Q_N VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08755 pd=0.89385 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X616 a_7113_13395# a_6862_13645# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5830,267 d=13600,536
X617 a_12323_5825# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X618 a_12978_1793# VDPWR a_12227_2049# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X619 a_14908_5467# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X620 a_12568_23237# a_12129_22871# a_12483_22871# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.07505 ps=0.76615 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X621 a_12655_4919# VDPWR a_12559_4919# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X622 VDPWR VDPWR a_14545_5467# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X623 VGND sky130_fd_sc_hd__inv_16_0.A uo_out[0] VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X624 a_12823_4553# a_12769_4809# a_12430_4527# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X625 VGND VGND a_10986_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X626 a_14771_4803# a_13709_4553# a_15188_4913# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X627 VDPWR a_15239_23241# a_15407_23143# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X628 a_9631_11547# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X629 a_4477_5409# a_3229_5051# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X630 a_4329_2043# a_3199_1791# a_4746_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X631 a_11255_13773# a_10717_13773# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X632 a_5363_5043# a_4423_5299# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X633 a_4423_5299# a_3229_5051# a_4840_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X634 a_24774_14701# ui_in[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X635 a_4309_5043# VDPWR a_4213_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X636 a_17521_23241# a_16657_22875# a_17264_22987# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.07862 ps=0.77179 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X637 VGND VGND a_11222_5837# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X638 a_17191_23241# a_16657_22875# a_17096_23241# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X639 a_23677_14701# a_23133_17137# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.36 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X640 a_8073_1793# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X641 a_4383_1787# a_4329_2043# a_3990_1761# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X642 VGND VDPWR a_14825_4913# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X643 a_16485_5729# a_15431_5467# a_16902_5473# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X644 a_18667_31552# a_18667_31684# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14038 pd=1.37821 as=0.15033 ps=1.4282 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X645 a_17264_22987# a_17096_23241# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.12659 pd=1.2736 as=0.12379 ps=1.28732 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X646 VGND VGND a_4505_13107# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X647 VGND VDPWR a_2706_5417# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X648 VGND a_21491_17145# a_20877_17147# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X649 a_18693_34175# a_18667_33636# a_18667_34470# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X650 a_18671_29942# a_18671_29108# a_18671_29306# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.07121 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X651 a_9896_1767# a_9223_1793# a_10121_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X652 VDPWR a_5942_1761# a_5890_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X653 VGND a_9317_5049# a_18846_5265# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=4514,209
X654 VDPWR sky130_fd_sc_hd__inv_12_0.A sky130_fd_sc_hd__inv_16_0.A VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X655 VGND sky130_fd_sc_hd__dfxbp_1_9.Q a_18667_33731# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X656 a_9577_15377# VGND a_9491_15377# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X657 a_10993_13773# a_9703_16093# a_10887_13773# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X658 VDPWR VGND a_8337_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X659 sky130_fd_sc_hd__dfxbp_1_0.CLK a_24962_14701# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X660 a_2145_1791# VDPWR a_2049_1791# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X661 VDPWR a_17264_22987# a_17191_23241# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X662 a_8038_5023# a_7315_5043# a_8263_5415# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X663 a_10525_5471# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X664 a_15239_23241# a_14375_22875# a_14982_22987# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.07862 ps=0.77179 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X665 a_5809_14763# a_4849_11293# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X666 sky130_fd_sc_hd__inv_16_0.A sky130_fd_sc_hd__inv_12_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X667 VGND VDPWR a_8431_5415# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X668 a_10550_22991# a_10382_23245# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14038 pd=1.37821 as=0.15033 ps=1.4282 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X669 VDPWR VGND a_16847_4529# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X670 a_18667_24874# a_18667_25006# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.12659 pd=1.2736 as=0.12379 ps=1.28732 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X671 a_5942_1761# a_5269_1787# a_6167_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X672 VGND a_13161_23139# a_13592_23193# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=3880,195
X673 VDPWR sky130_fd_sc_hd__dfxbp_1_9.CLK a_18667_31449# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.12828 pd=1.21873 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X674 a_18689_26867# sky130_fd_sc_hd__dfxbp_1_7.Q_N VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X675 VGND sky130_fd_sc_hd__dfxbp_1_2.CLK a_12129_22871# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X676 VDPWR a_4837_16089# a_6635_15235# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X677 VGND a_20877_17147# a_20109_17157# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X678 a_13473_5459# a_12533_5715# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X679 a_12533_5715# a_11411_5471# a_12950_5459# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X680 VGND VGND a_7032_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X681 a_15711_4547# a_14771_4803# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X682 a_12559_4553# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X683 sky130_fd_sc_hd__inv_12_0.A sky130_fd_sc_hd__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X684 a_19059_31529# a_18667_31354# a_18667_31684# VGND sky130_fd_pr__special_nfet_01v8 ad=0.06425 pd=0.70615 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X685 a_8304_22987# a_8136_23241# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.12659 pd=1.2736 as=0.12379 ps=1.28732 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X686 a_6792_5409# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X687 a_12419_5459# VDPWR a_12323_5459# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X688 a_12281_2159# a_11175_1793# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X689 a_18667_31354# a_18667_31449# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.12828 ps=1.21873 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X690 VDPWR a_8729_23143# a_8645_23241# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X691 a_14377_5833# VDPWR a_14281_5833# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X692 VDPWR a_14152_5441# a_14100_5467# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X693 a_10235_2049# a_9223_1793# a_10652_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X694 a_14930_1793# VDPWR a_14179_2049# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X695 a_16994_1793# VDPWR a_16243_2049# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X696 VDPWR VGND a_9463_11547# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X697 a_6429_5409# a_5363_5043# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X698 a_7315_5043# a_6375_5299# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X699 a_2313_2157# a_2187_1765# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X700 VDPWR sky130_fd_sc_hd__inv_16_0.A uo_out[0] VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X701 VGND a_18671_29306# a_19063_29283# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.07495 ps=0.82385 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X702 sky130_fd_sc_hd__dfxbp_1_5.CLK a_17689_23143# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X703 VDPWR VDPWR a_9501_13813# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X704 a_14065_1793# VDPWR a_13969_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X705 a_16129_1793# VDPWR a_16033_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X706 a_22274_16171# a_21506_16181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X707 a_4505_13107# VDPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X708 a_14281_5467# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X709 VDPWR sky130_fd_sc_hd__inv_6_0.A sky130_fd_sc_hd__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X710 VGND a_7944_1767# a_7892_1793# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X711 a_6635_15235# a_6629_15387# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X712 VGND VDPWR a_4713_12141# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X713 a_6261_5043# VDPWR a_6165_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X714 VGND sky130_fd_sc_hd__inv_6_0.A sky130_fd_sc_hd__inv_8_0.A VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=7020,368
X715 a_18667_31552# a_18667_31684# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.12659 pd=1.2736 as=0.12379 ps=1.28732 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X716 VGND VGND a_4515_11543# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X717 VGND sky130_fd_sc_hd__inv_12_0.A sky130_fd_sc_hd__inv_16_0.A VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X718 VGND a_4084_5017# a_4032_5043# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X719 VGND a_18667_25510# a_18667_25299# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X720 a_4840_5043# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X721 VGND a_18667_24874# a_19059_24851# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.07495 ps=0.82385 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X722 sky130_fd_sc_hd__dfxbp_1_5.Q_N a_18667_25879# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=6160,267 d=10400,504
X723 a_8051_22875# sky130_fd_sc_hd__dfxbp_1_0.Q_N VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X724 VGND a_16146_5447# a_16094_5473# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X725 a_9034_2159# VDPWR a_8283_2049# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X726 a_9769_15349# a_9491_15377# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X727 VGND VDPWR a_4746_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X728 a_14825_4913# a_13709_4553# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X729 VDPWR a_18663_27545# a_18663_28125# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.12828 pd=1.21873 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=6160,267
X730 a_18689_27047# a_18663_27017# a_18663_27252# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X731 VGND a_23133_17137# a_22365_17147# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X732 a_2676_1791# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X733 VGND sky130_fd_sc_hd__inv_8_0.A sky130_fd_sc_hd__inv_12_0.A VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X734 a_11671_15239# a_9713_14529# a_11583_15239# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X735 a_9779_13785# a_9501_13813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X736 a_4215_1787# VDPWR a_4119_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X737 uo_out[0] sky130_fd_sc_hd__inv_16_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X738 a_11195_12931# a_10841_12931# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=5266,228 d=6760,364
X739 a_4837_16089# VDPWR a_4753_16089# VGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X740 a_16539_5473# a_15431_5467# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X741 VDPWR a_18663_27120# a_18689_27047# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X742 a_4913_13781# a_4635_13809# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X743 VDPWR a_4839_12857# a_5975_12927# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0805 ps=0.94333 w=0.42 l=0.15
**devattr s=2646,147 d=5689,267
X744 a_6329_12927# a_5975_12927# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5689,267 d=10400,504
X745 VGND a_1950_5025# a_1898_5051# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X746 a_8167_5415# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X747 VGND VDPWR a_10652_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X748 a_4477_5409# a_4423_5299# a_4084_5017# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X749 a_14233_2159# a_13167_1793# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X750 a_12736_22983# a_12568_23237# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.12659 pd=1.2736 as=0.12379 ps=1.28732 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X751 VGND VDPWR a_10888_5837# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X752 a_16539_5839# a_16485_5729# a_16146_5447# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X753 a_11439_4597# a_10499_4853# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X754 a_24234_14385# ui_in[0] a_24241_14651# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1274 pd=1.16667 as=0.10855 ps=1.36 w=0.42 l=0.15
**devattr s=4316,272 d=2268,138
X755 a_16297_2159# a_15119_1793# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X756 sky130_fd_sc_hd__inv_16_0.A sky130_fd_sc_hd__inv_12_0.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X757 sky130_fd_sc_hd__inv_8_0.A sky130_fd_sc_hd__inv_6_0.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X758 a_6281_11907# a_6003_11935# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X759 a_10955_11939# a_9715_11297# a_10869_11939# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X760 a_10471_5727# VGND a_10888_5837# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X761 VGND a_12194_5433# a_12142_5459# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X762 a_18553_4938# a_18371_4938# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X763 VGND sky130_fd_sc_hd__inv_16_0.A uo_out[0] VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X764 a_10160_4571# VDPWR a_10385_4597# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X765 VDPWR a_4905_12113# a_6003_11935# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X766 a_9501_13813# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X767 a_4847_14525# a_4513_14775# a_4763_14775# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X768 a_11147_11911# a_10869_11939# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X769 VGND a_13161_23139# a_13119_22871# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.07108 ps=0.80231 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X770 a_14982_22987# a_14814_23241# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14038 pd=1.37821 as=0.15033 ps=1.4282 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X771 VGND a_9896_1767# a_9844_1793# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X772 sky130_fd_sc_hd__dfxbp_1_9.Q a_18667_31977# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X773 a_4515_11543# VDPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X774 sky130_fd_sc_hd__inv_6_0.A sky130_fd_sc_hd__inv_4_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X775 VDPWR a_9715_11297# a_10841_12931# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0805 ps=0.94333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X776 a_17544_4529# VDPWR a_16793_4785# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X777 sky130_fd_sc_hd__dfxbp_1_8.Q_N a_18667_34839# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3880,195 d=6760,364
X778 VDPWR a_11888_1767# a_11836_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X779 a_14596_1793# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X780 a_16660_1793# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X781 VGND sky130_fd_sc_hd__inv_16_0.A uo_out[0] VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X782 sky130_fd_sc_hd__inv_2_0.A a_18667_34259# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X783 a_24241_14651# a_6208_2817# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.36 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X784 VGND sky130_fd_sc_hd__inv_8_0.A sky130_fd_sc_hd__inv_12_0.A VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X785 a_12993_23237# a_12129_22871# a_12736_22983# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.07862 ps=0.77179 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X786 VGND a_17689_23143# a_17647_22875# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.07108 ps=0.80231 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X787 a_12017_1793# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X788 VGND VDPWR a_6698_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X789 a_8262_22875# a_7863_22875# a_8136_23241# VGND sky130_fd_pr__special_nfet_01v8 ad=0.06425 pd=0.70615 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X790 a_12663_23237# a_12129_22871# a_12568_23237# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X791 VDPWR a_18667_34259# a_18667_34839# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.12828 pd=1.21873 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=6160,267
X792 a_9453_13111# VDPWR a_9371_13111# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X793 a_6021_13769# a_4903_15345# a_5933_13769# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X794 VDPWR a_1920_1765# a_1868_1791# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X795 a_18693_33761# a_18667_33731# a_18667_33966# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X796 a_14814_23241# a_14541_22875# a_14729_22875# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X797 a_11501_15239# a_10953_14739# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X798 VGND a_6238_6077# a_24152_14385# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.10855 ps=1.36 w=0.42 l=0.15
**devattr s=4316,272 d=2268,138
X799 a_6127_13769# a_4837_16089# a_6021_13769# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X800 uo_out[0] sky130_fd_sc_hd__inv_16_0.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X801 a_18693_33581# sky130_fd_sc_hd__dfxbp_1_8.Q_N VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=4368,272 d=2310,139
X802 VGND a_15407_23143# a_15838_23197# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=3880,195
X803 VDPWR VDPWR a_9621_13111# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X804 a_4627_12141# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X805 a_8377_5305# a_7315_5043# a_8794_5049# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X806 VDPWR sky130_fd_sc_hd__inv_6_0.A sky130_fd_sc_hd__inv_8_0.A VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X807 a_9713_14529# a_9379_14779# a_9629_14779# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X808 a_6429_5409# a_6375_5299# a_6036_5017# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X809 a_7944_1767# a_7221_1787# a_8169_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X810 a_18667_33966# a_18667_33636# a_18693_33581# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X811 VDPWR a_12736_22983# a_12663_23237# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X812 a_10887_13773# a_9769_15349# a_10799_13773# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X813 a_4746_1787# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X814 sky130_fd_sc_hd__dfxbp_1_0.Q_N a_9160_23197# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=6160,267 d=10400,504
X815 a_10761_14767# a_9715_11297# a_10675_14767# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X816 a_4637_10577# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X817 VDPWR a_6238_6077# a_2217_5025# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X818 VDPWR VDPWR a_12281_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X819 VGND VDPWR a_8337_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X820 a_13969_2159# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X821 sky130_fd_sc_hd__inv_8_0.A sky130_fd_sc_hd__inv_6_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X822 VGND a_18667_31552# a_19059_31529# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.07495 ps=0.82385 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X823 VGND ui_in[0] a_23731_14309# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X824 VDPWR a_19235_17155# a_18113_17153# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X825 a_6003_11935# a_4849_11293# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X826 VDPWR VDPWR a_4477_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X827 VDPWR VGND a_9034_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X828 a_12823_4919# a_12769_4809# a_12430_4527# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X829 VGND sky130_fd_sc_hd__inv_4_0.A sky130_fd_sc_hd__inv_6_0.A VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X830 a_7831_14003# a_4915_10549# a_7749_14003# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2772,150
X831 a_16486_16197# a_15641_17149# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X832 VGND VDPWR a_4721_13809# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X833 a_4423_5299# a_3229_5051# a_4840_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X834 a_4383_2153# a_3199_1791# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X835 a_10499_4853# VDPWR a_10916_4963# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X836 VGND a_8729_23143# a_8687_22875# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.07108 ps=0.80231 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X837 sky130_fd_sc_hd__inv_12_0.A sky130_fd_sc_hd__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X838 a_4309_5409# VDPWR a_4213_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X839 sky130_fd_sc_hd__inv_12_0.A sky130_fd_sc_hd__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X840 sky130_fd_sc_hd__inv_6_0.A sky130_fd_sc_hd__inv_4_0.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X841 VGND a_12993_23237# a_13161_23139# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X842 sky130_fd_sc_hd__dfxbp_1_5.CLK a_17689_23143# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X843 a_16485_5729# a_15431_5467# a_16902_5839# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X844 a_9223_1793# a_8283_2049# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X845 VDPWR VGND a_17544_4529# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X846 VDPWR sky130_fd_sc_hd__inv_2_0.A sky130_fd_sc_hd__inv_4_0.A VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X847 a_12281_1793# a_12227_2049# a_11888_1767# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X848 a_2343_5051# a_2217_5025# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X849 a_7927_14003# a_6281_11907# a_7831_14003# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X850 a_10289_4597# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X851 a_7173_15235# a_6635_15235# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X852 a_12039_15239# a_11501_15239# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X853 a_10525_5837# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X854 VDPWR a_13840_1767# a_13788_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X855 a_8283_2049# a_7221_1787# a_8700_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X856 a_14432_4521# a_13709_4553# a_14657_4547# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X857 a_24234_14385# a_24774_14701# a_24962_14701# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1274 pd=1.16667 as=0.09209 ps=0.99 w=0.42 l=0.15
**devattr s=3683,198 d=10752,424
X858 a_15365_22875# a_14375_22875# a_15239_23241# VGND sky130_fd_pr__special_nfet_01v8 ad=0.06092 pd=0.68769 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X859 a_14152_5441# a_13473_5459# a_14377_5833# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X860 a_2313_1791# a_2259_2047# a_1920_1765# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X861 a_17733_4529# a_16793_4785# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X862 a_9771_12117# a_9493_12145# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X863 VGND a_9771_12117# a_10955_11939# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X864 a_16454_4503# a_15711_4547# a_16679_4529# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X865 a_12694_22871# a_12295_22871# a_12568_23237# VGND sky130_fd_pr__special_nfet_01v8 ad=0.06425 pd=0.70615 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X866 a_9128_5415# VDPWR a_8377_5305# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X867 a_18689_27461# a_18663_26922# a_18663_27756# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X868 VGND a_17521_23241# a_17689_23143# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X869 a_11777_15239# a_10953_14739# a_11671_15239# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X870 a_17210_4529# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X871 a_15188_4547# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X872 VDPWR sky130_fd_sc_hd__inv_12_0.A sky130_fd_sc_hd__inv_16_0.A VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X873 VDPWR a_9705_12861# a_10717_13773# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X874 a_10357_5471# VDPWR a_10261_5471# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X875 VDPWR VDPWR a_12587_5459# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X876 a_11175_1793# a_10235_2049# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X877 VDPWR VGND a_10553_4597# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X878 a_9781_10553# a_9503_10581# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X879 a_14233_2159# a_14179_2049# a_13840_1767# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X880 a_16297_2159# a_16243_2049# a_15904_1767# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X881 a_13840_1767# a_13167_1793# a_14065_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X882 VGND sky130_fd_sc_hd__inv_12_0.A sky130_fd_sc_hd__inv_16_0.A VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X883 a_17605_23241# a_16823_22875# a_17521_23241# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X884 a_8193_13753# a_7749_14003# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4075,198 d=7020,368
X885 a_4755_12857# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X886 a_12978_2159# VDPWR a_12227_2049# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X887 VGND a_4515_11543# a_4849_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X888 a_6036_5017# a_5363_5043# a_6261_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X889 VDPWR a_9705_12861# a_10841_12931# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0805 ps=0.94333 w=0.42 l=0.15
**devattr s=2646,147 d=5689,267
X890 a_13709_4553# a_12769_4809# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X891 a_12559_4919# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X892 VDPWR a_3990_1761# a_3938_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X893 a_4585_16339# VDPWR a_4503_16339# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X894 a_12430_4527# a_11439_4597# a_12655_4553# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X895 a_18671_29306# a_18671_29438# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.12659 pd=1.2736 as=0.12379 ps=1.28732 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X896 a_10953_14739# a_10675_14767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X897 VDPWR a_7113_13395# a_7999_14003# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=5930,268
X898 VGND a_8038_5023# a_7986_5049# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X899 VDPWR VDPWR a_6429_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X900 a_7032_1787# VDPWR a_6281_2043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X901 VGND a_18667_25299# a_18667_25879# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=3880,195
X902 VDPWR VDPWR a_16297_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X903 sky130_fd_sc_hd__dfxbp_1_9.CLK a_18671_29731# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X904 a_10289_1793# a_9223_1793# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X905 sky130_fd_sc_hd__dfxbp_1_9.Q_N a_18667_32557# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=6160,267 d=10400,504
X906 VDPWR a_4839_12857# a_5809_14763# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X907 a_6335_2153# a_5269_1787# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X908 a_13077_23237# a_12295_22871# a_12993_23237# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3528,168
X909 a_4595_14775# VDPWR a_4513_14775# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X910 a_7999_14003# a_7173_15235# a_7927_14003# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X911 a_5269_1787# a_4329_2043# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X912 a_8073_2159# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X913 a_13186_4553# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X914 a_3990_1761# a_3199_1791# a_4215_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X915 a_8431_5049# a_7315_5043# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X916 VDPWR a_18671_29731# a_18671_30311# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.12828 pd=1.21873 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=6160,267
X917 a_18671_29108# a_18671_29203# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X918 VGND a_20109_17157# a_19235_17155# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X919 VGND a_8561_23241# a_8729_23143# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X920 a_12295_22871# a_12129_22871# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X921 VGND VGND a_8337_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X922 a_18846_5265# a_17733_4529# a_18625_4938# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
**devattr s=3990,179 d=2772,150
X923 a_6261_5409# VDPWR a_6165_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X924 a_2049_1791# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X925 a_2145_2157# VDPWR a_2049_2157# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X926 a_19059_34232# a_18667_33731# a_18667_34470# VGND sky130_fd_pr__special_nfet_01v8 ad=0.06092 pd=0.68769 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X927 a_18663_27756# a_18663_27017# a_18663_27120# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.07862 ps=0.77179 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X928 VDPWR sky130_fd_sc_hd__inv_16_0.A uo_out[0] VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X929 sky130_fd_sc_hd__inv_16_0.A sky130_fd_sc_hd__inv_12_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X930 a_4840_5409# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X931 VDPWR VGND a_4477_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X932 a_10807_23245# a_10109_22879# a_10550_22991# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.07121 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X933 sky130_fd_sc_hd__inv_16_0.A sky130_fd_sc_hd__inv_12_0.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X934 VDPWR VDPWR a_4383_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X935 VDPWR a_10975_23147# a_11406_23201# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.12828 pd=1.21873 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=6160,267
X936 a_6389_13769# a_5851_13769# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X937 a_4839_12857# a_4505_13107# a_4755_13107# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X938 VGND VDPWR a_16847_4895# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X939 a_10553_4963# VDPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X940 a_19510_16177# a_18742_16187# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X941 VGND a_4839_12857# a_6127_13769# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X942 VDPWR a_9769_15349# a_10717_13773# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X943 VGND VGND a_9128_5415# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X944 VDPWR a_17689_23143# a_18120_23197# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.12828 pd=1.21873 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=6160,267
X945 VGND a_18671_29942# a_18671_29731# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X946 a_14729_22875# sky130_fd_sc_hd__dfxbp_1_3.Q_N VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08755 pd=0.89385 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X947 a_16539_5839# a_15431_5467# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X948 a_12113_1793# VDPWR a_12017_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X949 a_3010_1791# VDPWR a_2259_2047# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X950 VGND a_9705_12861# a_10993_13773# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X951 VDPWR a_16454_4503# a_16402_4529# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X952 VDPWR a_14432_4521# a_14380_4547# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X953 a_14657_4913# VDPWR a_14561_4913# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X954 a_17425_5473# a_16485_5729# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X955 sky130_fd_sc_hd__dfxbp_1_4.Q_N a_18120_23197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3880,195 d=6760,364
X956 a_23511_14335# ui_in[0] a_23761_14335# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.09322 ps=1.07 w=0.42 l=0.15
**devattr s=3409,185 d=4368,272
X957 VDPWR VDPWR a_8700_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X958 a_4765_11293# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X959 VGND a_10132_5445# a_10080_5471# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X960 a_21506_16181# a_20384_16179# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X961 a_14930_2159# VDPWR a_14179_2049# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X962 a_16994_2159# VDPWR a_16243_2049# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X963 a_10235_2049# a_9223_1793# a_10652_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X964 VGND sky130_fd_sc_hd__inv_8_0.A sky130_fd_sc_hd__inv_12_0.A VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X965 VDPWR sky130_fd_sc_hd__dfxbp_1_7.Q a_18671_29203# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.12828 pd=1.21873 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X966 a_16583_4529# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X967 a_14561_4547# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X968 a_16371_5473# VDPWR a_16275_5473# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X969 a_4903_15345# a_4625_15373# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X970 VDPWR a_6036_5017# a_5984_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X971 a_19055_27097# a_18663_26922# a_18663_27252# VGND sky130_fd_pr__special_nfet_01v8 ad=0.06425 pd=0.70615 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X972 VDPWR VGND a_12587_5459# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X973 uo_out[0] sky130_fd_sc_hd__inv_16_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X974 a_14065_2159# VDPWR a_13969_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X975 a_16129_2159# VDPWR a_16033_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X976 VDPWR VGND a_14825_4547# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X977 uo_out[0] sky130_fd_sc_hd__inv_16_0.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X978 VGND a_11255_13773# a_11728_13649# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4010,197
X979 a_10382_23245# a_10109_22879# a_10297_22879# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X980 a_6165_5043# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X981 VGND VGND a_14545_5833# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X982 VGND a_10975_23147# a_11406_23201# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=3880,195
X983 a_2343_5051# a_2289_5307# a_1950_5025# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X984 a_16033_1793# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X985 a_6281_2043# a_5269_1787# a_6698_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X986 VDPWR a_12430_4527# a_12378_4553# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X987 a_18697_29053# sky130_fd_sc_hd__dfxbp_1_6.Q_N VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08755 pd=0.89385 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X988 a_7863_22875# a_7697_22875# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X989 VGND a_22365_17147# a_21491_17145# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X990 VDPWR VGND a_6429_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X991 VDPWR a_6389_13769# a_6944_13645# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5830,267
X992 VDPWR VGND a_16297_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X993 a_11250_4597# VDPWR a_10499_4853# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X994 VGND a_18667_34259# a_19059_34232# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.07108 ps=0.80231 w=0.42 l=0.15
**devattr s=2640,149 d=4368,272
X995 a_18667_24676# a_18667_24771# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X996 VDPWR a_12993_23237# a_13161_23139# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X997 VDPWR VDPWR a_6335_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X998 a_24407_14651# a_23731_14309# a_24234_14385# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.09013 pd=0.995 as=0.1274 ps=1.16667 w=0.42 l=0.15
**devattr s=2268,138 d=3605,199
X999 VGND a_4839_12857# a_6129_12927# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5266,228
X1000 a_2676_2157# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X1001 a_18667_25006# a_18667_24771# a_18693_24621# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.07505 ps=0.76615 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X1002 a_7863_22875# a_7697_22875# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.12828 ps=1.21873 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X1003 a_4119_1787# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X1004 a_18667_33834# a_18667_33966# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14038 pd=1.37821 as=0.15033 ps=1.4282 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X1005 a_9369_16343# VDPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X1006 VGND a_9703_16093# a_11777_15239# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X1007 VDPWR VGND a_12823_4553# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X1008 VGND sky130_fd_sc_hd__dfxbp_1_4.CLK a_16657_22875# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X1009 a_9703_16093# VDPWR a_9619_16093# VGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X1010 VGND a_9705_12861# a_10995_12931# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5266,228
X1011 VDPWR a_16471_17161# a_15693_17123# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X1012 VDPWR a_18667_25299# a_18693_25215# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X1013 VDPWR sky130_fd_sc_hd__dfxbp_1_7.CLK a_18663_27017# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.12828 pd=1.21873 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X1014 a_10289_1793# a_10235_2049# a_9896_1767# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X1015 VDPWR VDPWR a_14908_5467# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X1016 sky130_fd_sc_hd__dfxbp_1_7.Q a_18663_27545# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X1017 sky130_fd_sc_hd__dfxbp_1_1.CLK a_8729_23143# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X1018 VDPWR a_17521_23241# a_17689_23143# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X1019 a_10841_12931# a_9779_13785# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0805 pd=0.94333 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2646,147
X1020 VDPWR VGND a_4383_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X1021 a_14491_5723# a_13473_5459# a_14908_5467# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X1022 VGND a_8304_22987# a_8262_22875# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.07495 ps=0.82385 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X1023 sky130_fd_sc_hd__dfxbp_1_3.Q_N a_15838_23197# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=6160,267 d=10400,504
X1024 VDPWR sky130_fd_sc_hd__dfxbp_1_4.CLK a_16657_22875# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.12828 pd=1.21873 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X1025 a_12644_1793# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X1026 VDPWR a_9317_5049# a_18371_4938# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2772,150
X1027 a_15239_23241# a_14541_22875# a_14982_22987# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.07121 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X1028 a_18742_16187# a_18128_16189# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X1029 a_6335_2153# a_6281_2043# a_5942_1761# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X1030 VGND VDPWR a_9579_12145# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X1031 a_6329_12927# a_5975_12927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=5266,228 d=6760,364
X1032 VGND VDPWR a_4477_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X1033 VGND VDPWR a_12950_5825# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X1034 VGND sky130_fd_sc_hd__dfxbp_1_5.CLK a_18667_24771# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X1035 a_5174_5043# VDPWR a_4423_5299# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X1036 VGND VDPWR a_15188_4913# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X1037 a_8431_5049# a_8377_5305# a_8038_5023# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X1038 a_11583_15239# a_8193_13753# a_11501_15239# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
X1039 a_11728_13649# a_11195_12931# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X1040 a_12587_5825# a_11411_5471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X1041 a_18663_27252# a_18663_26922# a_18689_26867# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
**devattr s=2310,139 d=2730,149
X1042 VGND VDPWR a_9589_10581# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X1043 a_19059_33811# a_18667_33636# a_18667_33966# VGND sky130_fd_pr__special_nfet_01v8 ad=0.06425 pd=0.70615 as=0.0621 ps=0.705 w=0.36 l=0.15
**devattr s=2484,141 d=2784,153
X1044 a_17236_5473# VDPWR a_16485_5729# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X1045 a_23133_17137# a_22274_16171# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X1046 a_11979_13399# a_11728_13649# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4010,197 d=6760,364
X1047 VDPWR VGND a_9453_13111# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X1048 a_18667_33636# a_18667_33731# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.12828 ps=1.21873 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X1049 VGND sky130_fd_sc_hd__dfxbp_1_0.CLK a_7697_22875# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X1050 a_24318_14385# a_6208_2817# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10858 pd=1.36 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X1051 a_10717_13773# a_9715_11297# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X1052 a_10923_12931# a_9715_11297# a_10841_12931# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X1053 a_14596_2159# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X1054 VGND a_15904_1767# a_15852_1793# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X1055 a_16660_2159# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X1056 a_17264_22987# a_17096_23241# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14038 pd=1.37821 as=0.15033 ps=1.4282 w=0.75 l=0.15
**devattr s=7155,252 d=4380,215
X1057 VDPWR VDPWR a_4627_12141# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X1058 a_6281_11907# a_6003_11935# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X1059 a_18667_34470# a_18667_33731# a_18667_33834# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.07862 ps=0.77179 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X1060 a_18663_27120# a_18663_27252# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.12659 pd=1.2736 as=0.12379 ps=1.28732 w=0.64 l=0.15
**devattr s=4838,217 d=3956,199
X1061 VDPWR a_8561_23241# a_8729_23143# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X1062 VGND a_9705_12861# a_10761_14767# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X1063 a_4915_10549# a_4637_10577# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X1064 a_2343_5417# a_2217_5025# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X1065 VGND VDPWR a_8794_5415# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X1066 VDPWR VGND a_11250_4597# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X1067 sky130_fd_sc_hd__inv_16_0.A sky130_fd_sc_hd__inv_12_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X1068 a_24318_14385# a_23731_14309# a_24234_14385# VGND sky130_fd_pr__nfet_01v8 ad=0.10858 pd=1.36 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=4318,272
X1069 a_12615_14007# a_9781_10553# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4368,272 d=2772,150
X1070 a_11147_11911# a_10869_11939# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X1071 a_3229_5051# a_2289_5307# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X1072 VDPWR sky130_fd_sc_hd__inv_16_0.A uo_out[0] VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X1073 VDPWR a_10975_23147# a_10891_23245# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X1074 a_6087_14735# a_5809_14763# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X1075 VDPWR VDPWR a_4637_10577# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X1076 a_10553_4963# a_10499_4853# a_10160_4571# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X1077 VDPWR a_18663_27756# a_18663_27545# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X1078 VDPWR sky130_fd_sc_hd__dfxbp_1_0.CLK a_7697_22875# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.12828 pd=1.21873 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X1079 a_12017_2159# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X1080 VDPWR VGND a_14930_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X1081 sky130_fd_sc_hd__dfxbp_1_7.Q_N a_18663_28125# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3880,195 d=6760,364
X1082 a_4753_16339# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X1083 a_9619_16093# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X1084 VGND VGND a_8431_5415# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X1085 VGND a_18667_31977# a_18667_32557# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=3880,195
X1086 a_2175_5051# VDPWR a_2079_5051# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X1087 a_6071_1787# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X1088 a_4763_14775# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X1089 a_10357_5837# VDPWR a_10261_5837# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X1090 a_13284_5459# VDPWR a_12533_5715# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X1091 a_10916_4597# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X1092 VDPWR VGND a_6335_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X1093 a_15522_4547# VDPWR a_14771_4803# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X1094 sky130_fd_sc_hd__dfxbp_1_3.CLK a_13161_23139# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X1095 a_18128_16189# a_17254_16187# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X1096 a_10525_5471# a_10471_5727# a_10132_5445# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X1097 VDPWR VDPWR a_10553_4597# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X1098 VGND VDPWR a_12281_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X1099 VDPWR sky130_fd_sc_hd__inv_8_0.A sky130_fd_sc_hd__inv_12_0.A VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X1100 a_8561_23241# a_7697_22875# a_8304_22987# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.07862 ps=0.77179 w=0.42 l=0.15
**devattr s=4380,215 d=2268,138
X1101 VGND a_12736_22983# a_12694_22871# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.07495 ps=0.82385 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X1102 a_6036_5017# a_5363_5043# a_6261_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X1103 a_15242_5833# VDPWR a_14491_5723# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X1104 a_8231_23241# a_7697_22875# a_8136_23241# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
**devattr s=2730,149 d=3066,157
X1105 VDPWR sky130_fd_sc_hd__dfxbp_1_9.Q a_18667_33731# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.12828 pd=1.21873 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X1106 a_10995_12931# a_9779_13785# a_10923_12931# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=1764,126
X1107 a_9579_12145# VGND a_9493_12145# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X1108 a_9381_11547# VDPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X1109 a_10986_1793# VDPWR a_10235_2049# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X1110 VDPWR VGND a_12978_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X1111 VGND VGND a_9034_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X1112 a_12430_4527# a_11439_4597# a_12655_4919# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X1113 VDPWR a_18113_17153# a_17345_17163# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X1114 VGND VDPWR a_6429_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X1115 a_7126_5043# VDPWR a_6375_5299# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X1116 a_9715_11297# VDPWR a_9631_11297# VGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X1117 VDPWR sky130_fd_sc_hd__inv_12_0.A sky130_fd_sc_hd__inv_16_0.A VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X1118 a_9589_10581# VGND a_9503_10581# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X1119 VDPWR VGND a_5174_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X1120 uo_out[0] sky130_fd_sc_hd__inv_16_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X1121 uo_out[0] sky130_fd_sc_hd__inv_16_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X1122 VDPWR a_8304_22987# a_8231_23241# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X1123 a_18693_31299# sky130_fd_sc_hd__dfxbp_1_9.Q_N VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08755 pd=0.89385 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X1124 VGND sky130_fd_sc_hd__inv_12_0.A sky130_fd_sc_hd__inv_16_0.A VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X1125 a_13167_1793# a_12227_2049# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X1126 a_13186_4919# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X1127 a_18663_27756# a_18663_26922# a_18663_27120# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.07121 ps=0.7164 w=0.36 l=0.15
**devattr s=3956,199 d=2736,148
X1128 a_10297_22879# sky130_fd_sc_hd__dfxbp_1_1.Q_N VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08755 pd=0.89385 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4368,272 d=3252,166
X1129 a_9317_5049# a_8377_5305# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X1130 a_14545_5467# a_13473_5459# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X1131 a_12281_2159# a_12227_2049# a_11888_1767# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X1132 a_11888_1767# a_11175_1793# a_12113_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X1133 a_13520_4553# VDPWR a_12769_4809# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X1134 a_10799_13773# a_9715_11297# a_10717_13773# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
X1135 a_5363_5043# a_4423_5299# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X1136 a_6167_2153# VDPWR a_6071_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X1137 sky130_fd_sc_hd__inv_16_0.A sky130_fd_sc_hd__inv_12_0.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X1138 a_4839_12857# VDPWR a_4755_12857# VGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X1139 a_4084_5017# a_3229_5051# a_4309_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X1140 a_8283_2049# a_7221_1787# a_8700_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X1141 a_3199_1791# a_2259_2047# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X1142 VGND VGND a_4477_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X1143 VDPWR a_18667_31977# a_18693_31893# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X1144 VDPWR a_18671_29306# a_18697_29233# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X1145 a_2313_2157# a_2259_2047# a_1920_1765# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X1146 a_8263_5049# VDPWR a_8167_5049# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X1147 VDPWR a_21491_17145# a_20877_17147# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X1148 VDPWR ui_in[0] a_23731_14309# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.1083 ps=1.36 w=0.42 l=0.15
**devattr s=4332,272 d=4316,272
X1149 a_1920_1765# a_2187_1765# a_2145_1791# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X1150 uo_out[0] sky130_fd_sc_hd__inv_16_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X1151 VDPWR a_18667_24874# a_18693_24801# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7155,252
X1152 VDPWR VGND a_4585_16339# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X1153 a_5080_1787# VDPWR a_4329_2043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X1154 a_16146_5447# a_15431_5467# a_16371_5473# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X1155 sky130_fd_sc_hd__inv_12_0.A sky130_fd_sc_hd__inv_8_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X1156 sky130_fd_sc_hd__inv_2_0.A a_18667_34259# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=6760,364
X1157 VGND a_9369_16343# a_9703_16093# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X1158 a_16902_5473# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X1159 sky130_fd_sc_hd__inv_12_0.A sky130_fd_sc_hd__inv_8_0.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X1160 VDPWR VGND a_4595_14775# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X1161 a_13840_1767# a_13167_1793# a_14065_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X1162 VDPWR VDPWR a_16539_5473# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X1163 a_19055_27518# a_18663_27017# a_18663_27756# VGND sky130_fd_pr__special_nfet_01v8 ad=0.06092 pd=0.68769 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X1164 VGND a_5942_1761# a_5890_1787# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X1165 a_16847_4895# a_16793_4785# a_16454_4503# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X1166 VDPWR VGND a_13284_5459# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X1167 VDPWR VDPWR a_2313_1791# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X1168 a_9621_12861# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X1169 VDPWR VGND a_15522_4547# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X1170 VDPWR sky130_fd_sc_hd__inv_16_0.A uo_out[0] VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X1171 a_2706_5051# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X1172 a_12587_5825# a_12533_5715# a_12194_5433# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X1173 VDPWR a_10160_4571# a_10108_4597# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X1174 a_10385_4963# VDPWR a_10289_4963# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X1175 a_17254_16187# a_16486_16197# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X1176 VDPWR a_9713_14529# a_11501_15239# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X1177 VGND VGND a_15242_5833# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X1178 a_14825_4913# a_14771_4803# a_14432_4521# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X1179 VGND sky130_fd_sc_hd__inv_16_0.A uo_out[0] VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X1180 a_9556_17271# a_12615_14007# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5930,268 d=10800,508
X1181 sky130_fd_sc_hd__dfxbp_1_1.CLK a_8729_23143# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X1182 a_6635_15235# a_6087_14735# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X1183 VGND VDPWR a_16297_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X1184 sky130_fd_sc_hd__dfxbp_1_2.Q_N a_13592_23193# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=3880,195 d=6760,364
X1185 VDPWR a_20877_17147# a_20109_17157# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X1186 a_9703_16093# a_9369_16343# a_9619_16343# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X1187 a_13473_5459# a_12533_5715# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X1188 a_16371_5839# VDPWR a_16275_5839# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X1189 a_10289_2159# a_9223_1793# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X1190 VDPWR a_13161_23139# a_13077_23237# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X1191 a_14814_23241# a_14375_22875# a_14729_22875# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.07505 ps=0.76615 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X1192 a_23761_14335# a_23731_14309# a_23511_14701# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X1193 a_18839_4938# a_17425_5473# a_18625_4938# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
**devattr s=7728,268 d=3066,157
X1194 a_15711_4547# a_14771_4803# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X1195 VDPWR VDPWR a_10916_4597# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X1196 VGND a_18663_27120# a_19055_27097# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.07495 ps=0.82385 w=0.42 l=0.15
**devattr s=2784,153 d=4838,217
X1197 a_10933_22879# a_9943_22879# a_10807_23245# VGND sky130_fd_pr__special_nfet_01v8 ad=0.06092 pd=0.68769 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2640,149
X1198 VDPWR a_15407_23143# a_15323_23241# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0882 ps=0.84 w=0.42 l=0.15
**devattr s=3528,168 d=4452,274
X1199 VDPWR VGND a_7126_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X1200 a_12194_5433# a_11411_5471# a_12419_5459# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X1201 VGND sky130_fd_sc_hd__inv_6_0.A sky130_fd_sc_hd__inv_8_0.A VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X1202 VDPWR VGND a_16994_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X1203 a_12950_5459# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X1204 a_11411_5471# a_10471_5727# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X1205 a_15119_1793# a_14179_2049# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X1206 a_24962_14701# ui_in[1] a_23761_14335# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.09209 pd=0.99 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=3683,198
X1207 a_8337_1793# a_8283_2049# a_7944_1767# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X1208 a_6165_5409# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X1209 a_7315_5043# a_6375_5299# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X1210 a_14908_5833# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X1211 a_2049_2157# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X1212 VGND sky130_fd_sc_hd__dfxbp_1_1.CLK a_9943_22879# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X1213 a_2343_5417# a_2289_5307# a_1950_5025# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X1214 a_6208_2817# a_16243_2049# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X1215 VDPWR VGND a_13520_4553# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X1216 VGND a_18667_32188# a_18667_31977# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X1217 VGND a_11147_11911# a_12615_14007# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2772,150 d=2268,138
X1218 VGND VDPWR a_14545_5833# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X1219 a_10652_1793# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X1220 a_14179_2049# a_13167_1793# a_14596_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X1221 VDPWR sky130_fd_sc_hd__inv_4_0.A sky130_fd_sc_hd__inv_6_0.A VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X1222 VGND a_6208_2817# a_2187_1765# VGND sky130_fd_pr__nfet_01v8 ad=0.12573 pd=1.30744 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X1223 sky130_fd_sc_hd__dfxbp_1_1.Q_N a_11406_23201# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=6160,267 d=10400,504
X1224 VGND VGND a_6429_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X1225 a_15904_1767# a_15119_1793# a_16129_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X1226 a_11439_4597# a_10499_4853# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X1227 a_4849_11293# VDPWR a_4765_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X1228 uo_out[0] sky130_fd_sc_hd__inv_16_0.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X1229 VDPWR a_18667_34470# a_18667_34259# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.27 ps=2.54 w=1 l=0.15
**devattr s=10800,508 d=5400,254
X1230 VDPWR sky130_fd_sc_hd__dfxbp_1_1.CLK a_9943_22879# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.12828 pd=1.21873 as=0.1664 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X1231 VDPWR a_4084_5017# a_4032_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X1232 VDPWR VDPWR a_14233_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X1233 VDPWR VGND a_5080_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X1234 a_6698_2153# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08124 ps=0.84481 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X1235 a_12113_2159# VDPWR a_12017_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X1236 a_3010_2157# VDPWR a_2259_2047# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X1237 VGND VGND a_12823_4919# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X1238 a_8794_5049# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X1239 a_7173_15235# a_6635_15235# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X1240 VDPWR a_16146_5447# a_16094_5473# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X1241 a_5851_13769# a_4837_16089# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X1242 a_4849_11293# a_4515_11543# a_4765_11543# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X1243 VGND a_4905_12113# a_6089_11935# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X1244 VGND VDPWR a_8700_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08124 pd=0.84481 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X1245 VDPWR a_23133_17137# a_22365_17147# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X1246 a_4213_5043# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X1247 a_4329_2043# a_3199_1791# a_4746_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X1248 sky130_fd_sc_hd__inv_8_0.A sky130_fd_sc_hd__inv_6_0.A VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.20043 ps=1.90427 w=1 l=0.15
**devattr s=17200,572 d=5400,254
X1249 a_9461_14779# VDPWR a_9379_14779# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X1250 a_20384_16179# a_19510_16177# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12573 ps=1.30744 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X1251 a_6911_15235# a_6087_14735# a_6805_15235# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X1252 VDPWR a_4839_12857# a_5851_13769# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X1253 a_16275_5473# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08418 ps=0.79979 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X1254 a_10382_23245# a_9943_22879# a_10297_22879# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.07505 ps=0.76615 w=0.36 l=0.15
**devattr s=3252,166 d=2484,141
X1255 VDPWR VDPWR a_9629_14779# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X1256 VDPWR a_1950_5025# a_1898_5051# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20043 pd=1.90427 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X1257 VDPWR VDPWR a_2676_1791# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08418 pd=0.79979 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
C0 a_10132_5445# a_10471_5727# 0.04737f
C1 a_15119_1793# a_6208_2817# 0.00767f
C2 a_17733_4529# a_18625_4938# 0.19558f
C3 a_18663_28125# a_18671_29108# 0
C4 a_5942_1761# a_6167_2153# 0.00559f
C5 a_4913_13781# a_4635_13809# 0.1205f
C6 a_11222_5471# a_10471_5727# 0.00682f
C7 a_10916_4963# VDPWR 0.05811f
C8 a_18667_32557# a_18667_31977# 0.10805f
C9 a_7113_13395# a_4849_11293# 0.00118f
C10 a_24241_14651# sky130_fd_sc_hd__dfxbp_1_0.CLK 0
C11 a_7113_13395# a_5851_13769# 0
C12 a_13167_1793# a_13969_1793# 0
C13 a_10717_13773# a_9705_12861# 0.13054f
C14 a_9705_12861# a_10887_13773# 0
C15 a_4753_16339# a_4837_16089# 0.07445f
C16 a_16454_4503# a_16793_4785# 0.04737f
C17 a_7697_22875# a_8231_23241# 0.0027f
C18 a_16679_4895# a_16847_4895# 0
C19 a_10160_4571# a_10553_4963# 0.02301f
C20 a_11810_13649# a_9715_11297# 0
C21 a_8304_22987# a_8729_23143# 0
C22 a_4383_1787# a_4215_1787# 0
C23 a_6281_11907# a_7831_14003# 0.00377f
C24 a_9371_13111# a_9779_13785# 0
C25 a_10841_12931# a_9771_12117# 0
C26 a_7944_1767# a_8169_2159# 0.00559f
C27 a_23731_14309# a_6238_6077# 0.106f
C28 a_15188_4547# a_14825_4547# 0.00985f
C29 a_10953_14739# a_9705_12861# 0.02465f
C30 a_10357_5471# a_10471_5727# 0
C31 a_12697_14007# a_11147_11911# 0.00377f
C32 a_2259_2047# a_2145_1791# 0
C33 a_4477_5043# a_4213_5043# 0
C34 a_5269_1787# a_6335_2153# 0.04534f
C35 a_6089_11935# a_4915_10549# 0
C36 VDPWR a_18697_29233# 0.00347f
C37 a_15431_5467# a_13473_5459# 0
C38 a_10499_4853# a_10916_4597# 0.03016f
C39 VDPWR a_8645_23241# 0.00627f
C40 a_4084_5017# a_3229_5051# 0.11874f
C41 a_15365_22875# VDPWR 0
C42 a_4837_16089# a_4913_13781# 0.01745f
C43 a_8283_2049# a_8337_2159# 0.03622f
C44 a_9317_5049# a_16793_4785# 0
C45 a_2187_1765# a_2049_2157# 0
C46 a_18671_29438# sky130_fd_sc_hd__dfxbp_1_7.Q_N 0
C47 a_17425_5473# VDPWR 0.27512f
C48 a_4763_14525# a_4903_15345# 0
C49 a_9769_15349# a_10993_13773# 0
C50 a_17733_4529# a_17544_4895# 0
C51 a_6238_6077# a_10888_5471# 0
C52 a_12323_5459# a_12194_5433# 0.00758f
C53 VDPWR a_10993_13773# 0.0014f
C54 a_8136_23241# a_8262_22875# 0.00553f
C55 a_9703_16093# a_9771_12117# 0
C56 a_14596_2159# a_13167_1793# 0.03325f
C57 a_10652_1793# a_11175_1793# 0
C58 a_5895_14763# a_5809_14763# 0.00658f
C59 a_14545_5467# a_14281_5467# 0
C60 a_18663_27017# a_18667_24676# 0
C61 a_7221_1787# a_8169_1793# 0
C62 a_16539_5839# a_14491_5723# 0
C63 a_16454_4503# a_16847_4895# 0.02301f
C64 a_16679_4895# a_6238_6077# 0
C65 a_6911_15235# a_4837_16089# 0.00241f
C66 sky130_fd_sc_hd__dfxbp_1_6.Q_N sky130_fd_sc_hd__dfxbp_1_7.Q_N 0
C67 a_1950_5025# a_2217_5025# 0.08244f
C68 a_9371_13111# a_9621_12861# 0.00723f
C69 a_18667_25006# a_18667_24874# 0.23675f
C70 a_18671_29942# a_18671_29108# 0.19462f
C71 sky130_fd_sc_hd__dfxbp_1_8.Q_N a_18667_33834# 0.05782f
C72 a_18693_33581# a_18667_33834# 0
C73 a_19059_24851# sky130_fd_sc_hd__dfxbp_1_7.CLK 0
C74 a_16485_5729# a_16371_5839# 0
C75 a_8377_5305# a_8431_5415# 0.03622f
C76 a_9317_5049# a_14152_5441# 0
C77 a_4585_16339# a_4503_16339# 0.00641f
C78 sky130_fd_sc_hd__dfxbp_1_3.CLK a_13161_23139# 0.12322f
C79 a_14179_2049# a_14233_1793# 0.00386f
C80 a_4849_11293# a_6862_13645# 0
C81 a_6862_13645# a_5851_13769# 0
C82 a_10235_2049# VDPWR 0.45025f
C83 a_9317_5049# a_16847_4895# 0
C84 a_6208_2817# a_14657_4547# 0
C85 a_8700_1793# VDPWR 0.21795f
C86 a_15407_23143# a_15838_23197# 0.10805f
C87 a_9317_5049# a_12533_5715# 0
C88 a_14814_23241# sky130_fd_sc_hd__dfxbp_1_2.Q_N 0
C89 a_9369_16343# a_9619_16093# 0.00723f
C90 a_18128_16189# a_16486_16197# 0
C91 a_2706_5051# VDPWR 0.21783f
C92 a_23677_14701# a_9556_17271# 0
C93 a_16793_4785# a_16847_4895# 0.03622f
C94 sky130_fd_sc_hd__dfxbp_1_7.Q_N a_18663_27252# 0.04247f
C95 a_2343_5417# a_2079_5417# 0
C96 a_16454_4503# a_6238_6077# 0
C97 VDPWR a_18671_29108# 0.31436f
C98 a_17264_22987# a_16823_22875# 0.11299f
C99 a_17191_23241# a_17096_23241# 0.00772f
C100 a_4477_5043# a_2217_5025# 0
C101 a_7113_13395# a_6635_15235# 0
C102 uo_out[2] uo_out[3] 0.03102f
C103 a_6238_6077# a_23677_14335# 0
C104 a_5269_1787# a_4746_1787# 0
C105 a_9621_13111# a_9371_13111# 0.02504f
C106 a_9453_13111# a_4915_10549# 0
C107 a_9493_12145# a_9501_13813# 0
C108 a_17689_23143# a_17264_22987# 0
C109 a_15431_5467# a_14491_5723# 0.13739f
C110 VDPWR a_11836_1793# 0.16681f
C111 a_10975_23147# a_9943_22879# 0.04808f
C112 sky130_fd_sc_hd__dfxbp_1_9.CLK a_18671_29942# 0.0039f
C113 a_9317_5049# a_6238_6077# 0.0245f
C114 a_9705_12861# a_11195_12931# 0.08252f
C115 a_4839_12857# a_5933_13769# 0
C116 sky130_fd_sc_hd__dfxbp_1_1.Q_N sky130_fd_sc_hd__dfxbp_1_1.CLK 0.0174f
C117 a_14380_4547# VDPWR 0.16838f
C118 a_9713_14529# a_10675_14767# 0.00524f
C119 a_18689_27461# sky130_fd_sc_hd__dfxbp_1_7.Q_N 0
C120 a_9713_14529# a_9379_14779# 0.1679f
C121 a_20384_16179# VDPWR 0.45257f
C122 a_9629_14529# a_4915_10549# 0
C123 a_14825_4913# VDPWR 0.01165f
C124 a_16793_4785# a_6238_6077# 0
C125 a_16402_4529# a_16583_4895# 0
C126 a_10717_13773# a_9769_15349# 0.16757f
C127 a_9769_15349# a_10887_13773# 0.00818f
C128 a_14152_5441# a_12533_5715# 0.00359f
C129 a_16471_17161# a_17345_17163# 0.1036f
C130 a_15711_4547# a_16902_5839# 0
C131 VDPWR a_10887_13773# 0
C132 a_9781_10553# a_9503_10581# 0.1296f
C133 a_10717_13773# VDPWR 0.44659f
C134 sky130_fd_sc_hd__dfxbp_1_9.CLK a_19063_29704# 0
C135 a_10499_4853# a_11250_4597# 0.00682f
C136 a_4905_12113# a_4913_13781# 0.00627f
C137 a_7173_15235# a_5809_14763# 0
C138 a_6238_6077# a_12823_4919# 0
C139 a_10953_14739# a_9769_15349# 0
C140 a_10499_4853# a_12559_4919# 0
C141 a_4721_13809# a_4913_13781# 0.00222f
C142 a_10953_14739# VDPWR 0.62612f
C143 a_18667_31552# VDPWR 0.19117f
C144 a_18671_29203# a_18697_29233# 0.0027f
C145 sky130_fd_sc_hd__dfxbp_1_9.CLK VDPWR 0.27403f
C146 a_12430_4527# VDPWR 0.36701f
C147 a_6127_13769# VDPWR 0.0014f
C148 a_9943_22879# a_12483_22871# 0
C149 a_7863_22875# a_8729_23143# 0.03136f
C150 a_12559_4553# VDPWR 0.00126f
C151 a_9713_14529# a_8193_13753# 0.30236f
C152 a_11411_5471# a_10471_5727# 0.13964f
C153 a_14545_5833# a_13473_5459# 0.04534f
C154 sky130_fd_sc_hd__dfxbp_1_8.Q_N VDPWR 0.60759f
C155 a_9943_22879# VDPWR 0.66221f
C156 a_6635_15235# a_6862_13645# 0
C157 a_18693_33581# VDPWR 0.07701f
C158 a_6238_6077# a_14152_5441# 0.0052f
C159 a_6208_2817# a_10289_2159# 0
C160 sky130_fd_sc_hd__dfxbp_1_1.Q_N a_10807_23245# 0.09273f
C161 a_7927_14003# a_6281_11907# 0.00264f
C162 sky130_fd_sc_hd__dfxbp_1_7.CLK a_18663_26922# 0.01405f
C163 a_24234_14385# a_23761_14335# 0.22643f
C164 a_16823_22875# sky130_fd_sc_hd__dfxbp_1_3.Q_N 0.00105f
C165 a_6208_2817# a_14233_1793# 0
C166 a_16847_4895# a_6238_6077# 0
C167 a_17425_5473# a_9317_5049# 0.24941f
C168 a_9943_22879# a_9160_23197# 0
C169 a_14179_2049# a_14065_2159# 0
C170 a_18667_31552# sky130_fd_sc_hd__dfxbp_1_9.Q 0
C171 a_4837_16089# a_5933_13769# 0
C172 a_12793_14007# VDPWR 0
C173 a_11671_15239# a_9713_14529# 0.00624f
C174 a_12950_5459# VDPWR 0.21528f
C175 sky130_fd_sc_hd__dfxbp_1_9.Q sky130_fd_sc_hd__dfxbp_1_9.CLK 0.00137f
C176 a_18693_25215# VDPWR 0.00627f
C177 a_6238_6077# a_12533_5715# 0.00752f
C178 a_15711_4547# a_16485_5729# 0
C179 a_9713_14529# a_9779_13785# 0.0012f
C180 a_10385_4963# a_6238_6077# 0
C181 a_18667_24874# a_18667_25299# 0
C182 a_23761_14335# a_24318_14385# 0.04391f
C183 a_17264_22987# a_17011_22875# 0
C184 a_4753_16339# a_4625_15373# 0
C185 a_17425_5473# a_16793_4785# 0
C186 sky130_fd_sc_hd__dfxbp_1_7.Q a_18671_29306# 0
C187 sky130_fd_sc_hd__dfxbp_1_8.Q_N sky130_fd_sc_hd__dfxbp_1_9.Q 0.01744f
C188 a_2259_2047# a_2676_1791# 0.03016f
C189 a_12950_5825# VDPWR 0.01932f
C190 a_18693_33581# sky130_fd_sc_hd__dfxbp_1_9.Q 0
C191 a_10382_23245# a_10109_22879# 0.07715f
C192 a_10869_11939# a_9779_13785# 0
C193 a_8794_5415# a_8431_5415# 0.00847f
C194 a_5851_13769# a_4913_13781# 0.00386f
C195 a_2289_5307# VDPWR 0.44913f
C196 a_4849_11293# a_4913_13781# 0.26133f
C197 a_18667_31552# a_18667_31977# 0
C198 a_18693_24621# VDPWR 0.07699f
C199 sky130_fd_sc_hd__dfxbp_1_9.CLK a_18667_31977# 0
C200 a_7113_13395# a_9501_13813# 0
C201 a_10652_2159# VDPWR 0.02101f
C202 a_8431_5415# a_8263_5415# 0
C203 a_14561_4547# a_14825_4547# 0
C204 a_10289_4963# a_6238_6077# 0
C205 a_12823_4553# a_12769_4809# 0.00386f
C206 ui_in[1] VDPWR 0.28112f
C207 a_2175_5051# VDPWR 0.00105f
C208 a_17191_23241# VDPWR 0.00345f
C209 VDPWR a_14233_2159# 0.00967f
C210 a_18671_29108# a_18671_29203# 0.96835f
C211 a_6281_11907# a_7999_14003# 0
C212 sky130_fd_sc_hd__dfxbp_1_8.Q_N a_18667_31977# 0
C213 a_9556_17271# a_22274_16171# 0
C214 a_13473_5459# VDPWR 1.37069f
C215 a_11147_11911# a_9493_12145# 0
C216 a_15188_4547# VDPWR 0.22144f
C217 a_2259_2047# a_2187_1765# 0.25757f
C218 a_8431_5415# VDPWR 0.00982f
C219 a_16297_1793# a_16660_1793# 0.00985f
C220 sky130_fd_sc_hd__dfxbp_1_4.CLK a_17264_22987# 0
C221 a_18742_16187# a_18113_17153# 0.00293f
C222 a_6329_12927# a_6281_11907# 0.00298f
C223 a_12281_2159# a_12017_2159# 0
C224 a_12823_4553# a_13186_4553# 0.00985f
C225 a_6208_2817# a_8169_2159# 0
C226 a_12323_5825# a_12587_5825# 0
C227 a_9715_11297# a_10993_13773# 0
C228 a_9493_12145# a_9771_12117# 0.12057f
C229 a_14825_4547# a_12769_4809# 0
C230 a_6238_6077# a_10916_4963# 0
C231 a_18667_33636# a_18667_33731# 0.96835f
C232 a_14545_5833# a_14491_5723# 0.03622f
C233 a_11195_12931# VDPWR 0.31272f
C234 a_16454_4503# a_14825_4913# 0
C235 a_11501_15239# a_11728_13649# 0
C236 a_18697_29647# a_18671_29306# 0
C237 a_12587_5825# a_12419_5825# 0
C238 a_23731_14309# ui_in[1] 0
C239 a_18693_31479# a_18693_31299# 0.00123f
C240 rst_n ui_in[0] 0.03102f
C241 a_8136_23241# sky130_fd_sc_hd__dfxbp_1_0.CLK 0
C242 a_23761_14335# a_24241_14651# 0
C243 a_2187_1765# a_2313_2157# 0.05199f
C244 a_17254_16187# a_18113_17153# 0
C245 sky130_fd_sc_hd__dfxbp_1_2.CLK sky130_fd_sc_hd__dfxbp_1_1.CLK 0.00137f
C246 a_17011_22875# sky130_fd_sc_hd__dfxbp_1_3.Q_N 0
C247 a_4585_16339# a_4837_16089# 0
C248 a_11439_4597# a_12378_4553# 0.04732f
C249 a_9629_14779# a_9501_13813# 0
C250 sky130_fd_sc_hd__dfxbp_1_9.CLK a_18671_29203# 0
C251 a_17521_23241# sky130_fd_sc_hd__dfxbp_1_4.Q_N 0.09273f
C252 a_17425_5473# a_6238_6077# 0.00921f
C253 a_17210_4529# a_14771_4803# 0
C254 a_9705_12861# a_10841_12931# 0.29952f
C255 a_4423_5299# a_4840_5043# 0.03016f
C256 a_6208_2817# a_14065_2159# 0
C257 a_4840_5043# VDPWR 0.21797f
C258 a_4503_16339# a_4903_15345# 0
C259 a_11222_5837# a_10471_5727# 0.00696f
C260 a_1920_1765# VDPWR 0.36056f
C261 uio_in[2] uio_in[3] 0.03102f
C262 a_10923_12931# a_10841_12931# 0.00517f
C263 a_1950_5025# a_2343_5051# 0.02283f
C264 ui_in[0] a_24962_14701# 0.02483f
C265 a_8337_1793# VDPWR 0.18609f
C266 a_15852_1793# VDPWR 0.16666f
C267 a_9379_14779# a_9491_15377# 0
C268 a_24407_14651# a_24774_14701# 0
C269 a_11583_15239# VDPWR 0
C270 a_8377_5305# a_10553_4963# 0
C271 sky130_fd_sc_hd__dfxbp_1_9.Q_N a_18667_32188# 0.09273f
C272 a_9317_5049# a_12430_4527# 0
C273 a_8051_22875# sky130_fd_sc_hd__dfxbp_1_0.CLK 0
C274 sky130_fd_sc_hd__dfxbp_1_1.Q_N a_10550_22991# 0.05782f
C275 a_8038_5023# a_8377_5305# 0.04737f
C276 a_10995_12931# a_9771_12117# 0
C277 VDPWR a_9844_1793# 0.17124f
C278 a_6389_13769# VDPWR 0.47192f
C279 a_9705_12861# a_9703_16093# 0.4639f
C280 a_10160_4571# a_10471_5727# 0
C281 a_14491_5723# VDPWR 0.45275f
C282 a_18846_5265# a_18625_4938# 0.00783f
C283 a_12142_5459# a_12194_5433# 0.1439f
C284 sky130_fd_sc_hd__dfxbp_1_4.CLK sky130_fd_sc_hd__dfxbp_1_3.Q_N 0.15089f
C285 a_4847_14525# a_4505_13107# 0
C286 sky130_fd_sc_hd__dfxbp_1_2.CLK a_10807_23245# 0.00393f
C287 a_17689_23143# a_17647_22875# 0
C288 a_6911_15235# a_6635_15235# 0.00119f
C289 a_8377_5305# a_7315_5043# 0.21187f
C290 VDPWR a_7831_14003# 0
C291 a_10525_5837# a_10261_5837# 0
C292 a_12430_4527# a_12823_4919# 0.02301f
C293 a_17733_4529# a_17210_4895# 0
C294 a_9491_15377# a_8193_13753# 0
C295 a_18663_27017# a_18667_25510# 0
C296 a_18663_27756# VDPWR 0.19985f
C297 a_10986_1793# VDPWR 0
C298 a_5895_14763# a_6087_14735# 0
C299 a_1898_5051# a_2217_5025# 0.0073f
C300 a_10508_22879# a_10382_23245# 0.00553f
C301 a_17236_5473# a_16485_5729# 0.00682f
C302 VDPWR a_8729_23143# 0.51269f
C303 a_11501_15239# a_8193_13753# 0.1684f
C304 a_18667_31449# a_18671_29731# 0
C305 a_4840_5409# a_3229_5051# 0.03325f
C306 a_24234_14385# a_24152_14385# 0.04662f
C307 a_16583_4895# VDPWR 0
C308 a_9715_11297# a_10887_13773# 0
C309 a_10717_13773# a_9715_11297# 0.17512f
C310 a_6165_5043# a_6036_5017# 0.00758f
C311 a_9160_23197# a_8729_23143# 0.10805f
C312 a_14375_22875# a_12993_23237# 0
C313 sky130_fd_sc_hd__dfxbp_1_9.Q_N a_18667_34470# 0
C314 a_4849_11293# a_5933_13769# 0
C315 a_5851_13769# a_5933_13769# 0.00578f
C316 sky130_fd_sc_hd__dfxbp_1_2.CLK sky130_fd_sc_hd__dfxbp_1_3.CLK 0.00105f
C317 a_10499_4853# a_12378_4553# 0
C318 a_10382_23245# a_10297_22879# 0.03733f
C319 a_16129_2159# VDPWR 0
C320 a_9556_17271# VDPWR 1.27647f
C321 a_14596_1793# a_13167_1793# 0.08907f
C322 a_11671_15239# a_11501_15239# 0.00167f
C323 a_4329_2043# a_3199_1791# 0.21188f
C324 a_11439_4597# a_13709_4553# 0
C325 a_24152_14385# a_24318_14385# 0.05583f
C326 a_10953_14739# a_9715_11297# 0.00179f
C327 a_12430_4527# a_12533_5715# 0
C328 a_4839_12857# a_4595_14775# 0
C329 a_9317_5049# a_13473_5459# 0.04695f
C330 a_18667_24771# sky130_fd_sc_hd__dfxbp_1_7.CLK 0
C331 a_3199_1791# a_4746_2153# 0.03325f
C332 a_14380_4547# a_6238_6077# 0
C333 a_4905_12113# a_6089_11935# 0
C334 a_18667_33731# a_18667_33834# 0.14145f
C335 a_6261_5409# a_6375_5299# 0
C336 a_10385_4597# VDPWR 0.00132f
C337 a_6238_6077# a_14825_4913# 0
C338 a_12950_5459# a_14152_5441# 0
C339 a_4847_14525# a_5809_14763# 0.00524f
C340 a_13592_23193# sky130_fd_sc_hd__dfxbp_1_3.Q_N 0
C341 a_5363_5043# a_6261_5043# 0
C342 a_12129_22871# a_12993_23237# 0.03218f
C343 sky130_fd_sc_hd__dfxbp_1_9.Q_N a_19059_31529# 0.00188f
C344 a_8431_5049# a_8263_5049# 0
C345 a_12950_5459# a_12533_5715# 0.03016f
C346 sky130_fd_sc_hd__dfxbp_1_8.Q_N a_18667_32557# 0
C347 a_1920_1765# a_2145_2157# 0.00559f
C348 a_11255_13773# a_12039_15239# 0.00147f
C349 sky130_fd_sc_hd__dfxbp_1_5.Q_N a_18663_27545# 0
C350 a_5975_12927# a_6329_12927# 0.09582f
C351 a_6087_14735# a_5809_14763# 0.1109f
C352 sky130_fd_sc_hd__dfxbp_1_5.CLK a_18693_24621# 0
C353 VDPWR a_15838_23197# 0.21273f
C354 a_11255_13773# a_12615_14007# 0.00184f
C355 a_6238_6077# a_12430_4527# 0
C356 a_15242_5467# VDPWR 0
C357 sky130_fd_sc_hd__dfxbp_1_1.CLK a_8262_22875# 0
C358 a_17210_4529# a_6208_2817# 0
C359 a_12950_5825# a_12533_5715# 0.06611f
C360 a_9769_15349# a_10841_12931# 0
C361 a_7749_14003# a_4915_10549# 0.07615f
C362 a_10841_12931# VDPWR 0.23989f
C363 a_1920_1765# a_1868_1791# 0.1439f
C364 a_4847_14525# a_7173_15235# 0
C365 a_14561_4547# VDPWR 0.00119f
C366 a_18667_31449# sky130_fd_sc_hd__dfxbp_1_9.Q_N 0.11931f
C367 a_19063_29283# sky130_fd_sc_hd__dfxbp_1_9.CLK 0
C368 uo_out[0] uio_in[7] 0.03102f
C369 a_14152_5441# a_13473_5459# 0.11881f
C370 a_23133_17137# a_24962_14701# 0
C371 a_10916_4963# a_12430_4527# 0
C372 a_12950_5459# a_6238_6077# 0
C373 a_7113_13395# a_6281_11907# 0.19569f
C374 a_9503_10581# a_9631_11547# 0
C375 a_4839_12857# a_4903_15345# 0.1369f
C376 a_9769_15349# a_9703_16093# 0.50561f
C377 a_12533_5715# a_13473_5459# 0.1374f
C378 a_15711_4547# a_13709_4553# 0
C379 a_8231_23241# VDPWR 0.00345f
C380 a_6087_14735# a_7173_15235# 0.00327f
C381 a_4849_11293# a_6089_11935# 0
C382 a_10132_5445# a_10261_5837# 0.00792f
C383 a_9703_16093# VDPWR 1.32189f
C384 a_9781_10553# a_10869_11939# 0
C385 a_14375_22875# sky130_fd_sc_hd__dfxbp_1_3.Q_N 0.11931f
C386 a_12697_14007# VDPWR 0
C387 a_18667_24874# a_18667_24676# 0.1111f
C388 a_10525_5471# a_10471_5727# 0.00386f
C389 a_6238_6077# a_12950_5825# 0.00186f
C390 a_8038_5023# a_8263_5415# 0.00559f
C391 a_7221_1787# a_8700_2159# 0.03325f
C392 sky130_fd_sc_hd__dfxbp_1_4.CLK a_17647_22875# 0
C393 a_10717_13773# a_10993_13773# 0.00119f
C394 sky130_fd_sc_hd__dfxbp_1_2.CLK a_10550_22991# 0
C395 a_2079_5051# a_2343_5051# 0
C396 a_12769_4809# VDPWR 0.45983f
C397 uo_out[0] VDPWR 1.72112f
C398 a_12227_2049# a_13167_1793# 0.13739f
C399 VDPWR a_4597_11543# 0.02521f
C400 a_11255_13773# a_11979_13399# 0.06148f
C401 a_9317_5049# a_14491_5723# 0
C402 a_19059_25272# sky130_fd_sc_hd__dfxbp_1_7.CLK 0
C403 a_18663_27756# a_18671_29203# 0
C404 a_4903_15345# a_4635_13809# 0.00159f
C405 a_6238_6077# ui_in[1] 0
C406 a_11195_12931# a_9715_11297# 0.00976f
C407 a_6261_5409# a_6036_5017# 0.00559f
C408 a_8794_5415# a_7315_5043# 0.03325f
C409 a_10553_4963# VDPWR 0.05574f
C410 sky130_fd_sc_hd__dfxbp_1_6.Q_N a_18663_27545# 0
C411 a_17096_23241# a_17222_22875# 0.00553f
C412 a_9223_1793# a_11175_1793# 0
C413 a_16583_4895# a_16454_4503# 0.00792f
C414 a_18128_16189# a_18113_17153# 0.01375f
C415 a_5174_5409# a_5363_5043# 0
C416 a_10235_2049# a_11836_1793# 0
C417 a_8038_5023# VDPWR 0.34968f
C418 a_19059_24851# VDPWR 0
C419 a_18667_33636# sky130_fd_sc_hd__inv_2_0.A 0
C420 a_6238_6077# a_13473_5459# 0.00671f
C421 a_14179_2049# a_13167_1793# 0.21187f
C422 a_8431_5415# a_6238_6077# 0
C423 a_11439_4597# a_13186_4919# 0.03325f
C424 a_13186_4553# VDPWR 0.21831f
C425 a_9379_14779# a_4915_10549# 0
C426 VDPWR a_18667_33731# 0.66159f
C427 sky130_fd_sc_hd__dfxbp_1_7.Q sky130_fd_sc_hd__dfxbp_1_7.CLK 0.00137f
C428 a_7927_14003# VDPWR 0
C429 ui_in[0] a_24774_14701# 0.022f
C430 a_13077_23237# a_12736_22983# 0
C431 a_18667_33636# a_18667_33966# 0.07715f
C432 a_4837_16089# a_4903_15345# 0.50561f
C433 a_10297_22879# a_10477_23245# 0.00123f
C434 a_6129_12927# a_4913_13781# 0
C435 a_17733_4529# VDPWR 0.4178f
C436 a_15641_17149# a_15693_17123# 0.11638f
C437 uio_in[4] uio_in[5] 0.03102f
C438 a_7315_5043# VDPWR 1.39221f
C439 a_12129_22871# a_10109_22879# 0
C440 a_6021_13769# VDPWR 0
C441 a_6862_13645# a_6281_11907# 0.00254f
C442 a_12694_22871# a_12736_22983# 0
C443 a_16902_5473# a_16485_5729# 0.03016f
C444 a_6717_15235# VDPWR 0
C445 sky130_fd_sc_hd__dfxbp_1_0.CLK a_24962_14701# 0.14425f
C446 a_8073_1793# VDPWR 0.00115f
C447 a_18693_31299# VDPWR 0.07702f
C448 a_6281_2043# a_7032_2153# 0.00696f
C449 a_14152_5441# a_14491_5723# 0.04737f
C450 sky130_fd_sc_hd__dfxbp_1_9.Q_N a_18667_31684# 0.04247f
C451 sky130_fd_sc_hd__dfxbp_1_9.Q a_18667_33731# 0.25126f
C452 a_9705_12861# a_9493_12145# 0
C453 a_8193_13753# a_4915_10549# 0.14315f
C454 a_15641_17149# VDPWR 0.67139f
C455 sky130_fd_sc_hd__dfxbp_1_9.CLK a_18671_29108# 0
C456 a_6281_2043# a_7221_1787# 0.13739f
C457 a_18671_29438# a_18697_29053# 0.03733f
C458 sky130_fd_sc_hd__dfxbp_1_4.Q_N a_16657_22875# 0.11931f
C459 a_18667_25006# sky130_fd_sc_hd__dfxbp_1_7.CLK 0
C460 a_14179_2049# a_15904_1767# 0.00358f
C461 VDPWR a_7999_14003# 0
C462 a_10132_5445# a_10080_5471# 0.1439f
C463 sky130_fd_sc_hd__dfxbp_1_9.Q a_18693_31299# 0
C464 a_18689_26867# a_18663_27017# 0.06222f
C465 a_13077_23237# VDPWR 0.00627f
C466 a_18667_31977# a_18667_33731# 0
C467 a_9779_13785# a_4915_10549# 0.00435f
C468 a_18663_27756# a_18663_27120# 0.03684f
C469 a_5942_1761# a_6167_1787# 0.00487f
C470 a_3229_5051# a_3040_5417# 0
C471 a_16275_5839# a_16539_5839# 0
C472 a_9371_13111# a_9631_11547# 0
C473 a_18667_24771# a_18667_25879# 0
C474 a_7697_22875# a_10109_22879# 0
C475 sky130_fd_sc_hd__dfxbp_1_6.Q_N a_18697_29053# 0.142f
C476 a_10717_13773# a_10887_13773# 0.00167f
C477 a_16583_4895# a_16847_4895# 0
C478 a_6329_12927# VDPWR 0.31272f
C479 a_12694_22871# VDPWR 0
C480 a_8337_2159# a_8700_2159# 0.00847f
C481 a_21506_16181# a_23133_17137# 0
C482 a_6238_6077# a_14491_5723# 0.00768f
C483 sky130_fd_sc_hd__dfxbp_1_4.CLK a_14541_22875# 0
C484 a_10235_2049# a_10652_2159# 0.06611f
C485 a_6375_5299# a_5363_5043# 0.21187f
C486 sky130_fd_sc_hd__dfxbp_1_5.Q_N a_18663_27017# 0.00248f
C487 a_10717_13773# a_10953_14739# 0
C488 a_1950_5025# VDPWR 0.36044f
C489 a_9896_1767# a_8283_2049# 0.00419f
C490 a_2289_5307# a_2706_5051# 0.03016f
C491 a_17605_23241# a_16823_22875# 0
C492 a_9705_12861# a_10995_12931# 0.00312f
C493 a_4753_16089# VDPWR 0.00472f
C494 a_3199_1791# a_5269_1787# 0
C495 a_12587_5825# a_12194_5433# 0.02301f
C496 a_11175_1793# a_10986_2159# 0
C497 a_9461_14779# a_9379_14779# 0.00641f
C498 a_17733_4529# a_16679_4895# 0
C499 a_18663_27545# sky130_fd_sc_hd__dfxbp_1_7.Q_N 0.12218f
C500 VDPWR a_18663_26922# 0.31445f
C501 a_9621_12861# a_4915_10549# 0
C502 a_18667_31552# sky130_fd_sc_hd__dfxbp_1_9.CLK 0
C503 VDPWR a_7032_2153# 0
C504 a_4329_2043# VDPWR 0.45087f
C505 a_16243_2049# VDPWR 0.43625f
C506 a_6208_2817# a_13167_1793# 0.00283f
C507 a_4711_15373# a_4625_15373# 0.00658f
C508 a_17222_22875# VDPWR 0
C509 a_16297_2159# a_15904_1767# 0.02301f
C510 a_6281_2043# a_7892_1793# 0
C511 a_12430_4527# a_12559_4553# 0.00758f
C512 a_9381_11547# a_9771_12117# 0
C513 a_4839_12857# a_7749_14003# 0
C514 a_12663_23237# a_12568_23237# 0.00772f
C515 a_5975_12927# a_7113_13395# 0
C516 a_8431_5049# a_8794_5049# 0.00985f
C517 a_16583_4895# a_6238_6077# 0
C518 a_9223_1793# a_9896_1767# 0.11878f
C519 a_14771_4803# a_15522_4913# 0.00696f
C520 sky130_fd_sc_hd__inv_2_0.A a_18667_33834# 0
C521 a_4746_2153# VDPWR 0.02101f
C522 a_7221_1787# VDPWR 1.39111f
C523 a_9317_5049# a_12769_4809# 0
C524 a_3990_1761# a_4119_2153# 0.00792f
C525 a_4423_5299# a_4477_5043# 0.00386f
C526 a_6238_6077# a_9556_17271# 0.0058f
C527 a_4477_5043# VDPWR 0.18614f
C528 a_21506_16181# a_21491_17145# 0.01682f
C529 a_6429_5043# a_6165_5043# 0
C530 a_12587_5459# a_12194_5433# 0.02283f
C531 a_18667_33966# a_18667_33834# 0.23675f
C532 a_18693_33581# sky130_fd_sc_hd__dfxbp_1_8.Q_N 0.142f
C533 a_17733_4529# a_16454_4503# 0
C534 a_23133_17137# a_24774_14701# 0
C535 a_9896_1767# a_10289_1793# 0.02283f
C536 a_14380_4547# a_13473_5459# 0
C537 a_12017_1793# a_6208_2817# 0
C538 a_2187_1765# a_4383_2153# 0
C539 a_9715_11297# a_10841_12931# 0.18585f
C540 VDPWR a_5890_1787# 0.17124f
C541 sky130_fd_sc_hd__inv_12_0.A VDPWR 1.65409f
C542 sky130_fd_sc_hd__dfxbp_1_1.CLK sky130_fd_sc_hd__dfxbp_1_0.CLK 0
C543 a_12823_4919# a_12769_4809# 0.03622f
C544 a_9621_13111# a_4915_10549# 0
C545 a_15407_23143# sky130_fd_sc_hd__dfxbp_1_3.Q_N 0.12218f
C546 a_6281_2043# a_8337_2159# 0
C547 a_17521_23241# a_16657_22875# 0.03218f
C548 a_15904_1767# a_6208_2817# 0.00324f
C549 a_6629_15387# VDPWR 1.52787f
C550 a_14545_5467# VDPWR 0.18447f
C551 a_9317_5049# a_7315_5043# 0
C552 a_5984_5043# a_6036_5017# 0.1439f
C553 a_9317_5049# a_17733_4529# 0.37402f
C554 a_8136_23241# a_7697_22875# 0.27314f
C555 a_14375_22875# a_14909_23241# 0.0027f
C556 a_9493_12145# VDPWR 0.44497f
C557 a_12113_2159# a_12281_2159# 0
C558 a_5363_5043# a_6036_5017# 0.11878f
C559 a_9715_11297# a_9703_16093# 0.03118f
C560 a_15904_1767# a_16033_2159# 0.00792f
C561 a_8337_1793# a_8700_1793# 0.00985f
C562 a_15242_5467# a_6238_6077# 0
C563 sky130_fd_sc_hd__dfxbp_1_7.CLK a_18667_25299# 0.12322f
C564 a_17733_4529# a_16793_4785# 0.14301f
C565 a_10382_23245# sky130_fd_sc_hd__dfxbp_1_1.CLK 0
C566 sky130_fd_sc_hd__dfxbp_1_7.Q_N a_18697_29053# 0
C567 a_5975_12927# a_6862_13645# 0
C568 a_19510_16177# VDPWR 0.45244f
C569 a_18663_27017# a_18663_27252# 0.27314f
C570 a_12533_5715# a_12769_4809# 0
C571 a_4903_15345# a_5851_13769# 0.16757f
C572 a_4849_11293# a_4903_15345# 0.30637f
C573 VDPWR a_7892_1793# 0.16676f
C574 a_4839_12857# a_6057_12927# 0.00148f
C575 a_16471_17161# a_15693_17123# 0.09786f
C576 a_10717_13773# a_11195_12931# 0
C577 a_9371_13111# a_9713_14529# 0
C578 a_13788_1793# VDPWR 0.16897f
C579 a_6335_2153# a_6071_2153# 0
C580 a_4847_14525# a_6087_14735# 0.3079f
C581 a_4625_15373# a_4903_15345# 0.12165f
C582 a_14375_22875# a_14541_22875# 0.96835f
C583 a_10953_14739# a_11195_12931# 0
C584 sky130_fd_sc_hd__dfxbp_1_4.CLK a_14729_22875# 0
C585 a_7697_22875# a_8051_22875# 0.06222f
C586 a_10385_4963# a_10553_4963# 0
C587 a_12950_5459# a_13473_5459# 0
C588 a_9705_12861# a_9629_14779# 0.00187f
C589 sky130_fd_sc_hd__dfxbp_1_6.Q_N a_18667_32188# 0
C590 a_12194_5433# a_11439_4597# 0
C591 a_10235_2049# a_10986_1793# 0.00682f
C592 a_12655_4553# a_11439_4597# 0
C593 a_3990_1761# a_4215_2153# 0.00559f
C594 a_16471_17161# VDPWR 0.43619f
C595 a_6165_5409# a_5984_5043# 0
C596 a_19059_31950# sky130_fd_sc_hd__dfxbp_1_9.Q_N 0.00125f
C597 a_18120_23197# VDPWR 0.20884f
C598 a_2175_5051# a_2289_5307# 0
C599 a_9619_16343# VDPWR 0.33721f
C600 a_10995_12931# VDPWR 0
C601 a_17733_4529# a_16847_4895# 0
C602 a_18663_27756# a_18671_29108# 0
C603 a_6238_6077# a_12769_4809# 0
C604 a_24774_14701# sky130_fd_sc_hd__dfxbp_1_0.CLK 0.01196f
C605 a_2187_1765# a_4119_1787# 0
C606 a_18671_29203# a_18663_26922# 0
C607 VDPWR a_8337_2159# 0.0097f
C608 sky130_fd_sc_hd__inv_2_0.A VDPWR 0.34513f
C609 a_10289_4963# a_10553_4963# 0
C610 uo_out[0] sky130_fd_sc_hd__inv_16_0.A 1.50114f
C611 a_6375_5299# a_6792_5409# 0.06611f
C612 a_4329_2043# a_5080_1787# 0.00682f
C613 a_18667_32557# a_18667_33731# 0
C614 a_6238_6077# a_10553_4963# 0
C615 a_12129_22871# a_14541_22875# 0
C616 a_2313_1791# a_2145_1791# 0
C617 a_11255_13773# a_11147_11911# 0.00254f
C618 a_8038_5023# a_6238_6077# 0.00209f
C619 sky130_fd_sc_hd__dfxbp_1_4.CLK a_15239_23241# 0.00387f
C620 a_6281_2043# a_5269_1787# 0.21187f
C621 a_24234_14385# VDPWR 0.28779f
C622 a_14940_22875# sky130_fd_sc_hd__dfxbp_1_3.Q_N 0.00188f
C623 a_10652_1793# a_6208_2817# 0
C624 a_12129_22871# a_12663_23237# 0.0027f
C625 VDPWR a_18667_33966# 0.25541f
C626 a_10953_14739# a_11583_15239# 0.00232f
C627 a_18667_24874# a_18667_25510# 0.03684f
C628 a_11888_1767# a_12281_2159# 0.02301f
C629 a_2079_5051# VDPWR 0.00123f
C630 a_16902_5839# a_16539_5839# 0.00847f
C631 a_2343_5417# a_2175_5417# 0
C632 sky130_fd_sc_hd__inv_2_0.A sky130_fd_sc_hd__dfxbp_1_9.Q 0.00149f
C633 a_10525_5837# a_12194_5433# 0
C634 a_18671_29306# a_18671_29731# 0
C635 VDPWR a_24318_14385# 0.00521f
C636 a_6127_13769# a_6389_13769# 0
C637 a_18663_27017# sky130_fd_sc_hd__dfxbp_1_7.Q_N 0.11931f
C638 a_10916_4963# a_10553_4963# 0.00847f
C639 a_6238_6077# a_7315_5043# 0.00286f
C640 a_7113_13395# VDPWR 0.49786f
C641 a_17733_4529# a_6238_6077# 0.01989f
C642 a_2187_1765# a_4746_1787# 0
C643 a_8136_23241# a_8304_22987# 0.23992f
C644 a_16994_1793# VDPWR 0
C645 a_17544_4529# a_6208_2817# 0
C646 a_17096_23241# a_17264_22987# 0.23992f
C647 a_9703_16093# a_10993_13773# 0.00702f
C648 sky130_fd_sc_hd__dfxbp_1_9.Q a_18667_33966# 0
C649 a_13077_23237# sky130_fd_sc_hd__dfxbp_1_2.Q_N 0
C650 a_6208_2817# a_16129_1793# 0
C651 a_6635_15235# a_4903_15345# 0
C652 a_20384_16179# a_9556_17271# 0
C653 VDPWR a_10471_5727# 0.46233f
C654 a_23761_14335# a_24962_14701# 0.09435f
C655 a_3229_5051# a_4213_5043# 0
C656 a_24234_14385# a_23731_14309# 0.12294f
C657 a_13119_22871# a_12736_22983# 0
C658 a_12694_22871# sky130_fd_sc_hd__dfxbp_1_2.Q_N 0.00188f
C659 a_6208_2817# ui_in[0] 0.0357f
C660 VDPWR a_18667_24771# 0.65217f
C661 a_18667_34839# VDPWR 0.21263f
C662 a_9781_10553# a_4915_10549# 0.00418f
C663 a_16485_5729# a_16539_5839# 0.03622f
C664 a_18667_31449# a_18671_29438# 0
C665 a_8167_5049# VDPWR 0.00115f
C666 a_8051_22875# a_8304_22987# 0
C667 sky130_fd_sc_hd__dfxbp_1_5.CLK a_17222_22875# 0
C668 a_9943_22879# a_8729_23143# 0
C669 a_9631_11297# VDPWR 0.00377f
C670 a_23731_14309# a_24318_14385# 0.02707f
C671 uo_out[5] uo_out[4] 0.03102f
C672 a_18663_27120# a_18663_26922# 0.1111f
C673 a_16902_5839# a_15431_5467# 0.03325f
C674 a_5975_12927# a_4913_13781# 0.08477f
C675 sky130_fd_sc_hd__dfxbp_1_7.Q a_18663_28125# 0.2081f
C676 a_5269_1787# VDPWR 1.3928f
C677 a_13709_4553# a_14908_5833# 0
C678 a_14375_22875# a_14729_22875# 0.06222f
C679 a_12295_22871# a_13161_23139# 0.03136f
C680 a_19055_27518# sky130_fd_sc_hd__dfxbp_1_7.CLK 0
C681 a_18667_31449# sky130_fd_sc_hd__dfxbp_1_6.Q_N 0.00248f
C682 a_2079_5417# a_2217_5025# 0
C683 a_8561_23241# sky130_fd_sc_hd__dfxbp_1_1.CLK 0.0039f
C684 a_16275_5839# VDPWR 0
C685 a_17425_5473# a_17733_4529# 0.39935f
C686 a_4032_5043# a_2217_5025# 0.00121f
C687 a_11411_5471# a_13186_4919# 0
C688 a_18846_5265# VDPWR 0
C689 a_3199_1791# a_3938_1787# 0.04946f
C690 a_13473_5459# a_14491_5723# 0.21187f
C691 a_24241_14651# VDPWR 0.27707f
C692 a_3990_1761# a_4383_1787# 0.02283f
C693 a_3229_5051# a_4477_5409# 0.04534f
C694 a_9629_14779# a_9769_15349# 0.00327f
C695 a_15188_4547# a_14491_5723# 0
C696 a_6862_13645# VDPWR 0.16013f
C697 a_9629_14779# VDPWR 0.33336f
C698 a_4913_13781# a_4513_14775# 0
C699 a_12993_23237# a_12736_22983# 0.03684f
C700 a_5942_1761# a_6335_2153# 0.02301f
C701 a_13119_22871# VDPWR 0
C702 a_15711_4547# a_14771_4803# 0.13762f
C703 a_7749_14003# a_5851_13769# 0
C704 a_12281_1793# a_12644_1793# 0.00985f
C705 a_4637_10577# a_4723_10577# 0.00658f
C706 a_10717_13773# a_10841_12931# 0
C707 a_12644_1793# VDPWR 0.21795f
C708 a_10888_5471# a_10471_5727# 0.03016f
C709 a_11888_1767# a_11175_1793# 0.11874f
C710 a_9781_10553# a_12865_14007# 0
C711 a_18689_26867# a_18689_27047# 0.00123f
C712 a_17096_23241# sky130_fd_sc_hd__dfxbp_1_3.Q_N 0
C713 uio_oe[5] uio_oe[4] 0.03102f
C714 sky130_fd_sc_hd__dfxbp_1_1.Q_N sky130_fd_sc_hd__dfxbp_1_0.Q_N 0
C715 a_18667_25879# a_18667_25299# 0.10805f
C716 a_10382_23245# a_10550_22991# 0.23992f
C717 a_14375_22875# a_15239_23241# 0.03218f
C718 a_16485_5729# a_15431_5467# 0.21187f
C719 a_14545_5467# a_14152_5441# 0.02283f
C720 a_5269_1787# a_6698_2153# 0.03325f
C721 a_14982_22987# sky130_fd_sc_hd__dfxbp_1_4.CLK 0
C722 a_3229_5051# a_2217_5025# 0.00481f
C723 a_15119_1793# a_13167_1793# 0
C724 a_1898_5051# VDPWR 0.17586f
C725 a_6003_11935# a_4913_13781# 0
C726 a_17236_5839# a_16485_5729# 0.00696f
C727 a_19055_27097# a_18663_27252# 0.00553f
C728 a_10717_13773# a_9703_16093# 0.08387f
C729 a_9703_16093# a_10887_13773# 0.00246f
C730 a_10761_14767# a_10675_14767# 0.00658f
C731 a_14380_4547# a_12769_4809# 0
C732 sky130_fd_sc_hd__dfxbp_1_7.Q a_18671_29942# 0
C733 a_9715_11297# a_9493_12145# 0.0022f
C734 a_23731_14309# a_24241_14651# 0.02645f
C735 a_9381_11547# a_9705_12861# 0
C736 a_19510_16177# a_19235_17155# 0.00704f
C737 a_19059_25272# VDPWR 0
C738 a_8193_13753# sky130_fd_sc_hd__dfxbp_1_0.CLK 0
C739 a_6281_11907# a_6089_11935# 0
C740 a_7173_15235# a_4915_10549# 0.09278f
C741 VDPWR a_18667_31354# 0.31446f
C742 a_10953_14739# a_9703_16093# 0.29394f
C743 a_12993_23237# VDPWR 0.19825f
C744 a_6208_2817# a_11439_4597# 0.00105f
C745 a_15407_23143# a_14541_22875# 0.03136f
C746 a_17264_22987# VDPWR 0.19112f
C747 a_9781_10553# a_9589_10581# 0
C748 a_17210_4895# a_16485_5729# 0
C749 a_16243_2049# a_16994_2159# 0.00696f
C750 a_8687_22875# a_8561_23241# 0.00617f
C751 sky130_fd_sc_hd__dfxbp_1_7.Q a_19063_29704# 0
C752 a_10916_4597# VDPWR 0.31232f
C753 a_4847_14525# a_4763_14525# 0.00206f
C754 sky130_fd_sc_hd__inv_12_0.A sky130_fd_sc_hd__inv_16_0.A 1.38086f
C755 sky130_fd_sc_hd__dfxbp_1_4.CLK sky130_fd_sc_hd__dfxbp_1_3.CLK 0.00137f
C756 a_10888_5837# a_10525_5837# 0.00847f
C757 a_18667_34259# a_19059_34232# 0
C758 a_12430_4527# a_12769_4809# 0.04737f
C759 a_12039_15239# a_10675_14767# 0
C760 a_6238_6077# a_14545_5467# 0
C761 a_2313_1791# a_2676_1791# 0.00985f
C762 a_8283_2049# a_7944_1767# 0.04737f
C763 a_8136_23241# a_7863_22875# 0.07715f
C764 sky130_fd_sc_hd__dfxbp_1_7.Q VDPWR 0.27299f
C765 sky130_fd_sc_hd__dfxbp_1_5.CLK a_18120_23197# 0.20225f
C766 sky130_fd_sc_hd__dfxbp_1_9.Q a_18667_31354# 0
C767 a_15904_1767# a_15119_1793# 0.11873f
C768 sky130_fd_sc_hd__dfxbp_1_6.Q_N a_18667_31684# 0
C769 a_4839_12857# a_4755_12857# 0.00208f
C770 a_4849_11293# a_6057_12927# 0.00146f
C771 a_11979_13399# a_11728_13649# 0.10945f
C772 a_2259_2047# a_3010_2157# 0.00696f
C773 a_6208_2817# a_23133_17137# 0
C774 sky130_fd_sc_hd__dfxbp_1_3.CLK a_12568_23237# 0
C775 a_9503_10581# a_4915_10549# 0.00102f
C776 a_9715_11297# a_10995_12931# 0
C777 a_6389_13769# a_7831_14003# 0
C778 a_18667_24676# sky130_fd_sc_hd__dfxbp_1_7.CLK 0
C779 a_9317_5049# a_10471_5727# 0
C780 a_6429_5043# a_5363_5043# 0.08312f
C781 a_5269_1787# a_6071_1787# 0
C782 a_18697_29647# a_18671_29942# 0.00851f
C783 a_18667_31977# a_18667_31354# 0.03136f
C784 a_4753_16339# VDPWR 0.33641f
C785 a_10975_23147# a_10109_22879# 0.03136f
C786 a_12039_15239# a_8193_13753# 0.00221f
C787 a_2313_1791# a_2187_1765# 0.08436f
C788 sky130_fd_sc_hd__dfxbp_1_7.Q_N a_19055_27097# 0.00188f
C789 a_8051_22875# a_7863_22875# 0.0967f
C790 a_18671_29731# a_18671_30311# 0.10805f
C791 a_6208_2817# a_10108_4597# 0
C792 sky130_fd_sc_hd__dfxbp_1_8.Q_N a_18667_33731# 0.11931f
C793 a_18667_25006# VDPWR 0.25526f
C794 a_10025_2159# VDPWR 0
C795 VDPWR a_10891_23245# 0.00629f
C796 a_18693_33581# a_18667_33731# 0.06222f
C797 sky130_fd_sc_hd__dfxbp_1_1.Q_N a_12295_22871# 0.00115f
C798 a_18667_31552# a_18693_31299# 0
C799 a_18693_31299# sky130_fd_sc_hd__dfxbp_1_9.CLK 0
C800 uio_out[7] uio_oe[0] 0.03102f
C801 a_12227_2049# a_12978_2159# 0.00696f
C802 uio_oe[7] uio_oe[6] 0.03102f
C803 a_10499_4853# a_6208_2817# 0
C804 a_15711_4547# a_6208_2817# 0.00103f
C805 a_11195_12931# a_10841_12931# 0.09582f
C806 a_5895_14763# a_4839_12857# 0
C807 VDPWR a_4913_13781# 0.75079f
C808 a_11671_15239# a_12039_15239# 0
C809 a_4839_12857# a_4505_13107# 0.16952f
C810 a_13592_23193# sky130_fd_sc_hd__dfxbp_1_3.CLK 0.20774f
C811 a_2676_2157# VDPWR 0.02202f
C812 a_18697_29647# VDPWR 0.00627f
C813 VDPWR sky130_fd_sc_hd__dfxbp_1_3.Q_N 0.60679f
C814 a_13473_5459# a_12769_4809# 0
C815 a_7221_1787# a_8700_1793# 0.08907f
C816 a_15188_4547# a_12769_4809# 0
C817 a_6335_1787# a_6167_1787# 0
C818 a_20109_17157# a_18113_17153# 0
C819 sky130_fd_sc_hd__dfxbp_1_5.Q_N a_18667_24874# 0.05782f
C820 a_18689_27047# a_18663_27252# 0.00772f
C821 uio_oe[2] uio_oe[1] 0.03102f
C822 a_23761_14335# a_24774_14701# 0.33858f
C823 a_4505_13107# a_4515_11543# 0.00102f
C824 a_14982_22987# a_14375_22875# 0.14145f
C825 a_16539_5473# a_16485_5729# 0.00386f
C826 a_6911_15235# VDPWR 0
C827 sky130_fd_sc_hd__dfxbp_1_5.CLK a_18667_24771# 0.24944f
C828 a_24234_14385# a_6238_6077# 0.07599f
C829 a_4505_13107# a_4635_13809# 0.00115f
C830 a_10109_22879# VDPWR 0.31445f
C831 a_9579_12145# a_4915_10549# 0
C832 a_8038_5023# a_8431_5415# 0.02301f
C833 a_6208_2817# a_16297_1793# 0
C834 a_4839_12857# a_6944_13645# 0
C835 a_16902_5839# VDPWR 0.01944f
C836 a_9381_11547# VDPWR 0.53681f
C837 a_6238_6077# a_24318_14385# 0.04268f
C838 a_6208_2817# sky130_fd_sc_hd__dfxbp_1_0.CLK 0
C839 a_15242_5467# a_14491_5723# 0.00682f
C840 a_18671_29203# a_18667_31354# 0
C841 uo_out[6] uo_out[5] 0.03102f
C842 a_9631_11297# a_9715_11297# 0.00206f
C843 a_11250_4597# VDPWR 0
C844 a_11501_15239# a_11777_15239# 0.00119f
C845 a_5895_14763# a_4837_16089# 0
C846 a_12559_4919# VDPWR 0
C847 a_9503_10581# a_9589_10581# 0.00658f
C848 a_14375_22875# sky130_fd_sc_hd__dfxbp_1_3.CLK 0.25091f
C849 a_8431_5415# a_7315_5043# 0.04534f
C850 a_9713_14529# a_9491_15377# 0.00215f
C851 a_12129_22871# a_10807_23245# 0
C852 a_18671_30311# sky130_fd_sc_hd__dfxbp_1_9.Q_N 0
C853 a_9705_12861# a_11255_13773# 0.04676f
C854 a_7697_22875# sky130_fd_sc_hd__dfxbp_1_1.CLK 0
C855 a_4839_12857# a_5809_14763# 0.21988f
C856 a_11411_5471# a_12194_5433# 0.11876f
C857 a_11583_15239# a_9703_16093# 0
C858 a_12281_2159# VDPWR 0.0097f
C859 a_6238_6077# a_10471_5727# 0.00739f
C860 a_9713_14529# a_11501_15239# 0.17824f
C861 a_7944_1767# a_8169_1793# 0.00487f
C862 a_15119_1793# a_16129_1793# 0
C863 sky130_fd_sc_hd__dfxbp_1_7.Q a_18671_29203# 0.25135f
C864 a_19059_34232# a_18667_34470# 0.00617f
C865 a_6208_2817# a_6335_2153# 0
C866 a_4084_5017# a_4309_5043# 0.00487f
C867 a_14233_1793# a_13167_1793# 0.08312f
C868 a_2217_5025# a_5984_5043# 0.00121f
C869 a_6208_2817# a_12017_2159# 0
C870 a_9715_11297# a_9629_14779# 0
C871 a_9371_13111# a_4915_10549# 0.00232f
C872 a_7986_5049# a_8167_5415# 0
C873 a_7749_14003# a_9501_13813# 0
C874 a_15407_23143# a_15239_23241# 0.31062f
C875 a_8167_5049# a_6238_6077# 0
C876 a_5363_5043# a_2217_5025# 0.00133f
C877 a_16371_5473# a_16146_5447# 0.00487f
C878 a_3938_1787# VDPWR 0.16677f
C879 a_13119_22871# sky130_fd_sc_hd__dfxbp_1_2.Q_N 0.00125f
C880 a_16485_5729# VDPWR 0.43937f
C881 a_12129_22871# sky130_fd_sc_hd__dfxbp_1_3.CLK 0
C882 a_4839_12857# a_7173_15235# 0.00585f
C883 a_1950_5025# a_2289_5307# 0.04737f
C884 a_16660_1793# VDPWR 0.21452f
C885 a_14825_4547# a_14432_4521# 0.02283f
C886 a_6238_6077# a_16275_5839# 0
C887 a_10499_4853# a_10553_4597# 0.00386f
C888 a_18846_5265# a_6238_6077# 0.00101f
C889 a_6238_6077# a_24241_14651# 0.03341f
C890 a_1950_5025# a_2175_5051# 0.00487f
C891 VDPWR a_18667_25299# 0.51563f
C892 sky130_fd_sc_hd__dfxbp_1_5.CLK a_17264_22987# 0
C893 a_5809_14763# a_4837_16089# 0.03093f
C894 a_18693_31893# VDPWR 0.00628f
C895 a_8136_23241# VDPWR 0.25517f
C896 a_20384_16179# a_19510_16177# 0.101f
C897 a_9369_16343# a_9769_15349# 0
C898 a_9631_11547# a_4915_10549# 0
C899 a_18663_27545# a_18697_29053# 0
C900 a_9556_17271# a_9703_16093# 0
C901 a_6208_2817# a_12978_2159# 0
C902 a_9781_10553# a_10955_11939# 0
C903 a_9369_16343# VDPWR 0.54727f
C904 a_6003_11935# a_6089_11935# 0.00658f
C905 a_14825_4547# a_13709_4553# 0.08312f
C906 a_6389_13769# a_6021_13769# 0
C907 a_8337_1793# a_8073_1793# 0
C908 a_6375_5299# a_6792_5043# 0.03016f
C909 a_12993_23237# sky130_fd_sc_hd__dfxbp_1_2.Q_N 0.09273f
C910 a_17647_22875# VDPWR 0
C911 sky130_fd_sc_hd__dfxbp_1_2.CLK a_12295_22871# 0.014f
C912 a_4477_5043# a_2289_5307# 0
C913 a_15431_5467# a_13709_4553# 0
C914 a_12194_5433# a_12419_5459# 0.00487f
C915 VDPWR a_5933_13769# 0
C916 sky130_fd_sc_hd__dfxbp_1_1.Q_N a_13161_23139# 0
C917 a_19059_33811# a_18667_33834# 0
C918 a_14814_23241# sky130_fd_sc_hd__dfxbp_1_3.Q_N 0.04247f
C919 a_7173_15235# a_4837_16089# 0.04212f
C920 a_9379_14779# a_9501_13813# 0.00144f
C921 sky130_fd_sc_hd__dfxbp_1_7.Q a_18663_27120# 0
C922 a_8051_22875# VDPWR 0.07692f
C923 sky130_fd_sc_hd__dfxbp_1_1.CLK a_8304_22987# 0
C924 a_12281_1793# a_11175_1793# 0.08312f
C925 a_10508_22879# VDPWR 0
C926 a_2259_2047# a_3990_1761# 0.00332f
C927 sky130_fd_sc_hd__dfxbp_1_0.Q_N a_8262_22875# 0.00188f
C928 a_4905_12113# a_4505_13107# 0
C929 a_11175_1793# VDPWR 1.39052f
C930 a_6208_2817# a_8283_2049# 0.00304f
C931 a_17425_5473# a_18846_5265# 0
C932 a_18667_25006# sky130_fd_sc_hd__dfxbp_1_5.CLK 0
C933 a_9705_12861# a_9453_13111# 0
C934 a_6208_2817# a_10289_4597# 0
C935 a_9703_16093# a_10841_12931# 0
C936 a_4849_11293# a_4755_12857# 0
C937 a_24152_14385# a_24774_14701# 0
C938 VDPWR a_10297_22879# 0.07696f
C939 a_13840_1767# VDPWR 0.34959f
C940 a_4847_14525# a_4503_16339# 0
C941 a_8193_13753# a_9501_13813# 0.00125f
C942 a_6389_13769# a_6329_12927# 0.20048f
C943 a_11255_13773# a_9769_15349# 0
C944 a_11255_13773# VDPWR 0.47196f
C945 a_8377_5305# a_10080_5471# 0
C946 a_14561_4913# VDPWR 0
C947 a_4637_10577# a_4915_10549# 0.1296f
C948 a_14545_5467# a_13473_5459# 0.08314f
C949 a_9223_1793# a_6208_2817# 0.00284f
C950 a_9705_12861# a_9629_14529# 0
C951 sky130_fd_sc_hd__inv_2_0.A sky130_fd_sc_hd__dfxbp_1_8.Q_N 0.14589f
C952 a_9556_17271# a_15641_17149# 0.03788f
C953 a_18663_27017# a_18663_27545# 0.04808f
C954 a_12644_2159# VDPWR 0.02101f
C955 a_14982_22987# a_15407_23143# 0
C956 a_18693_33581# sky130_fd_sc_hd__inv_2_0.A 0
C957 VDPWR a_14909_23241# 0.00347f
C958 sky130_fd_sc_hd__dfxbp_1_7.Q a_19063_29283# 0
C959 a_9779_13785# a_9501_13813# 0.1205f
C960 a_6281_2043# a_6698_1787# 0.03016f
C961 a_16454_4503# a_16485_5729# 0
C962 uio_oe[2] uio_oe[3] 0.03102f
C963 a_11147_11911# a_11728_13649# 0.00254f
C964 a_4905_12113# a_4713_12141# 0
C965 a_16146_5447# a_16371_5839# 0.00559f
C966 sky130_fd_sc_hd__dfxbp_1_8.Q_N a_18667_33966# 0.04247f
C967 a_4477_5043# a_4840_5043# 0.00985f
C968 sky130_fd_sc_hd__dfxbp_1_2.Q_N sky130_fd_sc_hd__dfxbp_1_3.Q_N 0
C969 a_18693_33581# a_18667_33966# 0.03733f
C970 a_7221_1787# a_8337_1793# 0.08313f
C971 a_6208_2817# a_10289_1793# 0
C972 a_3199_1791# a_2676_1791# 0
C973 VDPWR a_6089_11935# 0
C974 a_5895_14763# a_4849_11293# 0.00121f
C975 a_14908_5467# a_15431_5467# 0
C976 a_4849_11293# a_4505_13107# 0.00372f
C977 a_12823_4919# a_12559_4919# 0
C978 a_18671_29306# a_18671_29438# 0.23675f
C979 sky130_fd_sc_hd__inv_4_0.A sky130_fd_sc_hd__inv_8_0.A 0
C980 a_8687_22875# a_8304_22987# 0
C981 a_9317_5049# a_16485_5729# 0
C982 a_17345_17163# a_17254_16187# 0.01682f
C983 a_9781_10553# a_12039_15239# 0.09278f
C984 a_18663_27756# a_18663_26922# 0.19462f
C985 a_12663_23237# a_12483_22871# 0.00123f
C986 a_4585_16339# VDPWR 0.0252f
C987 a_9713_14529# a_4915_10549# 0
C988 a_15407_23143# sky130_fd_sc_hd__dfxbp_1_3.CLK 0
C989 a_18667_25510# sky130_fd_sc_hd__dfxbp_1_7.CLK 0.0039f
C990 a_14541_22875# VDPWR 0.31445f
C991 a_9781_10553# a_12615_14007# 0.07615f
C992 sky130_fd_sc_hd__inv_8_0.A sky130_fd_sc_hd__inv_6_0.A 0.59805f
C993 a_10160_4571# a_8794_5049# 0
C994 a_9381_11547# a_9715_11297# 0.16782f
C995 a_16793_4785# a_16485_5729# 0
C996 a_18671_29306# sky130_fd_sc_hd__dfxbp_1_6.Q_N 0.05782f
C997 a_12663_23237# VDPWR 0.00345f
C998 VDPWR a_10261_5837# 0
C999 a_19059_33811# VDPWR 0
C1000 a_19055_27518# VDPWR 0
C1001 a_12378_4553# VDPWR 0.18081f
C1002 a_3199_1791# a_2187_1765# 0.00474f
C1003 a_6429_5409# a_6261_5409# 0
C1004 a_4595_14775# a_4513_14775# 0.00641f
C1005 a_24234_14385# ui_in[1] 0.12911f
C1006 a_4849_11293# a_6944_13645# 0
C1007 a_13969_1793# VDPWR 0.00116f
C1008 a_13186_4553# a_12769_4809# 0.03016f
C1009 a_15522_4547# a_14771_4803# 0.00682f
C1010 a_6629_15387# a_6389_13769# 0
C1011 a_16129_2159# a_16243_2049# 0
C1012 a_11810_13649# a_11255_13773# 0.00183f
C1013 a_15323_23241# sky130_fd_sc_hd__dfxbp_1_3.Q_N 0
C1014 sky130_fd_sc_hd__dfxbp_1_8.Q_N a_18667_34839# 0.12801f
C1015 a_4849_11293# a_4713_12141# 0
C1016 a_12950_5459# a_10471_5727# 0
C1017 a_2145_1791# VDPWR 0.00107f
C1018 a_14545_5467# a_14491_5723# 0.00386f
C1019 a_14545_5833# a_13709_4553# 0
C1020 ui_in[1] a_24318_14385# 0.00197f
C1021 a_19059_33811# sky130_fd_sc_hd__dfxbp_1_9.Q 0
C1022 a_18663_27017# a_18697_29053# 0
C1023 VDPWR a_6698_1787# 0.21797f
C1024 a_4723_10577# a_4915_10549# 0
C1025 a_16679_4529# a_6208_2817# 0
C1026 a_6238_6077# a_16902_5839# 0.00192f
C1027 sky130_fd_sc_hd__dfxbp_1_4.Q_N a_16823_22875# 0.5114f
C1028 a_16847_4529# a_14771_4803# 0
C1029 a_15119_1793# a_16297_1793# 0.08312f
C1030 a_6165_5043# VDPWR 0.00119f
C1031 a_4849_11293# a_5809_14763# 0.10553f
C1032 a_5809_14763# a_5851_13769# 0
C1033 a_10553_4597# a_10289_4597# 0
C1034 a_8038_5023# a_7315_5043# 0.11881f
C1035 a_9896_1767# VDPWR 0.34957f
C1036 sky130_fd_sc_hd__dfxbp_1_2.CLK a_13161_23139# 0
C1037 a_9621_13111# a_9501_13813# 0
C1038 a_9781_10553# a_11979_13399# 0.2011f
C1039 a_6208_2817# a_8169_1793# 0
C1040 a_14940_22875# a_14982_22987# 0
C1041 a_6208_2817# a_23761_14335# 0.06557f
C1042 a_6238_6077# a_12559_4919# 0
C1043 a_6208_2817# a_10986_2159# 0
C1044 a_7749_14003# a_6281_11907# 0.19234f
C1045 sky130_fd_sc_hd__inv_4_0.A a_18667_34259# 0
C1046 a_14596_2159# VDPWR 0.02101f
C1047 sky130_fd_sc_hd__inv_4_0.A sky130_fd_sc_hd__inv_6_0.A 0.40684f
C1048 a_17689_23143# sky130_fd_sc_hd__dfxbp_1_4.Q_N 0.12218f
C1049 a_5975_12927# a_4903_15345# 0
C1050 sky130_fd_sc_hd__dfxbp_1_5.CLK a_18667_25299# 0
C1051 sky130_fd_sc_hd__dfxbp_1_1.CLK a_7863_22875# 0
C1052 a_14432_4521# VDPWR 0.35495f
C1053 a_9453_13111# VDPWR 0.02522f
C1054 a_15365_22875# sky130_fd_sc_hd__dfxbp_1_3.Q_N 0.00125f
C1055 a_18693_24621# a_18667_24771# 0.06222f
C1056 a_16094_5473# a_16146_5447# 0.1439f
C1057 sky130_fd_sc_hd__dfxbp_1_7.Q a_18671_29108# 0.014f
C1058 a_15188_4913# VDPWR 0.02568f
C1059 a_6629_15387# a_9556_17271# 0.10733f
C1060 a_4849_11293# a_7173_15235# 0
C1061 a_2313_2157# a_2049_2157# 0
C1062 a_12587_5459# a_12323_5459# 0
C1063 a_7173_15235# a_5851_13769# 0
C1064 a_4903_15345# a_4513_14775# 0.00566f
C1065 sky130_fd_sc_hd__dfxbp_1_5.CLK a_17647_22875# 0
C1066 a_18667_33636# sky130_fd_sc_hd__dfxbp_1_9.Q_N 0.00105f
C1067 a_9629_14529# a_9769_15349# 0
C1068 a_4847_14525# a_4839_12857# 0.2003f
C1069 a_9629_14529# VDPWR 0.00474f
C1070 a_8377_5305# a_8263_5049# 0
C1071 a_9461_14779# a_9713_14529# 0
C1072 a_16660_2159# VDPWR 0.0192f
C1073 a_2313_1791# a_2049_1791# 0
C1074 a_14940_22875# sky130_fd_sc_hd__dfxbp_1_3.CLK 0
C1075 a_12323_5825# VDPWR 0
C1076 a_2217_5025# a_3040_5051# 0
C1077 a_6238_6077# a_16485_5729# 0.00779f
C1078 a_13709_4553# VDPWR 1.40616f
C1079 a_15711_4547# a_16146_5447# 0
C1080 a_8283_2049# a_9034_1793# 0.00682f
C1081 a_9779_13785# a_9771_12117# 0.00627f
C1082 a_18667_31552# a_18667_31354# 0.1111f
C1083 a_3199_1791# a_4215_1787# 0
C1084 sky130_fd_sc_hd__dfxbp_1_9.CLK a_18667_31354# 0.01405f
C1085 a_12227_2049# a_12113_2159# 0
C1086 a_9556_17271# a_19510_16177# 0
C1087 a_4839_12857# a_6087_14735# 0.02465f
C1088 a_12419_5825# VDPWR 0
C1089 ui_in[1] a_24241_14651# 0.00151f
C1090 a_14814_23241# a_14909_23241# 0.00772f
C1091 a_9463_11547# a_4915_10549# 0
C1092 a_2343_5417# a_4084_5017# 0
C1093 VDPWR a_10080_5471# 0.17025f
C1094 a_4847_14525# a_4635_13809# 0
C1095 a_13840_1767# a_14065_1793# 0.00487f
C1096 a_16275_5473# a_16146_5447# 0.00758f
C1097 a_21506_16181# a_22274_16171# 0.1036f
C1098 a_2217_5025# a_5174_5043# 0
C1099 a_13969_2159# VDPWR 0
C1100 a_2079_5417# VDPWR 0
C1101 VDPWR a_24962_14701# 0.29265f
C1102 a_18671_29306# sky130_fd_sc_hd__dfxbp_1_7.Q_N 0
C1103 a_4032_5043# VDPWR 0.1668f
C1104 a_14729_22875# VDPWR 0.07696f
C1105 a_4711_15373# VDPWR 0.00333f
C1106 a_18667_24676# VDPWR 0.31434f
C1107 a_13520_4553# a_6208_2817# 0
C1108 a_4119_2153# a_4383_2153# 0
C1109 sky130_fd_sc_hd__dfxbp_1_7.Q sky130_fd_sc_hd__dfxbp_1_9.CLK 0.00105f
C1110 ui_in[0] a_23511_14335# 0.01792f
C1111 a_18697_29647# a_18671_29108# 0
C1112 a_7113_13395# a_6389_13769# 0.06148f
C1113 a_9223_1793# a_10025_1793# 0
C1114 a_6375_5299# a_7126_5043# 0.00682f
C1115 a_9556_17271# a_9619_16343# 0
C1116 sky130_fd_sc_hd__dfxbp_1_4.Q_N a_17011_22875# 0.142f
C1117 a_4637_10577# a_4515_11543# 0.00144f
C1118 a_14541_22875# a_14814_23241# 0.07715f
C1119 a_12978_1793# VDPWR 0
C1120 a_4847_14525# a_4837_16089# 0.46421f
C1121 a_6208_2817# a_10160_4571# 0
C1122 sky130_fd_sc_hd__dfxbp_1_0.Q_N sky130_fd_sc_hd__dfxbp_1_0.CLK 0.0158f
C1123 a_15522_4547# a_6208_2817# 0
C1124 a_4595_14775# VDPWR 0.02521f
C1125 a_17521_23241# a_16823_22875# 0.19462f
C1126 a_17605_23241# VDPWR 0.00627f
C1127 a_17425_5473# a_16485_5729# 0.13858f
C1128 a_7113_13395# a_7831_14003# 0.00223f
C1129 a_4423_5299# a_3229_5051# 0.21187f
C1130 a_11255_13773# a_9715_11297# 0.00488f
C1131 a_3229_5051# VDPWR 1.39976f
C1132 a_15239_23241# VDPWR 0.19826f
C1133 a_6261_5409# VDPWR 0
C1134 a_10025_1793# a_10289_1793# 0
C1135 a_8193_13753# a_6281_11907# 0.00288f
C1136 a_6087_14735# a_4837_16089# 0.29394f
C1137 sky130_fd_sc_hd__dfxbp_1_1.CLK a_10933_22879# 0
C1138 uo_out[0] sky130_fd_sc_hd__inv_12_0.A 0
C1139 a_23731_14309# a_24962_14701# 0
C1140 a_17521_23241# a_17689_23143# 0.31062f
C1141 a_16847_4529# a_6208_2817# 0
C1142 a_10382_23245# sky130_fd_sc_hd__dfxbp_1_0.Q_N 0
C1143 a_7173_15235# a_6635_15235# 0.08414f
C1144 a_14908_5467# VDPWR 0.21933f
C1145 a_12823_4553# a_12655_4553# 0
C1146 a_11888_1767# a_12227_2049# 0.04737f
C1147 a_6127_13769# a_4913_13781# 0
C1148 a_9223_1793# a_10121_1793# 0
C1149 sky130_fd_sc_hd__dfxbp_1_1.Q_N sky130_fd_sc_hd__dfxbp_1_2.CLK 0.15319f
C1150 sky130_fd_sc_hd__dfxbp_1_4.CLK sky130_fd_sc_hd__dfxbp_1_4.Q_N 0.01744f
C1151 a_10975_23147# sky130_fd_sc_hd__dfxbp_1_1.CLK 0
C1152 a_16454_4503# a_15188_4913# 0
C1153 a_7221_1787# a_8073_1793# 0
C1154 a_16033_1793# a_6208_2817# 0
C1155 a_6238_6077# a_14561_4913# 0
C1156 sky130_fd_sc_hd__dfxbp_1_6.Q_N a_18671_30311# 0.12801f
C1157 a_10841_12931# a_10995_12931# 0.00401f
C1158 a_6389_13769# a_6862_13645# 0.24537f
C1159 a_18667_34259# a_18667_34470# 0.31062f
C1160 a_6429_5409# a_5363_5043# 0.04534f
C1161 a_18689_26867# sky130_fd_sc_hd__dfxbp_1_7.CLK 0
C1162 a_18671_29731# a_18671_29942# 0.31062f
C1163 a_9317_5049# a_14432_4521# 0
C1164 VDPWR a_2676_1791# 0.22056f
C1165 a_18371_4938# VDPWR 0.15241f
C1166 sky130_fd_sc_hd__dfxbp_1_9.Q_N a_18667_33834# 0
C1167 a_10121_1793# a_10289_1793# 0
C1168 a_10807_23245# a_10933_22879# 0.00617f
C1169 a_4903_15345# VDPWR 0.38131f
C1170 a_4383_2153# a_4215_2153# 0
C1171 a_14541_22875# sky130_fd_sc_hd__dfxbp_1_2.Q_N 0.0011f
C1172 a_13186_4919# VDPWR 0.02137f
C1173 a_9619_16343# a_9703_16093# 0.07445f
C1174 a_18667_25006# a_18693_24621# 0.03733f
C1175 a_18663_27120# a_19055_27518# 0
C1176 a_18671_29731# a_19063_29704# 0
C1177 a_9943_22879# a_10109_22879# 0.96835f
C1178 a_4763_14775# a_4903_15345# 0.00327f
C1179 a_4755_13107# a_4505_13107# 0.02504f
C1180 sky130_fd_sc_hd__dfxbp_1_5.Q_N sky130_fd_sc_hd__dfxbp_1_7.CLK 0.15244f
C1181 a_6429_5043# a_6792_5043# 0.00985f
C1182 a_6208_2817# a_12113_2159# 0
C1183 a_14432_4521# a_12823_4919# 0
C1184 a_10975_23147# a_10807_23245# 0.31062f
C1185 a_9317_5049# a_13709_4553# 0.03427f
C1186 a_12430_4527# a_12559_4919# 0.00792f
C1187 a_18671_29731# VDPWR 0.51547f
C1188 sky130_fd_sc_hd__dfxbp_1_1.CLK VDPWR 0.2726f
C1189 a_2187_1765# VDPWR 1.68729f
C1190 a_11888_1767# a_12113_1793# 0.00487f
C1191 VDPWR a_6071_2153# 0
C1192 sky130_fd_sc_hd__dfxbp_1_1.CLK a_9160_23197# 0.20774f
C1193 a_2175_5417# a_2217_5025# 0
C1194 a_21506_16181# VDPWR 0.42312f
C1195 a_8263_5049# VDPWR 0
C1196 a_11255_13773# a_10993_13773# 0
C1197 a_10160_4571# a_10553_4597# 0.02283f
C1198 a_6238_6077# a_10261_5837# 0
C1199 a_9705_12861# a_11728_13649# 0.00327f
C1200 a_23511_14335# a_23133_17137# 0.05287f
C1201 a_14152_5441# a_14432_4521# 0
C1202 a_14729_22875# a_14814_23241# 0.03733f
C1203 a_6238_6077# a_12378_4553# 0
C1204 a_15323_23241# a_14541_22875# 0
C1205 a_16402_4529# a_14771_4803# 0
C1206 a_4329_2043# a_4746_2153# 0.06611f
C1207 a_7221_1787# a_7032_2153# 0
C1208 sky130_fd_sc_hd__dfxbp_1_3.CLK a_12736_22983# 0
C1209 a_14825_4547# a_14771_4803# 0.00386f
C1210 a_9715_11297# a_9453_13111# 0
C1211 sky130_fd_sc_hd__inv_2_0.A a_18667_33731# 0
C1212 a_10235_2049# a_11175_1793# 0.13739f
C1213 a_2259_2047# a_2313_2157# 0.03622f
C1214 VDPWR a_18693_33761# 0.00347f
C1215 a_15431_5467# a_14771_4803# 0
C1216 a_14982_22987# VDPWR 0.19114f
C1217 a_4765_11543# a_4505_13107# 0
C1218 sky130_fd_sc_hd__dfxbp_1_9.Q_N a_18671_29942# 0
C1219 a_7173_15235# a_9501_13813# 0
C1220 a_14377_5467# VDPWR 0
C1221 VDPWR a_10807_23245# 0.19828f
C1222 a_17521_23241# sky130_fd_sc_hd__dfxbp_1_4.CLK 0
C1223 VDPWR a_8073_2159# 0
C1224 a_16471_17161# a_15641_17149# 0
C1225 a_8377_5305# a_8794_5049# 0.03016f
C1226 a_18667_33966# a_18667_33731# 0.27314f
C1227 a_6335_2153# a_6167_2153# 0
C1228 a_5975_12927# a_6057_12927# 0.00517f
C1229 a_14152_5441# a_13709_4553# 0
C1230 a_4329_2043# a_5890_1787# 0
C1231 a_7986_5049# a_6375_5299# 0
C1232 a_6281_2043# a_7944_1767# 0.0035f
C1233 a_18667_31552# a_18693_31893# 0
C1234 sky130_fd_sc_hd__dfxbp_1_7.Q a_18663_27756# 0.00393f
C1235 a_9705_12861# a_10675_14767# 0.21988f
C1236 sky130_fd_sc_hd__dfxbp_1_3.CLK a_12483_22871# 0
C1237 a_4763_14525# a_4839_12857# 0
C1238 a_9705_12861# a_9379_14779# 0.00442f
C1239 a_10869_11939# a_10955_11939# 0.00658f
C1240 a_8687_22875# VDPWR 0
C1241 a_6238_6077# a_14432_4521# 0
C1242 a_9781_10553# a_11147_11911# 0.43338f
C1243 a_7113_13395# a_7927_14003# 0.00121f
C1244 a_3990_1761# a_4383_2153# 0.02301f
C1245 a_11888_1767# a_6208_2817# 0.00211f
C1246 VDPWR a_24774_14701# 0.22575f
C1247 a_12419_5825# a_12533_5715# 0
C1248 sky130_fd_sc_hd__dfxbp_1_5.CLK a_18667_24676# 0.01408f
C1249 a_11175_1793# a_11836_1793# 0.05012f
C1250 a_4847_14525# a_4849_11293# 0.00506f
C1251 a_5942_1761# a_6281_2043# 0.04737f
C1252 a_6238_6077# a_15188_4913# 0
C1253 a_4847_14525# a_5851_13769# 0
C1254 a_10025_2159# a_9844_1793# 0
C1255 sky130_fd_sc_hd__dfxbp_1_9.Q_N VDPWR 0.60837f
C1256 a_8136_23241# a_9943_22879# 0
C1257 a_8561_23241# sky130_fd_sc_hd__dfxbp_1_0.Q_N 0.09273f
C1258 sky130_fd_sc_hd__dfxbp_1_3.CLK VDPWR 0.27262f
C1259 a_13520_4919# VDPWR 0
C1260 a_2187_1765# a_3010_1791# 0
C1261 a_4032_5043# a_4213_5409# 0
C1262 a_9705_12861# a_10799_13773# 0
C1263 VDPWR a_4215_1787# 0
C1264 a_4847_14525# a_4625_15373# 0.00215f
C1265 a_6389_13769# a_4913_13781# 0
C1266 a_18663_27252# sky130_fd_sc_hd__dfxbp_1_7.CLK 0
C1267 a_8038_5023# a_8167_5049# 0.00758f
C1268 a_4849_11293# a_6087_14735# 0.00179f
C1269 a_9781_10553# a_9771_12117# 0.0298f
C1270 a_4423_5299# a_5984_5043# 0
C1271 a_14729_22875# sky130_fd_sc_hd__dfxbp_1_2.Q_N 0
C1272 a_6087_14735# a_5851_13769# 0
C1273 a_23511_14701# a_23511_14335# 0.00987f
C1274 a_10550_22991# a_10933_22879# 0
C1275 a_5984_5043# VDPWR 0.16491f
C1276 a_6238_6077# a_12323_5825# 0
C1277 a_9705_12861# a_8193_13753# 0.00341f
C1278 a_6238_6077# a_13709_4553# 0
C1279 a_4423_5299# a_5363_5043# 0.13739f
C1280 sky130_fd_sc_hd__dfxbp_1_5.CLK a_17605_23241# 0
C1281 a_5363_5043# VDPWR 1.39451f
C1282 a_18667_34839# a_18667_33731# 0
C1283 a_14380_4547# a_14561_4913# 0
C1284 a_6429_5409# a_6792_5409# 0.00847f
C1285 sky130_fd_sc_hd__dfxbp_1_9.Q sky130_fd_sc_hd__dfxbp_1_9.Q_N 0.15089f
C1286 a_14930_2159# VDPWR 0
C1287 a_7221_1787# a_7892_1793# 0.05007f
C1288 a_18667_31449# a_18667_32188# 0.03218f
C1289 a_2187_1765# a_2145_2157# 0
C1290 a_20109_17157# a_20877_17147# 0.10376f
C1291 a_6238_6077# a_12419_5825# 0
C1292 a_14657_4913# VDPWR 0
C1293 a_14561_4913# a_14825_4913# 0
C1294 a_18371_4938# a_9317_5049# 0.24923f
C1295 a_4849_11293# a_4637_10577# 0
C1296 a_11255_13773# a_10887_13773# 0
C1297 a_10717_13773# a_11255_13773# 0.07901f
C1298 a_6238_6077# a_10080_5471# 0.00331f
C1299 a_7113_13395# a_7999_14003# 0.00205f
C1300 a_8167_5049# a_7315_5043# 0
C1301 a_23731_14309# a_24774_14701# 0.00253f
C1302 a_12823_4553# a_6208_2817# 0
C1303 a_2187_1765# a_6071_1787# 0
C1304 a_4505_13107# a_4627_12141# 0.00144f
C1305 a_10975_23147# a_10550_22991# 0
C1306 a_9705_12861# a_9779_13785# 0.44871f
C1307 a_18671_29731# a_18671_29203# 0.04808f
C1308 a_2187_1765# a_5080_1787# 0
C1309 uo_out[6] uo_out[7] 0.03102f
C1310 a_7749_14003# VDPWR 0.13648f
C1311 a_1868_1791# a_2187_1765# 0.0073f
C1312 a_18371_4938# a_16793_4785# 0
C1313 a_14596_1793# VDPWR 0.21794f
C1314 a_10953_14739# a_11255_13773# 0.00214f
C1315 a_7944_1767# VDPWR 0.34956f
C1316 sky130_fd_sc_hd__dfxbp_1_9.Q_N a_18667_31977# 0.12218f
C1317 a_15239_23241# sky130_fd_sc_hd__dfxbp_1_2.Q_N 0
C1318 a_1950_5025# a_2079_5051# 0.00758f
C1319 a_18113_17153# sky130_fd_sc_hd__dfxbp_1_0.CLK 0.03683f
C1320 a_10121_2159# VDPWR 0
C1321 a_7113_13395# a_6329_12927# 0
C1322 a_16902_5839# a_14491_5723# 0
C1323 a_9943_22879# a_10297_22879# 0.06222f
C1324 a_8377_5305# a_9128_5415# 0.00696f
C1325 a_9223_1793# a_10289_2159# 0.04534f
C1326 a_9769_15349# a_11728_13649# 0
C1327 a_7221_1787# a_8337_2159# 0.04534f
C1328 a_16402_4529# a_6208_2817# 0
C1329 a_12039_15239# a_11777_15239# 0
C1330 VDPWR a_11728_13649# 0.16015f
C1331 a_13186_4919# a_12823_4919# 0.00847f
C1332 a_16657_22875# a_16823_22875# 0.96835f
C1333 a_5942_1761# VDPWR 0.35234f
C1334 a_6208_2817# a_14825_4547# 0
C1335 a_3990_1761# a_4119_1787# 0.00758f
C1336 a_10109_22879# a_8729_23143# 0
C1337 a_9587_13813# a_9779_13785# 0.00222f
C1338 a_10235_2049# a_9896_1767# 0.04737f
C1339 a_20109_17157# a_21491_17145# 0
C1340 a_18667_25510# VDPWR 0.1998f
C1341 a_18553_4938# a_18625_4938# 0
C1342 a_9713_14529# a_12039_15239# 0
C1343 a_9705_12861# a_9621_12861# 0.00208f
C1344 a_6261_5409# a_6238_6077# 0
C1345 sky130_fd_sc_hd__dfxbp_1_7.Q_N sky130_fd_sc_hd__dfxbp_1_7.CLK 0.0174f
C1346 a_17689_23143# a_16657_22875# 0.04808f
C1347 sky130_fd_sc_hd__dfxbp_1_5.Q_N a_18667_25879# 0.12801f
C1348 a_4713_12141# a_4627_12141# 0.00658f
C1349 a_15711_4547# a_17210_4529# 0.08907f
C1350 a_4119_1787# a_4383_1787# 0
C1351 a_16243_2049# a_16994_1793# 0.00682f
C1352 a_4847_14525# a_6635_15235# 0.17824f
C1353 a_18663_27017# a_18689_27047# 0.0027f
C1354 a_10550_22991# VDPWR 0.19115f
C1355 a_12194_5433# VDPWR 0.35512f
C1356 a_4505_13107# a_4587_13107# 0.00641f
C1357 a_12655_4553# VDPWR 0
C1358 ui_in[0] a_24407_14651# 0.00109f
C1359 a_15323_23241# a_15239_23241# 0.00851f
C1360 a_14982_22987# a_14814_23241# 0.23992f
C1361 a_14908_5467# a_6238_6077# 0
C1362 a_8283_2049# a_8169_2159# 0
C1363 a_20109_17157# sky130_fd_sc_hd__dfxbp_1_0.CLK 0.01979f
C1364 a_6087_14735# a_6635_15235# 0.08954f
C1365 a_9769_15349# a_10675_14767# 0.0039f
C1366 a_18667_33731# a_18667_31354# 0
C1367 a_13840_1767# a_14233_2159# 0.02301f
C1368 a_10675_14767# VDPWR 0.2094f
C1369 sky130_fd_sc_hd__dfxbp_1_3.Q_N a_15838_23197# 0.12801f
C1370 a_18667_24771# a_18663_26922# 0
C1371 a_9379_14779# a_9769_15349# 0.00566f
C1372 a_9379_14779# VDPWR 0.54114f
C1373 a_12295_22871# a_12568_23237# 0.07715f
C1374 a_6057_12927# VDPWR 0
C1375 a_12430_4527# a_12378_4553# 0.1439f
C1376 a_6944_13645# a_6281_11907# 0
C1377 a_9371_13111# a_9501_13813# 0.00115f
C1378 a_6208_2817# a_8700_2159# 0
C1379 a_6862_13645# a_6329_12927# 0.10646f
C1380 a_15119_1793# a_16033_1793# 0
C1381 a_4746_1787# a_4383_1787# 0.00985f
C1382 a_18693_31299# a_18667_31354# 0.0967f
C1383 sky130_fd_sc_hd__dfxbp_1_8.Q_N a_19059_33811# 0.00188f
C1384 a_9705_12861# a_9621_13111# 0.08134f
C1385 a_9769_15349# a_10799_13773# 0.0035f
C1386 a_18371_4938# a_6238_6077# 0.00367f
C1387 a_8794_5049# VDPWR 0.21794f
C1388 a_10799_13773# VDPWR 0
C1389 a_12281_1793# a_12227_2049# 0.00386f
C1390 a_16583_4529# a_6208_2817# 0
C1391 a_15904_1767# a_16129_1793# 0.00487f
C1392 a_14380_4547# a_14432_4521# 0.1439f
C1393 a_6238_6077# a_13186_4919# 0
C1394 a_15365_22875# a_15239_23241# 0.00617f
C1395 sky130_fd_sc_hd__dfxbp_1_3.CLK a_14814_23241# 0
C1396 a_4329_2043# a_5269_1787# 0.13739f
C1397 a_12227_2049# VDPWR 0.45036f
C1398 a_9769_15349# a_8193_13753# 0.00137f
C1399 a_11810_13649# a_11728_13649# 0.00477f
C1400 a_14432_4521# a_14825_4913# 0.02301f
C1401 a_11255_13773# a_11195_12931# 0.20048f
C1402 a_8193_13753# VDPWR 2.47419f
C1403 a_14771_4803# VDPWR 0.4846f
C1404 a_11411_5471# a_12323_5459# 0
C1405 a_15188_4913# a_14825_4913# 0.00847f
C1406 a_7221_1787# a_5269_1787# 0
C1407 a_6389_13769# a_5933_13769# 0
C1408 a_18667_25006# a_19059_24851# 0.00553f
C1409 a_4765_11293# a_4515_11543# 0.00723f
C1410 a_14377_5467# a_14152_5441# 0.00487f
C1411 a_13077_23237# a_12993_23237# 0.00851f
C1412 a_6792_5409# VDPWR 0.02103f
C1413 a_17011_22875# a_16657_22875# 0.06222f
C1414 a_1950_5025# a_1898_5051# 0.1439f
C1415 a_14380_4547# a_13709_4553# 0.05007f
C1416 a_9769_15349# a_9779_13785# 0.11601f
C1417 a_11671_15239# VDPWR 0.00152f
C1418 a_14179_2049# VDPWR 0.45001f
C1419 a_15407_23143# sky130_fd_sc_hd__dfxbp_1_4.Q_N 0
C1420 a_9779_13785# VDPWR 0.75079f
C1421 a_14982_22987# sky130_fd_sc_hd__dfxbp_1_2.Q_N 0
C1422 a_6238_6077# a_8263_5049# 0
C1423 a_13709_4553# a_14825_4913# 0.04534f
C1424 a_5269_1787# a_5890_1787# 0.0504f
C1425 a_7173_15235# a_6281_11907# 0.09952f
C1426 a_5942_1761# a_6071_1787# 0.00758f
C1427 sky130_fd_sc_hd__inv_2_0.A a_18667_33966# 0
C1428 a_18742_16187# VDPWR 0.43871f
C1429 a_9556_17271# a_9369_16343# 0
C1430 a_18667_24874# a_18663_27017# 0
C1431 a_17425_5473# a_18371_4938# 0.08028f
C1432 a_3229_5051# a_2706_5051# 0
C1433 a_7697_22875# sky130_fd_sc_hd__dfxbp_1_0.Q_N 0.11931f
C1434 a_6281_2043# a_6208_2817# 0.00307f
C1435 a_6021_13769# a_4913_13781# 0.00104f
C1436 a_6375_5299# a_6261_5043# 0
C1437 a_18667_31684# a_19059_31529# 0.00553f
C1438 a_12281_1793# a_12113_1793# 0
C1439 a_4839_12857# a_4915_10549# 0.00242f
C1440 a_12113_1793# VDPWR 0
C1441 sky130_fd_sc_hd__dfxbp_1_4.CLK a_16657_22875# 0.25126f
C1442 a_9579_12145# a_9771_12117# 0
C1443 a_14377_5467# a_6238_6077# 0
C1444 a_9621_12861# VDPWR 0.00415f
C1445 a_12295_22871# a_14375_22875# 0
C1446 sky130_fd_sc_hd__dfxbp_1_3.CLK sky130_fd_sc_hd__dfxbp_1_2.Q_N 0.15244f
C1447 a_24234_14385# a_24318_14385# 0.0296f
C1448 a_17264_22987# a_17222_22875# 0
C1449 a_17254_16187# VDPWR 0.46715f
C1450 a_10357_5837# a_10525_5837# 0
C1451 a_18667_32557# sky130_fd_sc_hd__dfxbp_1_9.Q_N 0.12801f
C1452 a_14982_22987# a_15323_23241# 0
C1453 a_4915_10549# a_4515_11543# 0
C1454 a_9128_5415# VDPWR 0
C1455 a_10297_22879# a_8729_23143# 0
C1456 sky130_fd_sc_hd__dfxbp_1_7.Q a_18663_26922# 0
C1457 a_16297_2159# VDPWR 0.00966f
C1458 a_14596_2159# a_14233_2159# 0.00847f
C1459 a_23133_17137# a_24407_14651# 0
C1460 a_18667_31449# a_18667_31684# 0.27314f
C1461 a_14432_4521# a_13473_5459# 0.00135f
C1462 a_6238_6077# a_24774_14701# 0
C1463 a_9317_5049# a_12194_5433# 0
C1464 a_10888_5837# VDPWR 0.02103f
C1465 sky130_fd_sc_hd__inv_2_0.A a_18667_34839# 0.20332f
C1466 sky130_fd_sc_hd__dfxbp_1_1.Q_N a_10382_23245# 0.04247f
C1467 a_5975_12927# a_4505_13107# 0
C1468 a_6238_6077# a_13520_4919# 0
C1469 a_12295_22871# a_12129_22871# 0.96835f
C1470 a_6329_12927# a_4913_13781# 0.0204f
C1471 a_18693_25215# a_18667_24676# 0
C1472 a_9371_13111# a_9771_12117# 0
C1473 a_12039_15239# a_11501_15239# 0.08415f
C1474 sky130_fd_sc_hd__dfxbp_1_7.Q_N a_18667_25879# 0
C1475 a_8136_23241# a_8231_23241# 0.00772f
C1476 a_9621_13111# VDPWR 0.33272f
C1477 a_14982_22987# a_15365_22875# 0
C1478 a_4837_16089# a_4915_10549# 0.01618f
C1479 a_13709_4553# a_13473_5459# 0.00111f
C1480 ui_in[2] ui_in[1] 0.03102f
C1481 a_6238_6077# a_5363_5043# 0.00183f
C1482 a_4505_13107# a_4513_14775# 0
C1483 a_9369_16343# a_9703_16093# 0.16891f
C1484 a_15188_4547# a_13709_4553# 0.08907f
C1485 a_12281_1793# a_6208_2817# 0
C1486 a_1920_1765# a_2145_1791# 0.00487f
C1487 sky130_fd_sc_hd__dfxbp_1_5.CLK a_18667_25510# 0
C1488 a_3040_5051# VDPWR 0
C1489 a_16454_4503# a_14771_4803# 0.00271f
C1490 a_9715_11297# a_11728_13649# 0
C1491 a_6208_2817# VDPWR 0.49985f
C1492 a_6208_2817# a_9034_2159# 0
C1493 a_4032_5043# a_2289_5307# 0
C1494 a_6238_6077# a_14657_4913# 0
C1495 a_2049_1791# VDPWR 0.00125f
C1496 a_9781_10553# a_9705_12861# 0.00242f
C1497 a_23761_14335# a_23511_14335# 0.08551f
C1498 a_9317_5049# a_8794_5049# 0
C1499 a_18667_24676# a_18693_24621# 0.0967f
C1500 sky130_fd_sc_hd__dfxbp_1_6.Q_N a_18663_28125# 0
C1501 ui_in[1] a_24962_14701# 0.03406f
C1502 a_18689_26867# VDPWR 0.07703f
C1503 a_18671_29731# a_18671_29108# 0.03136f
C1504 a_24234_14385# a_24241_14651# 0.13413f
C1505 a_18671_29306# a_18697_29053# 0
C1506 a_9713_14529# a_9501_13813# 0
C1507 a_13969_2159# a_14233_2159# 0
C1508 a_6261_5043# a_6036_5017# 0.00487f
C1509 a_16033_2159# VDPWR 0
C1510 a_4503_16339# a_4837_16089# 0.16891f
C1511 a_4423_5299# a_5174_5043# 0.00682f
C1512 a_18663_27756# a_19055_27518# 0.00617f
C1513 a_8231_23241# a_8051_22875# 0.00123f
C1514 a_5174_5043# VDPWR 0
C1515 a_9317_5049# a_14771_4803# 0
C1516 a_19059_31950# a_18667_32188# 0.00617f
C1517 sky130_fd_sc_hd__dfxbp_1_0.Q_N a_8304_22987# 0.05782f
C1518 a_15365_22875# sky130_fd_sc_hd__dfxbp_1_3.CLK 0
C1519 a_12533_5715# a_12194_5433# 0.04737f
C1520 a_17345_17163# a_18113_17153# 0.1017f
C1521 a_24241_14651# a_24318_14385# 0.01352f
C1522 a_9896_1767# a_9844_1793# 0.1439f
C1523 a_5975_12927# a_5809_14763# 0
C1524 sky130_fd_sc_hd__dfxbp_1_5.Q_N VDPWR 0.60771f
C1525 a_3229_5051# a_2289_5307# 0.13963f
C1526 a_24407_14651# sky130_fd_sc_hd__dfxbp_1_0.CLK 0
C1527 a_6629_15387# a_4753_16339# 0
C1528 a_7113_13395# a_6862_13645# 0.10945f
C1529 a_6375_5299# a_7126_5409# 0.00696f
C1530 a_13592_23193# a_13161_23139# 0.10805f
C1531 a_4309_5043# a_2217_5025# 0
C1532 a_11501_15239# a_11979_13399# 0
C1533 a_6127_13769# a_4903_15345# 0
C1534 a_6208_2817# a_6698_2153# 0
C1535 a_9715_11297# a_10675_14767# 0.10553f
C1536 a_23731_14309# a_6208_2817# 0
C1537 a_14432_4521# a_14491_5723# 0
C1538 a_9379_14779# a_9715_11297# 0.00146f
C1539 a_10357_5837# a_10132_5445# 0.00559f
C1540 a_15188_4913# a_14491_5723# 0
C1541 a_21506_16181# a_20384_16179# 0.1017f
C1542 a_14375_22875# a_16657_22875# 0
C1543 a_5809_14763# a_4513_14775# 0
C1544 a_4637_10577# a_4765_11543# 0
C1545 a_11255_13773# a_9703_16093# 0.00515f
C1546 a_11255_13773# a_12697_14007# 0
C1547 a_6238_6077# a_12194_5433# 0.0051f
C1548 sky130_fd_sc_hd__dfxbp_1_6.Q_N a_18671_29942# 0.09273f
C1549 a_9371_13111# a_6281_11907# 0
C1550 a_18671_29731# sky130_fd_sc_hd__dfxbp_1_9.CLK 0.12322f
C1551 a_14179_2049# a_14065_1793# 0
C1552 a_9715_11297# a_10799_13773# 0
C1553 a_4755_12857# VDPWR 0.00415f
C1554 a_13709_4553# a_14491_5723# 0.00129f
C1555 a_14908_5467# a_13473_5459# 0.08907f
C1556 a_18671_29438# VDPWR 0.25525f
C1557 a_15904_1767# a_16297_1793# 0.02283f
C1558 a_9943_22879# sky130_fd_sc_hd__dfxbp_1_1.CLK 0.25091f
C1559 sky130_fd_sc_hd__dfxbp_1_6.Q_N a_19063_29704# 0.00125f
C1560 a_12587_5825# a_11439_4597# 0
C1561 a_16146_5447# a_16539_5839# 0.02301f
C1562 a_3199_1791# a_3010_2157# 0
C1563 a_9317_5049# a_9128_5415# 0
C1564 a_17096_23241# sky130_fd_sc_hd__dfxbp_1_4.Q_N 0.04247f
C1565 a_14375_22875# a_13161_23139# 0
C1566 a_4849_11293# a_4765_11293# 0.00206f
C1567 sky130_fd_sc_hd__dfxbp_1_6.Q_N VDPWR 0.60833f
C1568 a_4905_12113# a_4915_10549# 0.0298f
C1569 a_6238_6077# a_8794_5049# 0
C1570 a_9715_11297# a_9779_13785# 0.26133f
C1571 uio_in[6] uio_in[5] 0.03102f
C1572 a_18742_16187# a_19235_17155# 0
C1573 a_10553_4597# VDPWR 0.27571f
C1574 sky130_fd_sc_hd__dfxbp_1_1.Q_N a_8561_23241# 0
C1575 a_9381_11547# a_9493_12145# 0
C1576 a_18663_28125# sky130_fd_sc_hd__dfxbp_1_7.Q_N 0.12801f
C1577 a_16243_2049# a_16660_1793# 0.03016f
C1578 a_3229_5051# a_4840_5043# 0.08907f
C1579 sky130_fd_sc_hd__dfxbp_1_2.CLK a_10382_23245# 0
C1580 a_5895_14763# VDPWR 0
C1581 a_4505_13107# VDPWR 0.54084f
C1582 a_18667_25299# a_18663_26922# 0
C1583 a_16454_4503# a_6208_2817# 0
C1584 a_14179_2049# a_14930_1793# 0.00682f
C1585 a_6238_6077# a_14771_4803# 0
C1586 a_13167_1793# a_12978_2159# 0
C1587 a_12587_5459# a_11439_4597# 0
C1588 a_18693_33581# a_18693_33761# 0.00123f
C1589 a_15711_4547# a_15522_4913# 0
C1590 a_4839_12857# a_4515_11543# 0
C1591 a_10235_2049# a_10121_2159# 0
C1592 a_6281_2043# a_6335_1787# 0.00386f
C1593 a_14825_4547# a_14657_4547# 0
C1594 a_23133_17137# a_22365_17147# 0.10345f
C1595 a_12129_22871# a_13161_23139# 0.04808f
C1596 a_9781_10553# VDPWR 0.67675f
C1597 a_20877_17147# a_22365_17147# 0
C1598 a_9943_22879# a_10807_23245# 0.03218f
C1599 sky130_fd_sc_hd__dfxbp_1_1.Q_N a_12568_23237# 0
C1600 a_4637_10577# a_4627_12141# 0
C1601 a_6792_5409# a_6238_6077# 0
C1602 VDPWR a_18663_27252# 0.25541f
C1603 a_4839_12857# a_4635_13809# 0.00246f
C1604 a_10869_11939# a_11147_11911# 0.11706f
C1605 ui_in[0] a_23133_17137# 0.01883f
C1606 a_18128_16189# VDPWR 0.35113f
C1607 a_4084_5017# a_4213_5043# 0.00758f
C1608 a_18667_31552# sky130_fd_sc_hd__dfxbp_1_9.Q_N 0.05782f
C1609 a_9621_12861# a_9715_11297# 0
C1610 a_15431_5467# a_16146_5447# 0.11891f
C1611 sky130_fd_sc_hd__dfxbp_1_9.CLK sky130_fd_sc_hd__dfxbp_1_9.Q_N 0.0174f
C1612 a_11411_5471# a_12142_5459# 0.04968f
C1613 a_14561_4547# a_14432_4521# 0.00758f
C1614 sky130_fd_sc_hd__dfxbp_1_6.Q_N a_18667_31977# 0
C1615 a_2175_5417# VDPWR 0
C1616 a_6944_13645# VDPWR 0.0014f
C1617 a_16793_4785# a_6208_2817# 0
C1618 sky130_fd_sc_hd__dfxbp_1_8.Q_N sky130_fd_sc_hd__dfxbp_1_9.Q_N 0
C1619 a_14657_4913# a_14825_4913# 0
C1620 a_5851_13769# a_4915_10549# 0.00192f
C1621 a_4849_11293# a_4915_10549# 0.00633f
C1622 a_14908_5467# a_14491_5723# 0.03016f
C1623 a_6208_2817# a_7032_1787# 0
C1624 a_18693_33581# sky130_fd_sc_hd__dfxbp_1_9.Q_N 0
C1625 a_10869_11939# a_9771_12117# 0.18489f
C1626 a_13119_22871# a_12993_23237# 0.00617f
C1627 a_4839_12857# a_4837_16089# 0.4639f
C1628 a_4713_12141# VDPWR 0.00297f
C1629 a_9034_1793# VDPWR 0
C1630 a_18689_27461# VDPWR 0.00629f
C1631 sky130_fd_sc_hd__dfxbp_1_0.Q_N a_7863_22875# 0.5114f
C1632 a_6208_2817# a_14065_1793# 0
C1633 sky130_fd_sc_hd__dfxbp_1_7.Q_N a_18671_29942# 0
C1634 a_10025_1793# VDPWR 0.00116f
C1635 a_9491_15377# a_9501_13813# 0
C1636 uo_out[2] uo_out[1] 0.03102f
C1637 a_5809_14763# VDPWR 0.2094f
C1638 a_21491_17145# a_22365_17147# 0.1036f
C1639 a_14561_4547# a_13709_4553# 0
C1640 a_4084_5017# a_2706_5417# 0
C1641 a_14377_5467# a_13473_5459# 0
C1642 uo_out[7] uio_out[0] 0.03102f
C1643 a_18667_25006# a_18667_24771# 0.27314f
C1644 a_10132_5445# a_10261_5471# 0.00758f
C1645 a_6375_5299# a_6036_5017# 0.04737f
C1646 a_4084_5017# a_4477_5409# 0.02301f
C1647 a_6389_13769# a_4903_15345# 0
C1648 a_14432_4521# a_12769_4809# 0.00352f
C1649 a_9621_13111# a_9715_11297# 0
C1650 a_9128_5415# a_6238_6077# 0
C1651 a_16486_16197# VDPWR 0.35942f
C1652 a_10717_13773# a_11728_13649# 0
C1653 ui_in[1] a_24774_14701# 0.29195f
C1654 VDPWR a_6335_1787# 0.18611f
C1655 a_1920_1765# a_2187_1765# 0.08244f
C1656 a_18671_29438# a_18671_29203# 0.27314f
C1657 a_4503_16339# a_4625_15373# 0.00144f
C1658 a_16129_1793# a_16297_1793# 0
C1659 a_9779_13785# a_10993_13773# 0
C1660 sky130_fd_sc_hd__dfxbp_1_7.Q_N VDPWR 0.60896f
C1661 a_6238_6077# a_10888_5837# 0.00192f
C1662 a_12865_14007# a_12039_15239# 0
C1663 a_22365_17147# sky130_fd_sc_hd__dfxbp_1_0.CLK 0.02379f
C1664 a_10953_14739# a_11728_13649# 0
C1665 sky130_fd_sc_hd__dfxbp_1_4.Q_N VDPWR 0.60276f
C1666 a_7173_15235# VDPWR 0.83685f
C1667 a_18689_26867# a_18663_27120# 0
C1668 a_18663_27545# sky130_fd_sc_hd__dfxbp_1_7.CLK 0
C1669 uio_oe[5] uio_oe[6] 0.03102f
C1670 a_12865_14007# a_12615_14007# 0.00876f
C1671 a_4084_5017# a_2217_5025# 0.0021f
C1672 a_13709_4553# a_12769_4809# 0.13741f
C1673 a_23511_14701# ui_in[0] 0.0029f
C1674 sky130_fd_sc_hd__dfxbp_1_6.Q_N a_18671_29203# 0.11931f
C1675 ui_in[0] sky130_fd_sc_hd__dfxbp_1_0.CLK 0.35686f
C1676 sky130_fd_sc_hd__dfxbp_1_5.Q_N sky130_fd_sc_hd__dfxbp_1_5.CLK 0.01521f
C1677 a_14930_1793# a_6208_2817# 0
C1678 a_17210_4529# a_16847_4529# 0.00985f
C1679 a_10121_1793# VDPWR 0
C1680 a_6862_13645# a_4913_13781# 0
C1681 a_15407_23143# a_16657_22875# 0
C1682 sky130_fd_sc_hd__dfxbp_1_5.Q_N a_18663_27120# 0
C1683 a_9705_12861# a_9371_13111# 0.16952f
C1684 a_12430_4527# a_12194_5433# 0
C1685 a_6238_6077# a_6208_2817# 0.91673f
C1686 a_10717_13773# a_10675_14767# 0
C1687 a_12655_4553# a_12430_4527# 0.00487f
C1688 sky130_fd_sc_hd__dfxbp_1_1.CLK a_8729_23143# 0.12322f
C1689 a_9381_11547# a_9631_11297# 0.00723f
C1690 a_13186_4553# a_13709_4553# 0
C1691 a_9369_16343# a_9619_16343# 0.02504f
C1692 a_15119_1793# VDPWR 1.38901f
C1693 a_12295_22871# a_11406_23201# 0
C1694 a_9943_22879# a_10550_22991# 0.14145f
C1695 a_18693_25215# a_18667_25510# 0.00851f
C1696 a_6792_5043# VDPWR 0.218f
C1697 a_9503_10581# VDPWR 0.43224f
C1698 a_10953_14739# a_10675_14767# 0.1109f
C1699 a_18667_31449# a_18671_29306# 0
C1700 sky130_fd_sc_hd__dfxbp_1_1.Q_N a_12129_22871# 0.0031f
C1701 a_10953_14739# a_9379_14779# 0
C1702 a_19059_34232# a_18667_33834# 0
C1703 a_10499_4853# a_11439_4597# 0.14008f
C1704 a_16539_5473# a_16146_5447# 0.02283f
C1705 a_14377_5467# a_14491_5723# 0
C1706 a_6429_5043# a_6261_5043# 0
C1707 a_10717_13773# a_10799_13773# 0.00578f
C1708 a_12865_14007# a_11979_13399# 0.00205f
C1709 a_9713_14529# a_9577_15377# 0
C1710 a_4839_12857# a_4905_12113# 0.04364f
C1711 a_13840_1767# a_13788_1793# 0.1439f
C1712 a_21506_16181# a_9556_17271# 0
C1713 sky130_fd_sc_hd__dfxbp_1_2.CLK a_12568_23237# 0
C1714 a_14771_4803# a_14825_4913# 0.03622f
C1715 a_6208_2817# a_16994_2159# 0
C1716 a_4839_12857# a_4721_13809# 0
C1717 a_2343_5417# a_2706_5417# 0.00847f
C1718 a_10975_23147# sky130_fd_sc_hd__dfxbp_1_0.Q_N 0
C1719 a_3990_1761# a_3199_1791# 0.11873f
C1720 a_10953_14739# a_8193_13753# 0.09734f
C1721 a_4905_12113# a_4515_11543# 0
C1722 a_12993_23237# sky130_fd_sc_hd__dfxbp_1_3.Q_N 0
C1723 a_18553_4938# VDPWR 0
C1724 a_9451_16343# VDPWR 0.0252f
C1725 a_17264_22987# sky130_fd_sc_hd__dfxbp_1_3.Q_N 0
C1726 a_5363_5043# a_4840_5043# 0
C1727 a_9779_13785# a_10887_13773# 0.00104f
C1728 a_10717_13773# a_9779_13785# 0.00386f
C1729 a_4721_13809# a_4635_13809# 0.00658f
C1730 a_5080_2153# VDPWR 0
C1731 a_3010_2157# VDPWR 0
C1732 a_7221_1787# a_6698_1787# 0
C1733 a_11195_12931# a_11728_13649# 0.10646f
C1734 a_18667_24771# a_18667_25299# 0.04808f
C1735 a_3199_1791# a_4383_1787# 0.08312f
C1736 a_20384_16179# a_18742_16187# 0
C1737 a_10953_14739# a_11671_15239# 0.00366f
C1738 a_17521_23241# VDPWR 0.19863f
C1739 a_10953_14739# a_9779_13785# 0
C1740 a_6165_5409# a_6036_5017# 0.00792f
C1741 a_6335_1787# a_6071_1787# 0
C1742 a_10499_4853# a_10525_5837# 0
C1743 a_2343_5417# a_2217_5025# 0.0517f
C1744 a_8687_22875# a_8729_23143# 0
C1745 a_4847_14525# a_4513_14775# 0.1679f
C1746 a_23133_17137# a_21491_17145# 0
C1747 a_9579_12145# VDPWR 0.00297f
C1748 a_20877_17147# a_21491_17145# 0.10446f
C1749 a_10652_1793# a_9223_1793# 0.08907f
C1750 a_2313_1791# a_2259_2047# 0.00386f
C1751 a_14657_4547# VDPWR 0
C1752 a_4119_2153# VDPWR 0
C1753 a_4905_12113# a_4837_16089# 0
C1754 sky130_fd_sc_hd__dfxbp_1_7.Q_N a_18671_29203# 0.0031f
C1755 a_4839_12857# a_4849_11293# 0.82006f
C1756 a_4839_12857# a_5851_13769# 0.13054f
C1757 a_9781_10553# a_9715_11297# 0.00634f
C1758 a_7944_1767# a_8337_1793# 0.02283f
C1759 a_19063_29283# a_18671_29438# 0.00553f
C1760 a_16146_5447# VDPWR 0.35339f
C1761 a_13186_4919# a_12769_4809# 0.06611f
C1762 a_6087_14735# a_4513_14775# 0
C1763 a_18663_27120# a_18663_27252# 0.23675f
C1764 a_6389_13769# a_7749_14003# 0.00184f
C1765 sky130_fd_sc_hd__dfxbp_1_0.Q_N VDPWR 0.60587f
C1766 a_16660_2159# a_16243_2049# 0.06611f
C1767 a_10235_2049# a_6208_2817# 0.00304f
C1768 a_6208_2817# a_8700_1793# 0
C1769 a_23511_14701# a_23133_17137# 0.08871f
C1770 a_1950_5025# a_2079_5417# 0.00792f
C1771 sky130_fd_sc_hd__dfxbp_1_0.Q_N a_9160_23197# 0.12801f
C1772 a_23133_17137# sky130_fd_sc_hd__dfxbp_1_0.CLK 0.00444f
C1773 a_4849_11293# a_4515_11543# 0.16782f
C1774 a_10652_1793# a_10289_1793# 0.00985f
C1775 a_20877_17147# sky130_fd_sc_hd__dfxbp_1_0.CLK 0.0164f
C1776 a_19063_29283# sky130_fd_sc_hd__dfxbp_1_6.Q_N 0.00188f
C1777 a_9501_13813# a_4915_10549# 0.00128f
C1778 a_5851_13769# a_4635_13809# 0
C1779 a_4849_11293# a_4635_13809# 0.00317f
C1780 a_9369_16343# a_9629_14779# 0
C1781 a_4084_5017# a_4309_5409# 0.00559f
C1782 a_7749_14003# a_7831_14003# 0.00695f
C1783 a_14771_4803# a_13473_5459# 0
C1784 a_15188_4547# a_14771_4803# 0.03016f
C1785 a_9371_13111# VDPWR 0.54084f
C1786 a_18371_4938# a_17733_4529# 0.15188f
C1787 a_18689_27461# a_18663_27120# 0
C1788 a_18671_29438# a_18697_29233# 0.00772f
C1789 a_4625_15373# a_4635_13809# 0
C1790 a_18663_27017# sky130_fd_sc_hd__dfxbp_1_7.CLK 0.25091f
C1791 VDPWR a_19059_34232# 0
C1792 a_6021_13769# a_4903_15345# 0.00818f
C1793 a_6281_2043# a_6167_2153# 0
C1794 a_10109_22879# a_10891_23245# 0
C1795 uio_in[6] uio_in[7] 0.03102f
C1796 a_14179_2049# a_14233_2159# 0.03622f
C1797 a_6805_15235# a_7173_15235# 0
C1798 sky130_fd_sc_hd__inv_2_0.A a_19059_33811# 0
C1799 a_6208_2817# a_11836_1793# 0.00121f
C1800 a_4837_16089# a_5851_13769# 0.08387f
C1801 a_12295_22871# a_10975_23147# 0
C1802 a_4849_11293# a_4837_16089# 0.03118f
C1803 a_8038_5023# a_8263_5049# 0.00487f
C1804 a_14380_4547# a_6208_2817# 0
C1805 a_12295_22871# a_12736_22983# 0.11299f
C1806 a_19059_25272# a_18667_25299# 0
C1807 a_15242_5833# a_15431_5467# 0
C1808 a_14545_5467# a_13709_4553# 0
C1809 a_10525_5837# a_10132_5445# 0.02301f
C1810 a_19059_33811# a_18667_33966# 0.00553f
C1811 sky130_fd_sc_hd__dfxbp_1_9.Q a_19059_34232# 0
C1812 sky130_fd_sc_hd__dfxbp_1_5.CLK sky130_fd_sc_hd__dfxbp_1_4.Q_N 0.14813f
C1813 a_4837_16089# a_4625_15373# 0
C1814 a_11411_5471# a_12587_5825# 0.04534f
C1815 a_18693_31893# a_18667_31354# 0
C1816 a_21491_17145# sky130_fd_sc_hd__dfxbp_1_0.CLK 0.02037f
C1817 sky130_fd_sc_hd__dfxbp_1_2.CLK a_12129_22871# 0.25135f
C1818 a_9705_12861# a_9713_14529# 0.20053f
C1819 a_10108_4597# a_10132_5445# 0
C1820 a_18671_29731# a_18693_31299# 0
C1821 sky130_fd_sc_hd__dfxbp_1_7.Q_N a_18663_27120# 0.05782f
C1822 VDPWR a_4215_2153# 0
C1823 a_11195_12931# a_9779_13785# 0.0204f
C1824 a_7315_5043# a_8263_5049# 0
C1825 uio_oe[4] uio_oe[3] 0.03102f
C1826 a_9631_11547# VDPWR 0.33144f
C1827 a_11175_1793# a_12644_1793# 0.08907f
C1828 a_6208_2817# a_12430_4527# 0
C1829 a_9705_12861# a_10869_11939# 0
C1830 a_10289_2159# VDPWR 0.00967f
C1831 a_6208_2817# a_12559_4553# 0
C1832 a_17264_22987# a_17647_22875# 0
C1833 a_14233_1793# VDPWR 0.18611f
C1834 a_4477_5043# a_3229_5051# 0.08312f
C1835 a_12295_22871# a_12483_22871# 0.0967f
C1836 a_18667_33731# a_18693_33761# 0.0027f
C1837 a_11250_4963# a_11439_4597# 0
C1838 a_17096_23241# a_16657_22875# 0.27314f
C1839 a_18553_4938# a_9317_5049# 0.00526f
C1840 a_18671_29438# a_18671_29108# 0.07715f
C1841 a_6375_5299# a_6429_5043# 0.00386f
C1842 a_12295_22871# VDPWR 0.31439f
C1843 a_9577_15377# a_9491_15377# 0.00658f
C1844 a_11411_5471# a_12587_5459# 0.08312f
C1845 a_18667_31449# a_18671_30311# 0
C1846 a_13520_4919# a_12769_4809# 0.00696f
C1847 a_4847_14525# VDPWR 0.482f
C1848 a_14771_4803# a_14491_5723# 0
C1849 a_13969_2159# a_13788_1793# 0
C1850 VDPWR a_6167_2153# 0
C1851 a_16454_4503# a_16146_5447# 0
C1852 a_14179_2049# a_15852_1793# 0
C1853 sky130_fd_sc_hd__dfxbp_1_6.Q_N a_18671_29108# 0.51145f
C1854 a_9503_10581# a_9715_11297# 0
C1855 a_4847_14525# a_4763_14775# 0.07979f
C1856 a_6087_14735# VDPWR 0.62614f
C1857 a_5174_5409# a_2217_5025# 0
C1858 a_12323_5459# VDPWR 0.00118f
C1859 a_10841_12931# a_11728_13649# 0
C1860 a_2289_5307# a_3040_5051# 0.00682f
C1861 sky130_fd_sc_hd__dfxbp_1_9.Q_N a_18667_33731# 0.00244f
C1862 a_6208_2817# a_10652_2159# 0
C1863 a_15904_1767# a_16033_1793# 0.00758f
C1864 a_23761_14335# ui_in[0] 0.05164f
C1865 a_9317_5049# a_16146_5447# 0
C1866 a_6208_2817# ui_in[1] 0.16407f
C1867 sky130_fd_sc_hd__dfxbp_1_5.Q_N a_18693_25215# 0
C1868 a_4637_10577# VDPWR 0.43224f
C1869 a_6635_15235# a_4837_16089# 0.232f
C1870 a_14908_5467# a_14545_5467# 0.00985f
C1871 a_6208_2817# a_14233_2159# 0
C1872 a_15188_4547# a_6208_2817# 0
C1873 a_9703_16093# a_11728_13649# 0
C1874 a_4840_5409# a_4477_5409# 0.00847f
C1875 a_18693_31299# sky130_fd_sc_hd__dfxbp_1_9.Q_N 0.142f
C1876 a_4329_2043# a_2187_1765# 0.00305f
C1877 VDPWR a_8169_2159# 0
C1878 a_9556_17271# a_8193_13753# 0.15228f
C1879 a_16902_5839# a_16485_5729# 0.06611f
C1880 a_4915_10549# a_9771_12117# 0.00452f
C1881 a_7126_5043# VDPWR 0
C1882 a_18671_29438# sky130_fd_sc_hd__dfxbp_1_9.CLK 0
C1883 a_6792_5043# a_6238_6077# 0
C1884 a_4849_11293# a_4905_12113# 0.25133f
C1885 a_5269_1787# a_6698_1787# 0.08907f
C1886 a_5363_5043# a_7315_5043# 0
C1887 a_24234_14385# a_24962_14701# 0.1456f
C1888 a_17521_23241# sky130_fd_sc_hd__dfxbp_1_5.CLK 0.00402f
C1889 a_10499_4853# a_11250_4963# 0.00696f
C1890 a_2187_1765# a_4746_2153# 0
C1891 a_17689_23143# a_16823_22875# 0.03136f
C1892 a_4913_13781# a_5933_13769# 0
C1893 sky130_fd_sc_hd__dfxbp_1_5.Q_N a_18693_24621# 0.142f
C1894 a_6629_15387# a_4903_15345# 0
C1895 a_11411_5471# a_11439_4597# 0
C1896 a_3990_1761# VDPWR 0.34976f
C1897 a_18667_33636# a_18667_34259# 0.03136f
C1898 a_10675_14767# a_10841_12931# 0
C1899 a_18663_27545# a_18663_28125# 0.10805f
C1900 a_18667_31552# sky130_fd_sc_hd__dfxbp_1_6.Q_N 0
C1901 a_7749_14003# a_7927_14003# 0.00412f
C1902 a_11777_15239# VDPWR 0
C1903 sky130_fd_sc_hd__dfxbp_1_9.CLK sky130_fd_sc_hd__dfxbp_1_6.Q_N 0.15244f
C1904 a_12587_5459# a_12419_5459# 0
C1905 a_6429_5043# a_6036_5017# 0.02283f
C1906 a_12865_14007# a_11147_11911# 0
C1907 a_4840_5409# a_2217_5025# 0
C1908 a_10160_4571# a_8431_5049# 0
C1909 a_10357_5471# a_10132_5445# 0.00487f
C1910 a_9579_12145# a_9715_11297# 0
C1911 a_2187_1765# a_5890_1787# 0.00121f
C1912 a_14065_2159# VDPWR 0
C1913 a_9713_14529# a_9769_15349# 0.15229f
C1914 VDPWR a_4383_1787# 0.1861f
C1915 a_9781_10553# a_10717_13773# 0.00192f
C1916 a_9713_14529# VDPWR 0.48168f
C1917 a_9556_17271# a_18742_16187# 0
C1918 a_23511_14335# VDPWR 0.00538f
C1919 a_6071_2153# a_5890_1787# 0
C1920 a_4423_5299# a_4309_5043# 0
C1921 sky130_fd_sc_hd__dfxbp_1_1.Q_N a_11406_23201# 0.12801f
C1922 a_12655_4553# a_12769_4809# 0
C1923 sky130_fd_sc_hd__dfxbp_1_3.CLK a_12694_22871# 0
C1924 a_9703_16093# a_10675_14767# 0.03093f
C1925 a_18553_4938# a_6238_6077# 0
C1926 a_4309_5043# VDPWR 0
C1927 a_4763_14525# a_4513_14775# 0.00723f
C1928 a_9379_14779# a_9703_16093# 0
C1929 a_7944_1767# a_8073_1793# 0.00758f
C1930 a_18663_27017# a_18667_25879# 0
C1931 a_13161_23139# a_12736_22983# 0
C1932 a_10869_11939# VDPWR 0.22392f
C1933 a_19055_27097# sky130_fd_sc_hd__dfxbp_1_7.CLK 0
C1934 a_1920_1765# a_2049_1791# 0.00758f
C1935 a_16657_22875# VDPWR 0.66128f
C1936 a_18667_24676# a_18667_24771# 0.96835f
C1937 a_6208_2817# a_8337_1793# 0
C1938 a_6208_2817# a_15852_1793# 0.00174f
C1939 a_4849_11293# a_5851_13769# 0.17512f
C1940 a_9703_16093# a_10799_13773# 0
C1941 a_12615_14007# a_12039_15239# 0.16707f
C1942 a_7749_14003# a_7999_14003# 0.00876f
C1943 sky130_fd_sc_hd__dfxbp_1_7.Q a_19055_27518# 0
C1944 a_9556_17271# a_17254_16187# 0
C1945 a_6208_2817# a_9844_1793# 0.00121f
C1946 VDPWR a_18113_17153# 0.45396f
C1947 a_10235_2049# a_10121_1793# 0
C1948 sky130_fd_sc_hd__dfxbp_1_7.Q_N a_18671_29108# 0.00115f
C1949 a_16297_2159# a_16129_2159# 0
C1950 a_8193_13753# a_9703_16093# 0.36685f
C1951 a_10109_22879# a_10297_22879# 0.0967f
C1952 a_9779_13785# a_10841_12931# 0.08477f
C1953 a_16033_2159# a_15852_1793# 0
C1954 a_4723_10577# VDPWR 0.00176f
C1955 a_9371_13111# a_9715_11297# 0.00372f
C1956 a_9781_10553# a_12793_14007# 0
C1957 a_21506_16181# a_19510_16177# 0
C1958 a_4329_2043# a_4215_1787# 0
C1959 a_4755_13107# a_4839_12857# 0.08134f
C1960 a_6281_11907# a_4915_10549# 0.43338f
C1961 a_6238_6077# a_16146_5447# 0.00525f
C1962 a_23731_14309# a_23511_14335# 0.0457f
C1963 a_12017_1793# a_11888_1767# 0.00758f
C1964 a_11411_5471# a_10499_4853# 0
C1965 a_17011_22875# a_16823_22875# 0.0967f
C1966 uio_oe[0] uio_oe[1] 0.03102f
C1967 a_14377_5467# a_14545_5467# 0
C1968 a_15242_5833# VDPWR 0
C1969 a_11671_15239# a_9703_16093# 0
C1970 a_11175_1793# a_12281_2159# 0.04534f
C1971 a_13161_23139# VDPWR 0.5127f
C1972 a_10986_1793# a_6208_2817# 0
C1973 a_9779_13785# a_9703_16093# 0.01745f
C1974 a_14233_1793# a_14065_1793# 0
C1975 a_8167_5415# VDPWR 0
C1976 a_18693_34175# a_18667_34470# 0.00851f
C1977 a_4755_13107# a_4635_13809# 0
C1978 a_8561_23241# sky130_fd_sc_hd__dfxbp_1_0.CLK 0
C1979 a_23761_14335# a_23133_17137# 0.06603f
C1980 a_2259_2047# a_3199_1791# 0.13962f
C1981 a_18663_27545# VDPWR 0.51574f
C1982 a_14541_22875# sky130_fd_sc_hd__dfxbp_1_3.Q_N 0.5114f
C1983 a_12039_15239# a_11979_13399# 0.41061f
C1984 a_7315_5043# a_8794_5049# 0.08907f
C1985 a_8073_2159# a_7892_1793# 0
C1986 a_4847_14525# a_6805_15235# 0.00624f
C1987 a_7113_13395# a_4903_15345# 0
C1988 a_4839_12857# a_6129_12927# 0.00312f
C1989 a_6208_2817# a_16129_2159# 0
C1990 a_20109_17157# VDPWR 0.44007f
C1991 a_12615_14007# a_11979_13399# 0.27996f
C1992 a_10525_5471# a_10261_5471# 0
C1993 a_9631_11547# a_9715_11297# 0.08177f
C1994 a_1898_5051# a_2079_5417# 0
C1995 a_2289_5307# a_2175_5417# 0
C1996 a_10382_23245# a_10477_23245# 0.00772f
C1997 a_15711_4547# a_16679_4529# 0
C1998 sky130_fd_sc_hd__dfxbp_1_5.Q_N a_18663_27756# 0
C1999 sky130_fd_sc_hd__dfxbp_1_4.CLK a_16823_22875# 0.01409f
C2000 a_12281_2159# a_12644_2159# 0.00847f
C2001 a_6087_14735# a_6805_15235# 0.00366f
C2002 a_7221_1787# a_7944_1767# 0.11881f
C2003 a_2049_2157# VDPWR 0
C2004 a_18667_34259# a_18667_33834# 0
C2005 sky130_fd_sc_hd__dfxbp_1_0.Q_N a_8645_23241# 0
C2006 a_4329_2043# a_5942_1761# 0.00419f
C2007 ui_in[0] a_24152_14385# 0.03419f
C2008 a_6208_2817# a_10385_4597# 0
C2009 a_2217_5025# a_6036_5017# 0
C2010 a_8136_23241# a_8051_22875# 0.03733f
C2011 a_9896_1767# a_10025_2159# 0.00792f
C2012 a_9463_11547# VDPWR 0.02521f
C2013 a_18667_33636# a_18667_34470# 0.19462f
C2014 a_4765_11543# a_4515_11543# 0.02504f
C2015 a_17689_23143# sky130_fd_sc_hd__dfxbp_1_4.CLK 0
C2016 a_17210_4529# VDPWR 0.21928f
C2017 sky130_fd_sc_hd__dfxbp_1_1.Q_N a_10933_22879# 0.00125f
C2018 a_16902_5473# a_15711_4547# 0
C2019 a_12295_22871# sky130_fd_sc_hd__dfxbp_1_2.Q_N 0.5114f
C2020 a_7986_5049# VDPWR 0.16479f
C2021 a_8073_2159# a_8337_2159# 0
C2022 a_18667_33966# a_18693_33761# 0.00772f
C2023 a_4763_14525# VDPWR 0.00474f
C2024 a_23511_14335# a_23677_14335# 0.00648f
C2025 a_8193_13753# a_7999_14003# 0
C2026 sky130_fd_sc_hd__inv_8_0.A VDPWR 1.19708f
C2027 a_18663_27017# a_18663_28125# 0
C2028 a_12559_4919# a_12378_4553# 0
C2029 sky130_fd_sc_hd__dfxbp_1_1.Q_N a_10975_23147# 0.12218f
C2030 sky130_fd_sc_hd__dfxbp_1_1.Q_N a_12736_22983# 0
C2031 a_14561_4547# a_6208_2817# 0
C2032 a_17345_17163# sky130_fd_sc_hd__dfxbp_1_0.CLK 0.02041f
C2033 a_5942_1761# a_5890_1787# 0.1439f
C2034 a_23761_14335# a_23511_14701# 0.05408f
C2035 a_17264_22987# a_17605_23241# 0
C2036 sky130_fd_sc_hd__dfxbp_1_2.CLK a_11406_23201# 0.2081f
C2037 a_4903_15345# a_6862_13645# 0
C2038 a_8262_22875# a_8304_22987# 0
C2039 a_23761_14335# sky130_fd_sc_hd__dfxbp_1_0.CLK 0.00101f
C2040 VDPWR a_18697_29053# 0.07699f
C2041 a_24234_14385# a_24774_14701# 0.17579f
C2042 a_7944_1767# a_7892_1793# 0.1439f
C2043 a_18667_31449# a_18693_31479# 0.0027f
C2044 a_9769_15349# a_9491_15377# 0.12165f
C2045 a_2187_1765# a_5269_1787# 0.00136f
C2046 a_9491_15377# VDPWR 0.4511f
C2047 a_12655_4919# VDPWR 0
C2048 sky130_fd_sc_hd__dfxbp_1_9.Q_N a_18667_33966# 0
C2049 a_11501_15239# a_9769_15349# 0
C2050 a_18667_33636# a_18667_31449# 0
C2051 a_4839_12857# a_4627_12141# 0
C2052 a_11501_15239# VDPWR 0.42363f
C2053 a_6238_6077# a_12323_5459# 0
C2054 a_18667_25006# a_18667_24676# 0.07715f
C2055 a_4423_5299# a_4084_5017# 0.04737f
C2056 a_24318_14385# a_24774_14701# 0.01242f
C2057 a_9223_1793# a_8283_2049# 0.13739f
C2058 a_4084_5017# VDPWR 0.34979f
C2059 a_6208_2817# a_12769_4809# 0
C2060 sky130_fd_sc_hd__dfxbp_1_1.Q_N a_12483_22871# 0
C2061 a_10160_4571# a_10108_4597# 0.1439f
C2062 a_15641_17149# a_17254_16187# 0
C2063 a_6389_13769# a_6944_13645# 0.00183f
C2064 a_2217_5025# a_3040_5417# 0
C2065 a_4627_12141# a_4515_11543# 0
C2066 sky130_fd_sc_hd__dfxbp_1_4.CLK a_17011_22875# 0
C2067 sky130_fd_sc_hd__dfxbp_1_1.Q_N VDPWR 0.60723f
C2068 a_10499_4853# a_10160_4571# 0.04737f
C2069 sky130_fd_sc_hd__inv_4_0.A VDPWR 0.63754f
C2070 a_16371_5473# a_15431_5467# 0
C2071 a_14729_22875# sky130_fd_sc_hd__dfxbp_1_3.Q_N 0.142f
C2072 a_18663_27545# a_18671_29203# 0
C2073 a_4627_12141# a_4635_13809# 0
C2074 a_11175_1793# a_12644_2159# 0.03325f
C2075 a_12142_5459# VDPWR 0.16775f
C2076 a_7944_1767# a_8337_2159# 0.02301f
C2077 sky130_fd_sc_hd__dfxbp_1_1.Q_N a_9160_23197# 0
C2078 a_6238_6077# a_7126_5043# 0
C2079 a_9713_14529# a_9715_11297# 0.00506f
C2080 a_13186_4553# a_6208_2817# 0
C2081 a_18667_34259# VDPWR 0.51525f
C2082 sky130_fd_sc_hd__dfxbp_1_5.CLK a_16657_22875# 0.0016f
C2083 VDPWR sky130_fd_sc_hd__inv_6_0.A 0.97191f
C2084 a_23677_14701# ui_in[0] 0.02125f
C2085 a_14375_22875# a_16823_22875# 0
C2086 a_9781_10553# a_9556_17271# 0.15958f
C2087 a_15711_4547# a_16847_4529# 0.08312f
C2088 a_10553_4597# a_10385_4597# 0
C2089 a_4839_12857# a_6281_11907# 0.02321f
C2090 a_17733_4529# a_6208_2817# 0
C2091 a_18693_24801# VDPWR 0.00347f
C2092 a_9705_12861# a_4915_10549# 0
C2093 a_10869_11939# a_9715_11297# 0.10273f
C2094 a_18667_24874# sky130_fd_sc_hd__dfxbp_1_7.CLK 0
C2095 a_1868_1791# a_2049_2157# 0
C2096 a_18689_27461# a_18663_27756# 0.00851f
C2097 a_9556_17271# a_18128_16189# 0
C2098 a_18113_17153# a_19235_17155# 0.101f
C2099 a_4839_12857# a_4587_13107# 0
C2100 a_11147_11911# a_10955_11939# 0
C2101 a_18671_29731# a_18667_31354# 0
C2102 sky130_fd_sc_hd__dfxbp_1_5.Q_N a_19059_24851# 0.00188f
C2103 a_6629_15387# a_8193_13753# 0.05689f
C2104 a_9223_1793# a_10289_1793# 0.08312f
C2105 a_6208_2817# a_8073_1793# 0
C2106 a_18667_33834# a_18667_34470# 0.03684f
C2107 a_10235_2049# a_10289_2159# 0.03622f
C2108 a_18663_27017# VDPWR 0.66226f
C2109 a_15239_23241# sky130_fd_sc_hd__dfxbp_1_3.Q_N 0.09273f
C2110 a_7113_13395# a_7749_14003# 0.27996f
C2111 sky130_fd_sc_hd__dfxbp_1_9.Q a_18667_34259# 0
C2112 a_9943_22879# sky130_fd_sc_hd__dfxbp_1_0.Q_N 0.00248f
C2113 a_6238_6077# a_23511_14335# 0.00544f
C2114 a_24241_14651# a_24774_14701# 0.0098f
C2115 a_6389_13769# a_7173_15235# 0.00147f
C2116 uio_out[5] uio_out[4] 0.03102f
C2117 a_4905_12113# a_6129_12927# 0
C2118 a_10955_11939# a_9771_12117# 0
C2119 a_4503_16339# a_4513_14775# 0.00102f
C2120 a_18839_4938# a_18625_4938# 0.00557f
C2121 a_18693_31479# a_18667_31684# 0.00772f
C2122 sky130_fd_sc_hd__dfxbp_1_7.Q a_18671_29731# 0
C2123 a_6003_11935# a_4915_10549# 0
C2124 a_9587_13813# a_4915_10549# 0
C2125 a_12227_2049# a_13788_1793# 0
C2126 a_16297_2159# a_16243_2049# 0.03622f
C2127 a_13119_22871# sky130_fd_sc_hd__dfxbp_1_3.CLK 0
C2128 sky130_fd_sc_hd__dfxbp_1_2.CLK a_10933_22879# 0
C2129 a_18663_27756# sky130_fd_sc_hd__dfxbp_1_7.Q_N 0.09273f
C2130 a_10357_5837# VDPWR 0
C2131 a_7697_22875# sky130_fd_sc_hd__dfxbp_1_0.CLK 0.24853f
C2132 a_4755_13107# a_4849_11293# 0
C2133 a_13840_1767# a_13969_1793# 0.00758f
C2134 a_16371_5839# a_16539_5839# 0
C2135 a_17210_4529# a_16793_4785# 0.03016f
C2136 sky130_fd_sc_hd__dfxbp_1_8.Q_N a_19059_34232# 0.00125f
C2137 sky130_fd_sc_hd__dfxbp_1_2.Q_N a_13161_23139# 0.12218f
C2138 a_10160_4571# a_10132_5445# 0
C2139 a_8283_2049# a_8169_1793# 0
C2140 a_8377_5305# a_8431_5049# 0.00386f
C2141 a_4903_15345# a_4913_13781# 0.11601f
C2142 a_15119_1793# a_15852_1793# 0.0495f
C2143 a_16033_1793# a_16297_1793# 0
C2144 a_20109_17157# a_19235_17155# 0.1036f
C2145 a_18663_27545# a_18663_27120# 0
C2146 a_18697_29053# a_18671_29203# 0.06222f
C2147 a_2343_5417# VDPWR 0.00939f
C2148 a_9556_17271# a_16486_16197# 0
C2149 a_4765_11293# VDPWR 0.00377f
C2150 a_18667_32188# VDPWR 0.1998f
C2151 sky130_fd_sc_hd__dfxbp_1_2.CLK a_10975_23147# 0.1234f
C2152 sky130_fd_sc_hd__dfxbp_1_2.CLK a_12736_22983# 0
C2153 a_24407_14651# VDPWR 0.00288f
C2154 a_13167_1793# VDPWR 1.38964f
C2155 a_9781_10553# a_9703_16093# 0.01618f
C2156 a_2259_2047# VDPWR 0.44946f
C2157 a_8193_13753# a_9619_16343# 0
C2158 a_9781_10553# a_12697_14007# 0
C2159 a_18667_25510# a_18667_24771# 0.03218f
C2160 a_18742_16187# a_19510_16177# 0.1036f
C2161 a_6238_6077# a_15242_5833# 0
C2162 a_12194_5433# a_10471_5727# 0.00291f
C2163 a_18667_24676# a_18667_25299# 0.03136f
C2164 sky130_fd_sc_hd__dfxbp_1_9.Q_N a_18667_31354# 0.51145f
C2165 a_6208_2817# a_7032_2153# 0
C2166 a_6208_2817# a_16243_2049# 0.15654f
C2167 a_4849_11293# a_6129_12927# 0
C2168 a_18689_26867# a_18663_26922# 0.0967f
C2169 a_12993_23237# sky130_fd_sc_hd__dfxbp_1_3.CLK 0.0039f
C2170 a_9705_12861# a_9461_14779# 0
C2171 a_8167_5415# a_6238_6077# 0
C2172 a_5942_1761# a_5269_1787# 0.11878f
C2173 a_2676_2157# a_2187_1765# 0.03547f
C2174 sky130_fd_sc_hd__dfxbp_1_9.Q a_18667_32188# 0.00387f
C2175 a_9463_11547# a_9715_11297# 0
C2176 a_9779_13785# a_10995_12931# 0
C2177 a_16539_5473# a_16371_5473# 0
C2178 a_4849_11293# a_4765_11543# 0.08177f
C2179 a_7221_1787# a_6208_2817# 0.00288f
C2180 a_14432_4521# a_14561_4913# 0.00792f
C2181 a_12281_1793# a_12017_1793# 0
C2182 a_10499_4853# a_10525_5471# 0
C2183 a_2313_2157# VDPWR 0.00827f
C2184 sky130_fd_sc_hd__dfxbp_1_2.CLK a_12483_22871# 0
C2185 a_12017_1793# VDPWR 0.00116f
C2186 a_22365_17147# a_22274_16171# 0.02069f
C2187 a_17254_16187# a_19510_16177# 0
C2188 a_12823_4553# a_11439_4597# 0.08312f
C2189 uio_out[2] uio_out[3] 0.03102f
C2190 a_18693_31299# sky130_fd_sc_hd__dfxbp_1_6.Q_N 0
C2191 a_12039_15239# a_11147_11911# 0.09952f
C2192 sky130_fd_sc_hd__dfxbp_1_1.CLK a_10109_22879# 0.01405f
C2193 a_7113_13395# a_8193_13753# 0.03478f
C2194 sky130_fd_sc_hd__dfxbp_1_5.Q_N a_18663_26922# 0.0011f
C2195 a_12823_4919# a_12655_4919# 0
C2196 sky130_fd_sc_hd__dfxbp_1_2.CLK VDPWR 0.27173f
C2197 VDPWR a_18667_34470# 0.1998f
C2198 a_4905_12113# a_4627_12141# 0.12057f
C2199 a_15904_1767# VDPWR 0.34924f
C2200 a_18667_32188# a_18667_31977# 0.31062f
C2201 a_23677_14701# a_23133_17137# 0.00696f
C2202 sky130_fd_sc_hd__dfxbp_1_4.Q_N a_15838_23197# 0
C2203 a_12295_22871# a_9943_22879# 0
C2204 a_12615_14007# a_11147_11911# 0.19234f
C2205 a_10807_23245# a_10891_23245# 0.00851f
C2206 a_6261_5043# VDPWR 0
C2207 VDPWR a_4915_10549# 0.84484f
C2208 a_14375_22875# sky130_fd_sc_hd__dfxbp_1_4.CLK 0
C2209 a_9621_13111# a_9493_12145# 0
C2210 a_9371_13111# a_11195_12931# 0
C2211 a_14982_22987# sky130_fd_sc_hd__dfxbp_1_3.Q_N 0.05782f
C2212 a_18663_27017# a_18671_29203# 0
C2213 a_7986_5049# a_6238_6077# 0.00121f
C2214 a_10652_2159# a_10289_2159# 0.00847f
C2215 a_13840_1767# a_13969_2159# 0.00792f
C2216 sky130_fd_sc_hd__dfxbp_1_9.Q a_18667_34470# 0
C2217 a_8304_22987# sky130_fd_sc_hd__dfxbp_1_0.CLK 0
C2218 a_18667_31449# a_18671_29942# 0
C2219 a_19059_31529# VDPWR 0
C2220 a_5975_12927# a_4839_12857# 0.29952f
C2221 a_16146_5447# a_14491_5723# 0.00354f
C2222 a_10160_4571# a_10289_4597# 0.00758f
C2223 a_9379_14779# a_9629_14779# 0.02504f
C2224 a_14375_22875# a_12568_23237# 0
C2225 a_11411_5471# a_12419_5459# 0
C2226 a_4503_16339# VDPWR 0.54671f
C2227 a_2259_2047# a_3010_1791# 0.00682f
C2228 a_6281_2043# a_6167_1787# 0
C2229 a_6429_5409# a_6375_5299# 0.03622f
C2230 a_4213_5409# a_4084_5017# 0.00792f
C2231 a_4905_12113# a_6281_11907# 0.03573f
C2232 a_10109_22879# a_10807_23245# 0.19462f
C2233 a_18667_25510# a_19059_25272# 0.00617f
C2234 a_6208_2817# a_7892_1793# 0.00121f
C2235 a_15711_4547# a_16539_5839# 0
C2236 sky130_fd_sc_hd__inv_8_0.A sky130_fd_sc_hd__inv_16_0.A 0
C2237 a_16371_5473# VDPWR 0
C2238 a_6208_2817# a_13788_1793# 0.00121f
C2239 a_4505_13107# a_6329_12927# 0
C2240 a_11147_11911# a_11979_13399# 0.19569f
C2241 sky130_fd_sc_hd__dfxbp_1_3.CLK sky130_fd_sc_hd__dfxbp_1_3.Q_N 0.0174f
C2242 a_4763_14775# a_4503_16339# 0
C2243 a_14729_22875# a_14909_23241# 0.00123f
C2244 a_2187_1765# a_3938_1787# 0.00121f
C2245 a_4839_12857# a_4513_14775# 0.00442f
C2246 a_2259_2047# a_2145_2157# 0
C2247 a_15407_23143# a_16823_22875# 0
C2248 a_12865_14007# VDPWR 0
C2249 a_10261_5471# VDPWR 0.00116f
C2250 a_4849_11293# a_4627_12141# 0.0022f
C2251 sky130_fd_sc_hd__dfxbp_1_9.Q a_19059_31529# 0
C2252 a_10953_14739# a_11777_15239# 0.00651f
C2253 a_18667_31449# VDPWR 0.6622f
C2254 a_10717_13773# a_9713_14529# 0
C2255 a_12823_4553# a_10499_4853# 0
C2256 sky130_fd_sc_hd__dfxbp_1_1.Q_N sky130_fd_sc_hd__dfxbp_1_2.Q_N 0
C2257 a_4213_5043# a_2217_5025# 0
C2258 sky130_fd_sc_hd__dfxbp_1_0.Q_N a_8729_23143# 0.12218f
C2259 a_10132_5445# a_10525_5471# 0.02283f
C2260 a_6238_6077# a_12655_4919# 0
C2261 a_12129_22871# a_12568_23237# 0.27314f
C2262 a_19055_27097# VDPWR 0
C2263 a_12227_2049# a_12644_1793# 0.03016f
C2264 a_11411_5471# a_11222_5837# 0
C2265 a_14100_5467# a_14281_5833# 0
C2266 a_13592_23193# a_14375_22875# 0
C2267 a_23677_14701# a_23511_14701# 0.05551f
C2268 a_10953_14739# a_9713_14529# 0.3079f
C2269 clk ena 0.03102f
C2270 a_16094_5473# a_15431_5467# 0.05029f
C2271 a_15522_4913# VDPWR 0
C2272 a_4635_13809# a_4513_14775# 0.00144f
C2273 a_4903_15345# a_5933_13769# 0.0035f
C2274 a_6208_2817# a_8337_2159# 0
C2275 a_4423_5299# a_5174_5409# 0.00696f
C2276 a_10652_1793# VDPWR 0.21795f
C2277 a_8136_23241# sky130_fd_sc_hd__dfxbp_1_1.CLK 0
C2278 a_5174_5409# VDPWR 0
C2279 a_6003_11935# a_4839_12857# 0
C2280 a_14541_22875# a_14729_22875# 0.0967f
C2281 a_18667_31449# sky130_fd_sc_hd__dfxbp_1_9.Q 0
C2282 a_5975_12927# a_4837_16089# 0
C2283 a_2313_2157# a_2145_2157# 0
C2284 a_10357_5471# a_10525_5471# 0
C2285 a_16402_4529# a_15711_4547# 0.0498f
C2286 a_10080_5471# a_10261_5837# 0
C2287 a_9461_14779# a_9769_15349# 0
C2288 a_18663_27252# a_18663_26922# 0.07715f
C2289 a_16486_16197# a_15641_17149# 0.10145f
C2290 a_18663_27545# a_18671_29108# 0
C2291 a_8431_5049# VDPWR 0.18609f
C2292 a_9461_14779# VDPWR 0.02521f
C2293 a_18663_27017# a_18663_27120# 0.14145f
C2294 a_9589_10581# VDPWR 0.00176f
C2295 a_11888_1767# a_12017_2159# 0.00792f
C2296 a_24234_14385# a_6208_2817# 0.04349f
C2297 a_7697_22875# a_8561_23241# 0.03218f
C2298 a_1950_5025# a_2175_5417# 0.00559f
C2299 a_7173_15235# a_6717_15235# 0
C2300 a_6281_11907# a_5851_13769# 0
C2301 a_4849_11293# a_6281_11907# 0.00683f
C2302 a_2217_5025# a_2706_5417# 0.0357f
C2303 a_6238_6077# a_12142_5459# 0.003f
C2304 a_15711_4547# a_15431_5467# 0
C2305 a_10888_5837# a_10471_5727# 0.06611f
C2306 a_17544_4529# VDPWR 0
C2307 a_4477_5409# a_2217_5025# 0
C2308 a_13592_23193# a_12129_22871# 0
C2309 a_8038_5023# a_6792_5043# 0
C2310 a_18697_29053# a_18697_29233# 0.00123f
C2311 VDPWR a_6167_1787# 0
C2312 a_4849_11293# a_4587_13107# 0
C2313 a_4837_16089# a_4513_14775# 0
C2314 a_18667_31449# a_18667_31977# 0.04808f
C2315 a_3199_1791# a_4383_2153# 0.04534f
C2316 a_6208_2817# a_24318_14385# 0.05111f
C2317 a_12587_5825# VDPWR 0.01034f
C2318 a_7126_5409# VDPWR 0
C2319 a_9703_16093# a_9451_16343# 0
C2320 a_22365_17147# VDPWR 0.35781f
C2321 a_16129_1793# VDPWR 0
C2322 a_6429_5409# a_6036_5017# 0.02301f
C2323 a_6208_2817# a_16994_1793# 0
C2324 sky130_fd_sc_hd__dfxbp_1_1.CLK a_8051_22875# 0
C2325 a_13167_1793# a_14065_1793# 0
C2326 a_8377_5305# a_10108_4597# 0
C2327 a_8262_22875# VDPWR 0
C2328 a_16275_5473# a_15431_5467# 0
C2329 a_14432_4521# a_13709_4553# 0.11874f
C2330 a_10550_22991# a_10891_23245# 0
C2331 a_18689_27461# a_18663_26922# 0
C2332 a_14541_22875# a_15239_23241# 0.19462f
C2333 a_10508_22879# sky130_fd_sc_hd__dfxbp_1_1.CLK 0
C2334 a_7173_15235# a_7999_14003# 0
C2335 clk rst_n 0.03102f
C2336 a_23133_17137# a_22274_16171# 0.10226f
C2337 a_15188_4913# a_13709_4553# 0.03325f
C2338 a_6792_5043# a_7315_5043# 0
C2339 ui_in[0] VDPWR 0.77926f
C2340 a_15711_4547# a_17210_4895# 0.03325f
C2341 a_4847_14525# a_6389_13769# 0
C2342 a_4423_5299# a_4840_5409# 0.06611f
C2343 a_20109_17157# a_20384_16179# 0.00293f
C2344 a_14065_2159# a_14233_2159# 0
C2345 a_6003_11935# a_4837_16089# 0
C2346 a_4840_5409# VDPWR 0.02103f
C2347 sky130_fd_sc_hd__dfxbp_1_1.CLK a_10297_22879# 0
C2348 uio_out[6] uio_out[5] 0.03102f
C2349 a_8794_5415# a_6375_5299# 0
C2350 a_18667_31684# VDPWR 0.25534f
C2351 a_18625_5265# VDPWR 0
C2352 a_12587_5459# VDPWR 0.18754f
C2353 a_6389_13769# a_6087_14735# 0.00238f
C2354 a_16679_4529# a_16847_4529# 0
C2355 a_14375_22875# a_12129_22871# 0
C2356 a_18693_31893# sky130_fd_sc_hd__dfxbp_1_9.Q_N 0
C2357 a_17191_23241# a_16657_22875# 0.0027f
C2358 a_15711_4547# a_16583_4529# 0
C2359 a_9619_16093# VDPWR 0.00495f
C2360 a_10550_22991# a_10109_22879# 0.11299f
C2361 sky130_fd_sc_hd__dfxbp_1_7.Q_N a_18663_26922# 0.51145f
C2362 a_10357_5837# a_6238_6077# 0
C2363 a_7863_22875# sky130_fd_sc_hd__dfxbp_1_0.CLK 0.01356f
C2364 a_9371_13111# a_10841_12931# 0
C2365 a_5269_1787# a_6208_2817# 0.00234f
C2366 a_6429_5409# a_6165_5409# 0
C2367 a_18553_4938# a_17733_4529# 0.00143f
C2368 a_18697_29053# a_18671_29108# 0.0967f
C2369 a_6375_5299# VDPWR 0.45147f
C2370 a_18689_27047# VDPWR 0.00349f
C2371 a_23731_14309# ui_in[0] 0.45726f
C2372 sky130_fd_sc_hd__dfxbp_1_9.Q a_18667_31684# 0
C2373 a_4839_12857# VDPWR 1.04909f
C2374 a_16371_5839# VDPWR 0
C2375 sky130_fd_sc_hd__dfxbp_1_4.Q_N a_17222_22875# 0.00188f
C2376 a_6208_2817# a_24241_14651# 0.03575f
C2377 a_18667_31449# a_18671_29203# 0
C2378 a_18128_16189# a_19510_16177# 0
C2379 sky130_fd_sc_hd__dfxbp_1_5.Q_N a_18667_24771# 0.11931f
C2380 a_6238_6077# a_24407_14651# 0
C2381 a_3199_1791# a_4119_1787# 0
C2382 a_15407_23143# sky130_fd_sc_hd__dfxbp_1_4.CLK 0.12293f
C2383 a_6629_15387# a_5809_14763# 0
C2384 a_4839_12857# a_4763_14775# 0.00187f
C2385 VDPWR a_4515_11543# 0.53681f
C2386 a_8561_23241# a_8304_22987# 0.03684f
C2387 a_5975_12927# a_4905_12113# 0
C2388 a_6208_2817# a_12644_1793# 0
C2389 VDPWR a_4635_13809# 0.43903f
C2390 sky130_fd_sc_hd__dfxbp_1_2.CLK sky130_fd_sc_hd__dfxbp_1_2.Q_N 0.01749f
C2391 a_9715_11297# a_4915_10549# 0
C2392 a_15119_1793# a_16243_2049# 0.21187f
C2393 a_8377_5305# a_10132_5445# 0
C2394 a_9713_14529# a_11583_15239# 0.00159f
C2395 a_11439_4597# VDPWR 1.62298f
C2396 a_8431_5415# a_8167_5415# 0
C2397 a_4763_14775# a_4635_13809# 0
C2398 a_23761_14335# a_24152_14385# 0.02235f
C2399 a_16539_5473# a_15711_4547# 0
C2400 a_6629_15387# a_7173_15235# 0.00221f
C2401 ui_in[3] ui_in[2] 0.03102f
C2402 a_3199_1791# a_4746_1787# 0.08907f
C2403 sky130_fd_sc_hd__dfxbp_1_9.CLK a_18697_29053# 0
C2404 a_4837_16089# VDPWR 1.33864f
C2405 a_18667_25510# a_18667_25299# 0.31062f
C2406 a_9128_5049# a_8377_5305# 0.00682f
C2407 a_14908_5467# a_13709_4553# 0
C2408 a_9705_12861# a_10761_14767# 0
C2409 a_4032_5043# a_3229_5051# 0.04911f
C2410 a_14432_4521# a_13186_4919# 0
C2411 a_12430_4527# a_12655_4919# 0.00559f
C2412 a_16539_5473# a_16275_5473# 0
C2413 a_6238_6077# a_6261_5043# 0
C2414 a_14982_22987# a_14541_22875# 0.11299f
C2415 a_10953_14739# a_11501_15239# 0.08954f
C2416 a_12227_2049# a_12281_2159# 0.03622f
C2417 a_6208_2817# a_10916_4597# 0
C2418 a_4477_5409# a_4309_5409# 0
C2419 a_17096_23241# a_16823_22875# 0.07715f
C2420 a_6003_11935# a_4905_12113# 0.18489f
C2421 a_18663_27017# a_18671_29108# 0
C2422 a_14545_5833# a_14377_5833# 0
C2423 a_4423_5299# a_6036_5017# 0.00419f
C2424 a_5975_12927# a_4849_11293# 0.18585f
C2425 a_5975_12927# a_5851_13769# 0
C2426 a_6036_5017# VDPWR 0.35121f
C2427 a_23133_17137# VDPWR 0.92242f
C2428 a_16471_17161# a_16486_16197# 0.02069f
C2429 a_20877_17147# VDPWR 0.35105f
C2430 a_16793_4785# a_17544_4529# 0.00682f
C2431 a_16094_5473# VDPWR 0.16911f
C2432 sky130_fd_sc_hd__dfxbp_1_5.Q_N a_19059_25272# 0.00125f
C2433 sky130_fd_sc_hd__dfxbp_1_7.Q a_18689_26867# 0
C2434 a_10525_5837# VDPWR 0.00694f
C2435 a_7113_13395# a_6944_13645# 0
C2436 a_4329_2043# a_5080_2153# 0.00696f
C2437 a_18663_27120# a_19055_27097# 0
C2438 a_9705_12861# a_12039_15239# 0.00585f
C2439 a_18667_24874# VDPWR 0.191f
C2440 a_9556_17271# a_23511_14335# 0.04403f
C2441 a_14281_5833# a_14545_5833# 0
C2442 a_4849_11293# a_4513_14775# 0.00146f
C2443 a_9503_10581# a_9493_12145# 0
C2444 a_18667_31449# a_18667_32557# 0
C2445 a_4309_5409# a_2217_5025# 0
C2446 a_9705_12861# a_12615_14007# 0
C2447 ui_in[3] ui_in[4] 0.03102f
C2448 a_14940_22875# sky130_fd_sc_hd__dfxbp_1_4.CLK 0
C2449 a_10108_4597# VDPWR 0.12354f
C2450 sky130_fd_sc_hd__dfxbp_1_1.Q_N a_9943_22879# 0.11931f
C2451 a_14541_22875# sky130_fd_sc_hd__dfxbp_1_3.CLK 0.01405f
C2452 a_9379_14779# a_9369_16343# 0.00102f
C2453 sky130_fd_sc_hd__dfxbp_1_4.Q_N a_18120_23197# 0.12801f
C2454 sky130_fd_sc_hd__dfxbp_1_8.Q_N sky130_fd_sc_hd__inv_4_0.A 0
C2455 a_15242_5833# a_14491_5723# 0.00696f
C2456 a_6238_6077# a_16371_5473# 0
C2457 a_4625_15373# a_4513_14775# 0
C2458 VDPWR a_10955_11939# 0
C2459 a_10499_4853# VDPWR 0.71029f
C2460 a_4711_15373# a_4903_15345# 0.00101f
C2461 a_15711_4547# VDPWR 1.46429f
C2462 a_11255_13773# a_11728_13649# 0.24537f
C2463 a_10508_22879# a_10550_22991# 0
C2464 a_4755_13107# a_4627_12141# 0
C2465 a_6238_6077# a_10261_5471# 0
C2466 a_6281_2043# a_6335_2153# 0.03622f
C2467 sky130_fd_sc_hd__dfxbp_1_8.Q_N a_18667_34259# 0.12218f
C2468 a_6208_2817# a_10025_2159# 0
C2469 uo_out[2] VDPWR 0
C2470 a_23731_14309# a_23133_17137# 0.08898f
C2471 a_4084_5017# a_2289_5307# 0.00286f
C2472 ui_in[5] ui_in[4] 0.03102f
C2473 a_1920_1765# a_2049_2157# 0.00792f
C2474 a_6165_5409# VDPWR 0
C2475 a_6003_11935# a_4849_11293# 0.10273f
C2476 a_15407_23143# a_14375_22875# 0.04808f
C2477 a_14377_5833# VDPWR 0
C2478 a_21491_17145# VDPWR 0.46902f
C2479 a_16275_5473# VDPWR 0.00116f
C2480 a_10550_22991# a_10297_22879# 0
C2481 a_9369_16343# a_8193_13753# 0.00258f
C2482 a_8283_2049# a_8700_2159# 0.06611f
C2483 a_15693_17123# sky130_fd_sc_hd__dfxbp_1_0.CLK 0.02023f
C2484 a_12587_5825# a_12533_5715# 0.03622f
C2485 a_6238_6077# a_15522_4913# 0
C2486 a_4595_14775# a_4903_15345# 0
C2487 a_18663_27756# a_18663_27545# 0.31062f
C2488 a_19059_31950# VDPWR 0
C2489 a_11147_11911# a_9771_12117# 0.03573f
C2490 a_23677_14701# a_23761_14335# 0.0594f
C2491 a_7113_13395# a_7173_15235# 0.41047f
C2492 a_4847_14525# a_6717_15235# 0.00159f
C2493 a_9705_12861# a_11979_13399# 0.00446f
C2494 a_16297_1793# VDPWR 0.18607f
C2495 VDPWR a_4383_2153# 0.0097f
C2496 sky130_fd_sc_hd__dfxbp_1_5.Q_N a_18667_25006# 0.04247f
C2497 a_14281_5833# VDPWR 0
C2498 sky130_fd_sc_hd__dfxbp_1_6.Q_N a_18667_31354# 0.0011f
C2499 a_23511_14701# VDPWR 0.10426f
C2500 a_6238_6077# a_8431_5049# 0
C2501 a_11777_15239# a_9703_16093# 0.00241f
C2502 sky130_fd_sc_hd__dfxbp_1_7.Q a_18671_29438# 0
C2503 a_8561_23241# a_7863_22875# 0.19462f
C2504 a_16657_22875# a_15838_23197# 0
C2505 a_6944_13645# a_6862_13645# 0.00477f
C2506 a_3040_5417# VDPWR 0
C2507 VDPWR sky130_fd_sc_hd__dfxbp_1_0.CLK 0.41675f
C2508 a_4905_12113# VDPWR 0.43561f
C2509 a_12587_5459# a_14152_5441# 0
C2510 a_8794_5415# a_10132_5445# 0
C2511 a_10869_11939# a_10841_12931# 0
C2512 a_9579_12145# a_9493_12145# 0.00658f
C2513 a_17096_23241# a_17011_22875# 0.03733f
C2514 a_4765_11543# a_4627_12141# 0
C2515 a_6087_14735# a_6717_15235# 0.00232f
C2516 a_18693_24801# a_18693_24621# 0.00123f
C2517 a_5363_5043# a_6165_5043# 0
C2518 a_11175_1793# a_12227_2049# 0.21187f
C2519 a_4721_13809# VDPWR 0.003f
C2520 a_9713_14529# a_9703_16093# 0.46421f
C2521 a_14545_5467# a_16146_5447# 0
C2522 sky130_fd_sc_hd__dfxbp_1_9.Q a_19059_31950# 0
C2523 a_6238_6077# a_12587_5825# 0.00113f
C2524 a_6238_6077# a_7126_5409# 0
C2525 a_12587_5459# a_12533_5715# 0.00386f
C2526 a_13077_23237# a_12295_22871# 0
C2527 a_10553_4597# a_10916_4597# 0.00985f
C2528 sky130_fd_sc_hd__dfxbp_1_7.Q sky130_fd_sc_hd__dfxbp_1_6.Q_N 0.01749f
C2529 a_18667_31552# a_18667_32188# 0.03684f
C2530 a_2343_5051# a_2217_5025# 0.0842f
C2531 sky130_fd_sc_hd__dfxbp_1_9.CLK a_18667_32188# 0
C2532 a_14982_22987# a_14729_22875# 0
C2533 a_6208_2817# a_11250_4597# 0
C2534 a_12227_2049# a_13840_1767# 0.00419f
C2535 a_9317_5049# a_11439_4597# 0.04997f
C2536 a_10761_14767# a_9769_15349# 0
C2537 a_11255_13773# a_10799_13773# 0
C2538 a_10761_14767# VDPWR 0
C2539 a_10869_11939# a_9703_16093# 0
C2540 VDPWR a_16823_22875# 0.31438f
C2541 a_10382_23245# VDPWR 0.25536f
C2542 a_5269_1787# a_6335_1787# 0.08312f
C2543 VDPWR a_6335_2153# 0.00967f
C2544 a_7944_1767# a_6698_1787# 0
C2545 a_6238_6077# ui_in[0] 0.07426f
C2546 VDPWR a_12017_2159# 0
C2547 a_10132_5445# VDPWR 0.35066f
C2548 ui_in[6] ui_in[5] 0.03102f
C2549 a_14432_4521# a_14657_4913# 0.00559f
C2550 a_13520_4919# a_13709_4553# 0
C2551 a_11222_5471# VDPWR 0
C2552 a_11255_13773# a_8193_13753# 0
C2553 a_6208_2817# a_12281_2159# 0
C2554 a_4329_2043# a_4215_2153# 0
C2555 a_19059_31950# a_18667_31977# 0
C2556 a_23731_14309# a_23511_14701# 0.00549f
C2557 a_17689_23143# VDPWR 0.51106f
C2558 a_23731_14309# sky130_fd_sc_hd__dfxbp_1_0.CLK 0
C2559 a_12227_2049# a_12644_2159# 0.06611f
C2560 a_9896_1767# a_10121_2159# 0.00559f
C2561 a_23133_17137# a_23677_14335# 0
C2562 sky130_fd_sc_hd__dfxbp_1_4.CLK a_17096_23241# 0
C2563 a_11501_15239# a_11583_15239# 0.00578f
C2564 a_18625_5265# a_6238_6077# 0
C2565 a_11439_4597# a_12823_4919# 0.04534f
C2566 a_14179_2049# a_13840_1767# 0.04737f
C2567 a_9371_13111# a_9493_12145# 0.00144f
C2568 a_24774_14701# a_24962_14701# 0.10432f
C2569 a_6238_6077# a_12587_5459# 0
C2570 a_6087_14735# a_6329_12927# 0
C2571 a_18839_4938# VDPWR 0.00182f
C2572 a_7697_22875# a_8304_22987# 0.14145f
C2573 sky130_fd_sc_hd__dfxbp_1_7.Q a_18663_27252# 0
C2574 a_9128_5049# VDPWR 0
C2575 a_12039_15239# a_9769_15349# 0
C2576 a_10357_5471# VDPWR 0
C2577 a_11255_13773# a_9779_13785# 0
C2578 a_14982_22987# a_15239_23241# 0.03684f
C2579 sky130_fd_sc_hd__dfxbp_1_3.CLK a_14729_22875# 0
C2580 a_12039_15239# VDPWR 0.83278f
C2581 a_6805_15235# a_4837_16089# 0
C2582 a_4849_11293# VDPWR 1.0316f
C2583 VDPWR a_5851_13769# 0.44659f
C2584 a_2343_5417# a_2289_5307# 0.03622f
C2585 a_12615_14007# VDPWR 0.13186f
C2586 a_2187_1765# a_2676_1791# 0.08982f
C2587 a_16902_5473# a_15431_5467# 0.08907f
C2588 VDPWR a_4119_1787# 0.00116f
C2589 a_18671_29306# a_18671_29942# 0.03684f
C2590 a_6208_2817# a_16660_1793# 0.00236f
C2591 a_15711_4547# a_16454_4503# 0.11874f
C2592 a_6698_2153# a_6335_2153# 0.00847f
C2593 a_12113_1793# a_11175_1793# 0
C2594 a_4625_15373# VDPWR 0.45106f
C2595 a_6375_5299# a_6238_6077# 0.00299f
C2596 a_18697_29647# sky130_fd_sc_hd__dfxbp_1_6.Q_N 0
C2597 a_18667_31449# a_18671_29108# 0
C2598 a_4849_11293# a_4763_14775# 0
C2599 a_6238_6077# a_16371_5839# 0
C2600 a_12978_2159# VDPWR 0
C2601 a_10652_1793# a_10235_2049# 0.03016f
C2602 a_12533_5715# a_11439_4597# 0
C2603 sky130_fd_sc_hd__dfxbp_1_8.Q_N a_18667_34470# 0.09273f
C2604 sky130_fd_sc_hd__dfxbp_1_2.CLK a_9943_22879# 0
C2605 a_4505_13107# a_4913_13781# 0
C2606 a_13167_1793# a_14233_2159# 0.04534f
C2607 a_18671_29306# a_19063_29704# 0
C2608 a_4763_14775# a_4625_15373# 0
C2609 a_18689_26867# a_18667_25299# 0
C2610 a_9317_5049# a_10499_4853# 0
C2611 a_9317_5049# a_15711_4547# 0.03484f
C2612 a_9631_11547# a_9493_12145# 0
C2613 a_15239_23241# sky130_fd_sc_hd__dfxbp_1_3.CLK 0
C2614 a_17236_5473# VDPWR 0
C2615 a_18667_31552# a_19059_31529# 0
C2616 a_18671_29306# VDPWR 0.19099f
C2617 sky130_fd_sc_hd__dfxbp_1_1.Q_N a_8729_23143# 0
C2618 sky130_fd_sc_hd__dfxbp_1_9.CLK a_19059_31529# 0
C2619 a_2187_1765# a_6071_2153# 0
C2620 a_17425_5473# a_18625_5265# 0.0056f
C2621 VDPWR a_4746_1787# 0.21795f
C2622 a_8038_5023# a_8167_5415# 0.00792f
C2623 a_15711_4547# a_16793_4785# 0.21188f
C2624 a_20877_17147# a_19235_17155# 0
C2625 sky130_fd_sc_hd__inv_2_0.A a_19059_34232# 0
C2626 a_17264_22987# sky130_fd_sc_hd__dfxbp_1_4.Q_N 0.05782f
C2627 uio_out[7] uio_out[6] 0.03102f
C2628 a_9769_15349# a_11979_13399# 0
C2629 a_4847_14525# a_6629_15387# 0.29596f
C2630 a_11250_4963# VDPWR 0
C2631 a_11979_13399# VDPWR 0.49382f
C2632 a_3229_5051# a_5363_5043# 0
C2633 sky130_fd_sc_hd__dfxbp_1_5.Q_N a_18667_25299# 0.12218f
C2634 a_6238_6077# a_11439_4597# 0
C2635 a_13284_5825# a_12533_5715# 0.00696f
C2636 a_17011_22875# VDPWR 0.07693f
C2637 sky130_fd_sc_hd__dfxbp_1_5.CLK a_18667_24874# 0
C2638 a_8283_2049# VDPWR 0.45035f
C2639 a_8283_2049# a_9034_2159# 0.00696f
C2640 a_12323_5825# a_12194_5433# 0.00792f
C2641 sky130_fd_sc_hd__dfxbp_1_7.Q sky130_fd_sc_hd__dfxbp_1_7.Q_N 0.15319f
C2642 a_12129_22871# a_11406_23201# 0
C2643 a_4627_12141# a_6281_11907# 0
C2644 a_4329_2043# a_3990_1761# 0.04737f
C2645 a_6629_15387# a_6087_14735# 0.09734f
C2646 a_10289_4597# VDPWR 0.00151f
C2647 a_5269_1787# a_5080_2153# 0
C2648 a_9705_12861# a_9501_13813# 0.00246f
C2649 a_18667_31449# a_18667_31552# 0.14145f
C2650 a_18667_31449# sky130_fd_sc_hd__dfxbp_1_9.CLK 0.25091f
C2651 a_6208_2817# a_11175_1793# 0.00288f
C2652 a_12419_5825# a_12194_5433# 0.00559f
C2653 a_18663_27017# a_18663_27756# 0.03218f
C2654 a_18667_24676# a_18667_25510# 0.19462f
C2655 a_12736_22983# a_12568_23237# 0.23992f
C2656 a_9379_14779# a_9629_14529# 0.00723f
C2657 a_9781_10553# a_9381_11547# 0
C2658 sky130_fd_sc_hd__dfxbp_1_1.CLK a_10807_23245# 0
C2659 a_11888_1767# a_12113_2159# 0.00559f
C2660 a_9223_1793# VDPWR 1.38873f
C2661 a_6208_2817# a_13840_1767# 0.00211f
C2662 a_5809_14763# a_4913_13781# 0
C2663 a_9223_1793# a_9034_2159# 0
C2664 a_15711_4547# a_16847_4895# 0.04534f
C2665 a_4329_2043# a_4383_1787# 0.00386f
C2666 a_14432_4521# a_14771_4803# 0.04737f
C2667 a_6635_15235# VDPWR 0.42362f
C2668 a_9715_11297# a_10955_11939# 0
C2669 a_2259_2047# a_1920_1765# 0.04737f
C2670 a_6238_6077# a_13284_5825# 0
C2671 a_6238_6077# a_6036_5017# 0
C2672 a_6238_6077# a_23133_17137# 0.00495f
C2673 a_8038_5023# a_7986_5049# 0.1439f
C2674 a_14771_4803# a_15188_4913# 0.06611f
C2675 a_10385_4963# a_10499_4853# 0
C2676 a_21491_17145# a_19235_17155# 0
C2677 VDPWR a_10477_23245# 0.00347f
C2678 a_14152_5441# a_14377_5833# 0.00559f
C2679 sky130_fd_sc_hd__dfxbp_1_4.CLK VDPWR 0.2713f
C2680 a_14179_2049# a_14596_2159# 0.06611f
C2681 a_18667_25879# sky130_fd_sc_hd__dfxbp_1_7.CLK 0.20774f
C2682 a_8687_22875# sky130_fd_sc_hd__dfxbp_1_1.CLK 0
C2683 a_6238_6077# a_16094_5473# 0.0031f
C2684 a_9587_13813# a_9501_13813# 0.00658f
C2685 a_8561_23241# VDPWR 0.19824f
C2686 a_6429_5043# VDPWR 0.18612f
C2687 a_6238_6077# a_10525_5837# 0.0014f
C2688 a_16275_5839# a_16146_5447# 0.00792f
C2689 a_6208_2817# a_12644_2159# 0
C2690 a_18671_29731# sky130_fd_sc_hd__dfxbp_1_9.Q_N 0
C2691 a_10289_4963# a_10108_4597# 0
C2692 a_8377_5305# a_10160_4571# 0
C2693 a_9317_5049# a_10132_5445# 0
C2694 a_9491_15377# a_9703_16093# 0
C2695 a_10289_1793# VDPWR 0.18611f
C2696 a_4755_13107# a_4513_14775# 0
C2697 a_12568_23237# a_12483_22871# 0.03733f
C2698 a_4477_5043# a_4309_5043# 0
C2699 a_17733_4529# a_17210_4529# 0
C2700 a_6238_6077# a_10108_4597# 0
C2701 a_7986_5049# a_7315_5043# 0.05015f
C2702 a_14771_4803# a_13709_4553# 0.21188f
C2703 a_11501_15239# a_9703_16093# 0.232f
C2704 a_2187_1765# a_4215_1787# 0
C2705 a_14281_5833# a_14152_5441# 0.00792f
C2706 VDPWR a_12568_23237# 0.25518f
C2707 a_19235_17155# sky130_fd_sc_hd__dfxbp_1_0.CLK 0.02511f
C2708 a_1920_1765# a_2313_2157# 0.02301f
C2709 ui_in[6] ui_in[7] 0.03102f
C2710 sky130_fd_sc_hd__dfxbp_1_4.Q_N sky130_fd_sc_hd__dfxbp_1_3.Q_N 0
C2711 a_16902_5473# a_16539_5473# 0.00985f
C2712 a_12655_4919# a_12769_4809# 0
C2713 a_10499_4853# a_6238_6077# 0
C2714 a_7697_22875# a_7863_22875# 0.96835f
C2715 a_9317_5049# a_18839_4938# 0.00688f
C2716 a_15711_4547# a_6238_6077# 0
C2717 a_11411_5471# VDPWR 1.42163f
C2718 a_5975_12927# a_6129_12927# 0.00401f
C2719 a_11810_13649# a_11979_13399# 0
C2720 a_14281_5467# VDPWR 0.00104f
C2721 a_6911_15235# a_7173_15235# 0
C2722 a_6238_6077# a_14377_5833# 0
C2723 a_15904_1767# a_15852_1793# 0.1439f
C2724 uo_out[3] uo_out[4] 0.03102f
C2725 a_6238_6077# a_16275_5473# 0
C2726 a_17521_23241# a_17264_22987# 0.03684f
C2727 a_4213_5043# VDPWR 0.00116f
C2728 sky130_fd_sc_hd__dfxbp_1_5.CLK a_16823_22875# 0
C2729 a_14982_22987# sky130_fd_sc_hd__dfxbp_1_3.CLK 0
C2730 a_15693_17123# a_17345_17163# 0
C2731 a_10499_4853# a_10916_4963# 0.06611f
C2732 a_18663_27545# a_18663_26922# 0.03136f
C2733 a_12227_2049# a_12978_1793# 0.00682f
C2734 a_16583_4529# a_16847_4529# 0
C2735 a_18667_31552# a_18667_31684# 0.23675f
C2736 sky130_fd_sc_hd__dfxbp_1_9.CLK a_18667_31684# 0
C2737 a_6208_2817# a_12378_4553# 0
C2738 a_13592_23193# VDPWR 0.21267f
C2739 a_6389_13769# a_4915_10549# 0.00248f
C2740 a_18671_29306# a_18671_29203# 0.14145f
C2741 a_10869_11939# a_9493_12145# 0
C2742 a_10761_14767# a_9715_11297# 0.00121f
C2743 a_12950_5825# a_12587_5825# 0.00847f
C2744 a_6208_2817# a_13969_1793# 0
C2745 a_8169_2159# a_8337_2159# 0
C2746 sky130_fd_sc_hd__dfxbp_1_5.CLK a_17689_23143# 0.12068f
C2747 a_14375_22875# a_12736_22983# 0
C2748 a_14281_5833# a_6238_6077# 0
C2749 a_6238_6077# a_23511_14701# 0.00106f
C2750 a_16679_4529# VDPWR 0
C2751 a_6238_6077# sky130_fd_sc_hd__dfxbp_1_0.CLK 0
C2752 a_17345_17163# VDPWR 0.42372f
C2753 a_9705_12861# a_11147_11911# 0.02321f
C2754 a_8169_1793# VDPWR 0
C2755 a_5942_1761# a_2187_1765# 0.001f
C2756 a_14545_5833# a_14908_5833# 0.00847f
C2757 a_4915_10549# a_7831_14003# 0
C2758 a_23761_14335# VDPWR 0.09737f
C2759 a_10986_2159# VDPWR 0
C2760 a_2706_5417# VDPWR 0.021f
C2761 a_6208_2817# a_6698_1787# 0
C2762 a_5942_1761# a_6071_2153# 0.00792f
C2763 a_4423_5299# a_4477_5409# 0.03622f
C2764 a_17425_5473# a_15711_4547# 0
C2765 a_12950_5459# a_12587_5459# 0.00985f
C2766 a_4477_5409# VDPWR 0.0096f
C2767 a_16660_2159# a_16297_2159# 0.00847f
C2768 a_11411_5471# a_10888_5471# 0
C2769 a_9769_15349# a_9501_13813# 0.00159f
C2770 a_6127_13769# a_4839_12857# 0.00253f
C2771 a_9896_1767# a_6208_2817# 0.00211f
C2772 a_16902_5473# VDPWR 0.21501f
C2773 VDPWR a_9501_13813# 0.43907f
C2774 a_12039_15239# a_9715_11297# 0
C2775 a_18667_34259# a_18667_33731# 0.04808f
C2776 ui_in[1] ui_in[0] 5.54574f
C2777 a_10975_23147# a_12129_22871# 0
C2778 a_9705_12861# a_9771_12117# 0.04364f
C2779 a_10550_22991# sky130_fd_sc_hd__dfxbp_1_1.CLK 0
C2780 a_12129_22871# a_12736_22983# 0.14145f
C2781 a_6208_2817# a_14596_2159# 0
C2782 a_15904_1767# a_16129_2159# 0.00559f
C2783 a_9381_11547# a_9503_10581# 0.00144f
C2784 a_7944_1767# a_8073_2159# 0.00792f
C2785 a_6208_2817# a_14432_4521# 0
C2786 a_6238_6077# a_10132_5445# 0.00451f
C2787 a_12419_5459# VDPWR 0
C2788 a_6238_6077# a_11222_5471# 0
C2789 a_14375_22875# VDPWR 0.66219f
C2790 a_2313_1791# VDPWR 0.18286f
C2791 a_18667_33636# a_18693_34175# 0
C2792 a_16657_22875# a_18120_23197# 0
C2793 a_4423_5299# a_2217_5025# 0.00303f
C2794 a_18671_30311# VDPWR 0.21282f
C2795 a_2217_5025# VDPWR 1.57816f
C2796 a_16471_17161# a_18113_17153# 0
C2797 a_9781_10553# a_11255_13773# 0.00248f
C2798 sky130_fd_sc_hd__dfxbp_1_7.Q_N a_18667_25299# 0
C2799 a_7863_22875# a_8304_22987# 0.11299f
C2800 a_17521_23241# sky130_fd_sc_hd__dfxbp_1_3.Q_N 0
C2801 a_5363_5043# a_5984_5043# 0.05065f
C2802 a_18839_4938# a_6238_6077# 0.0023f
C2803 a_23731_14309# a_23761_14335# 0.35203f
C2804 a_9128_5049# a_6238_6077# 0
C2805 a_18625_4938# VDPWR 0.11729f
C2806 a_12430_4527# a_11439_4597# 0.1189f
C2807 a_10357_5471# a_6238_6077# 0
C2808 a_16660_2159# a_6208_2817# 0.00205f
C2809 a_4755_13107# VDPWR 0.33272f
C2810 a_6208_2817# a_13709_4553# 0
C2811 a_12559_4553# a_11439_4597# 0
C2812 sky130_fd_sc_hd__dfxbp_1_4.CLK a_14814_23241# 0
C2813 a_14908_5833# VDPWR 0.02196f
C2814 a_6087_14735# a_6862_13645# 0
C2815 a_12129_22871# a_12483_22871# 0.06222f
C2816 a_8377_5305# a_10525_5471# 0
C2817 sky130_fd_sc_hd__dfxbp_1_5.CLK a_17011_22875# 0
C2818 a_11222_5837# VDPWR 0
C2819 a_20384_16179# a_20877_17147# 0.01375f
C2820 a_6127_13769# a_4837_16089# 0.00702f
C2821 a_20109_17157# a_19510_16177# 0
C2822 a_13520_4553# VDPWR 0
C2823 a_12129_22871# VDPWR 0.66338f
C2824 a_10550_22991# a_10807_23245# 0.03684f
C2825 sky130_fd_sc_hd__dfxbp_1_4.Q_N a_17647_22875# 0.00125f
C2826 a_9715_11297# a_11979_13399# 0.00118f
C2827 a_15119_1793# a_16660_1793# 0.08907f
C2828 a_6805_15235# a_6635_15235# 0.00167f
C2829 a_12950_5459# a_11439_4597# 0
C2830 a_6208_2817# a_13969_2159# 0
C2831 a_6208_2817# a_24962_14701# 0.00237f
C2832 a_6375_5299# a_8431_5415# 0
C2833 a_5975_12927# a_6281_11907# 0
C2834 a_12865_14007# a_9556_17271# 0
C2835 a_17544_4895# VDPWR 0
C2836 sky130_fd_sc_hd__inv_12_0.A sky130_fd_sc_hd__inv_8_0.A 0.96515f
C2837 a_12295_22871# a_12993_23237# 0.19462f
C2838 a_11411_5471# a_9317_5049# 0.05944f
C2839 a_10160_4571# VDPWR 0.4471f
C2840 uio_in[0] ui_in[7] 0.03102f
C2841 a_15431_5467# a_16539_5839# 0.04534f
C2842 a_6003_11935# a_4627_12141# 0
C2843 a_15522_4547# VDPWR 0
C2844 sky130_fd_sc_hd__dfxbp_1_0.Q_N a_10109_22879# 0.0011f
C2845 a_6129_12927# VDPWR 0
C2846 a_6238_6077# a_17236_5473# 0
C2847 a_18667_32188# a_18667_33731# 0
C2848 a_6208_2817# a_12978_1793# 0
C2849 sky130_fd_sc_hd__dfxbp_1_5.CLK sky130_fd_sc_hd__dfxbp_1_4.CLK 0.00149f
C2850 a_4084_5017# a_4477_5043# 0.02283f
C2851 a_4765_11543# VDPWR 0.33144f
C2852 a_13284_5459# VDPWR 0
C2853 a_16454_4503# a_16679_4529# 0.00487f
C2854 a_16847_4529# VDPWR 0.18786f
C2855 a_19063_29283# a_18671_29306# 0
C2856 a_20384_16179# a_21491_17145# 0
C2857 sky130_fd_sc_hd__dfxbp_1_5.Q_N a_18667_24676# 0.51145f
C2858 a_7697_22875# VDPWR 0.65176f
C2859 a_10499_4853# a_12430_4527# 0.00138f
C2860 a_11147_11911# VDPWR 0.29962f
C2861 a_9713_14529# a_9629_14779# 0.07979f
C2862 a_7697_22875# a_9160_23197# 0
C2863 a_23761_14335# a_23677_14335# 0
C2864 a_18693_25215# a_18667_24874# 0
C2865 a_10025_2159# a_10289_2159# 0
C2866 a_18663_27017# a_18663_26922# 0.96835f
C2867 a_16402_4529# a_15431_5467# 0
C2868 a_9381_11547# a_9371_13111# 0.00102f
C2869 a_16033_1793# VDPWR 0.00115f
C2870 a_6003_11935# a_6281_11907# 0.11706f
C2871 a_4119_2153# a_3938_1787# 0
C2872 VDPWR sky130_fd_sc_hd__dfxbp_1_7.CLK 0.27419f
C2873 a_9369_16343# a_9451_16343# 0.00641f
C2874 a_16793_4785# a_16679_4529# 0
C2875 ui_in[1] a_23133_17137# 0
C2876 VDPWR a_9771_12117# 0.43751f
C2877 a_18667_33731# a_18667_34470# 0.03218f
C2878 a_16485_5729# a_16146_5447# 0.04737f
C2879 a_14281_5467# a_14152_5441# 0.00758f
C2880 sky130_fd_sc_hd__dfxbp_1_2.Q_N a_12568_23237# 0.04247f
C2881 a_11411_5471# a_12533_5715# 0.21188f
C2882 a_13284_5825# a_13473_5459# 0
C2883 a_6389_13769# a_4839_12857# 0.04676f
C2884 a_18667_31552# a_19059_31950# 0
C2885 a_17425_5473# a_17236_5473# 0
C2886 a_18667_24874# a_18693_24621# 0
C2887 sky130_fd_sc_hd__inv_12_0.A sky130_fd_sc_hd__inv_6_0.A 0
C2888 a_19059_31950# sky130_fd_sc_hd__dfxbp_1_9.CLK 0
C2889 a_18693_34175# a_18667_33834# 0
C2890 a_7927_14003# a_4915_10549# 0
C2891 a_9556_17271# ui_in[0] 0.00107f
C2892 uio_in[0] uio_in[1] 0.03102f
C2893 a_18671_30311# a_18671_29203# 0
C2894 a_6429_5043# a_6238_6077# 0
C2895 a_24152_14385# VDPWR 0.00498f
C2896 a_1950_5025# a_2343_5417# 0.02301f
C2897 a_11836_1793# a_12017_2159# 0
C2898 a_4847_14525# a_4913_13781# 0.0012f
C2899 a_17521_23241# a_17647_22875# 0.00617f
C2900 a_14375_22875# a_14814_23241# 0.27314f
C2901 a_12113_2159# VDPWR 0
C2902 a_9381_11547# a_9631_11547# 0.02504f
C2903 a_9491_15377# a_9619_16343# 0
C2904 a_4423_5299# a_4309_5409# 0
C2905 a_8136_23241# sky130_fd_sc_hd__dfxbp_1_0.Q_N 0.04247f
C2906 sky130_fd_sc_hd__dfxbp_1_7.Q_N a_19055_27518# 0.00125f
C2907 a_4627_12141# VDPWR 0.445f
C2908 a_4309_5409# VDPWR 0
C2909 a_6087_14735# a_4913_13781# 0
C2910 a_17345_17163# a_19235_17155# 0
C2911 a_14771_4803# a_14657_4913# 0
C2912 a_11411_5471# a_6238_6077# 0.00691f
C2913 a_10025_1793# a_9896_1767# 0.00758f
C2914 a_9317_5049# a_18625_4938# 0.31816f
C2915 a_13592_23193# sky130_fd_sc_hd__dfxbp_1_2.Q_N 0.12801f
C2916 a_15711_4547# a_15188_4547# 0
C2917 a_10953_14739# a_10761_14767# 0
C2918 a_6792_5409# a_5363_5043# 0.03325f
C2919 a_13119_22871# a_13161_23139# 0
C2920 uio_in[4] uio_in[3] 0.03102f
C2921 a_6238_6077# a_14281_5467# 0
C2922 a_18667_33636# a_18667_33834# 0.1111f
C2923 a_8193_13753# a_7749_14003# 0.10797f
C2924 a_2187_1765# a_6208_2817# 0.11803f
C2925 a_14179_2049# a_14930_2159# 0.00696f
C2926 a_11810_13649# a_11147_11911# 0
C2927 a_4915_10549# a_7999_14003# 0
C2928 a_17264_22987# a_16657_22875# 0.14145f
C2929 a_18625_4938# a_16793_4785# 0
C2930 a_6698_1787# a_6335_1787# 0.00985f
C2931 a_6087_14735# a_6911_15235# 0.00651f
C2932 a_6389_13769# a_4837_16089# 0.00515f
C2933 a_23731_14309# a_24152_14385# 0.01881f
C2934 a_4213_5409# a_4477_5409# 0
C2935 sky130_fd_sc_hd__dfxbp_1_2.CLK a_12694_22871# 0
C2936 a_18667_31449# a_18667_33731# 0
C2937 a_10717_13773# a_12039_15239# 0
C2938 a_10382_23245# a_9943_22879# 0.27314f
C2939 sky130_fd_sc_hd__dfxbp_1_4.CLK a_15365_22875# 0
C2940 a_8561_23241# a_8645_23241# 0.00851f
C2941 a_18671_29306# a_18671_29108# 0.1111f
C2942 a_2289_5307# a_3040_5417# 0.00696f
C2943 a_9715_11297# a_9501_13813# 0.00317f
C2944 VDPWR a_8304_22987# 0.19095f
C2945 sky130_fd_sc_hd__dfxbp_1_0.Q_N a_8051_22875# 0.142f
C2946 a_15407_23143# VDPWR 0.51272f
C2947 sky130_fd_sc_hd__inv_2_0.A sky130_fd_sc_hd__inv_4_0.A 0.14042f
C2948 a_8283_2049# a_8700_1793# 0.03016f
C2949 a_10717_13773# a_12615_14007# 0
C2950 a_10525_5471# VDPWR 0.18051f
C2951 a_14179_2049# a_14596_1793# 0.03016f
C2952 a_10953_14739# a_12039_15239# 0.00327f
C2953 ui_in[1] sky130_fd_sc_hd__dfxbp_1_0.CLK 0.31497f
C2954 a_16454_4503# a_16847_4529# 0.02283f
C2955 a_8038_5023# a_8431_5049# 0.02283f
C2956 a_6281_11907# VDPWR 0.30386f
C2957 a_9317_5049# a_10160_4571# 0
C2958 sky130_fd_sc_hd__inv_2_0.A a_18667_34259# 0.12052f
C2959 a_18667_31449# a_18693_31299# 0.06222f
C2960 a_12533_5715# a_12419_5459# 0
C2961 a_12587_5825# a_12769_4809# 0
C2962 sky130_fd_sc_hd__inv_2_0.A sky130_fd_sc_hd__inv_6_0.A 0
C2963 a_6127_13769# a_4849_11293# 0
C2964 a_9379_14779# a_10675_14767# 0
C2965 a_6127_13769# a_5851_13769# 0.00119f
C2966 VDPWR a_4587_13107# 0.02522f
C2967 a_9896_1767# a_10121_1793# 0.00487f
C2968 a_12993_23237# a_13161_23139# 0.31062f
C2969 a_4213_5409# a_2217_5025# 0
C2970 a_16793_4785# a_17544_4895# 0.00696f
C2971 sky130_fd_sc_hd__dfxbp_1_0.Q_N a_10297_22879# 0
C2972 a_9779_13785# a_11728_13649# 0
C2973 a_15904_1767# a_16243_2049# 0.04737f
C2974 a_6238_6077# a_23761_14335# 0.07254f
C2975 a_14375_22875# sky130_fd_sc_hd__dfxbp_1_2.Q_N 0.00248f
C2976 a_9223_1793# a_10235_2049# 0.21187f
C2977 a_6208_2817# a_8073_2159# 0
C2978 a_9223_1793# a_8700_1793# 0
C2979 uo_out[0] uo_out[1] 0.03102f
C2980 a_16094_5473# a_14491_5723# 0
C2981 a_12281_1793# a_11888_1767# 0.02283f
C2982 a_8431_5049# a_7315_5043# 0.08313f
C2983 a_16902_5473# a_6238_6077# 0
C2984 a_11888_1767# VDPWR 0.34955f
C2985 uio_out[0] uio_out[1] 0.03102f
C2986 a_12533_5715# a_14908_5833# 0
C2987 a_12615_14007# a_12793_14007# 0.00412f
C2988 a_18693_34175# VDPWR 0.00627f
C2989 a_2343_5051# VDPWR 0.18537f
C2990 a_8193_13753# a_10675_14767# 0
C2991 a_9703_16093# a_9619_16093# 0.00234f
C2992 a_4503_16339# a_4753_16089# 0.00723f
C2993 a_16793_4785# a_16847_4529# 0.00386f
C2994 a_9379_14779# a_8193_13753# 0.00206f
C2995 a_6238_6077# a_12419_5459# 0
C2996 a_6208_2817# a_24774_14701# 0.00556f
C2997 a_12587_5459# a_12769_4809# 0
C2998 a_16539_5473# a_15431_5467# 0.08313f
C2999 a_23677_14701# VDPWR 0.20475f
C3000 a_9577_15377# a_9769_15349# 0.00101f
C3001 a_14100_5467# VDPWR 0.15904f
C3002 a_10235_2049# a_10289_1793# 0.00386f
C3003 a_10717_13773# a_11979_13399# 0
C3004 a_9577_15377# VDPWR 0.00333f
C3005 a_7315_5043# a_7126_5409# 0
C3006 a_18671_29306# sky130_fd_sc_hd__dfxbp_1_9.CLK 0
C3007 sky130_fd_sc_hd__dfxbp_1_7.Q a_18663_27545# 0.1234f
C3008 uio_out[1] uio_out[2] 0.03102f
C3009 a_12129_22871# sky130_fd_sc_hd__dfxbp_1_2.Q_N 0.11931f
C3010 a_13167_1793# a_13788_1793# 0.05049f
C3011 a_6238_6077# a_2217_5025# 0.11807f
C3012 a_8431_5415# a_10132_5445# 0
C3013 a_12142_5459# a_10471_5727# 0
C3014 a_16539_5839# VDPWR 0.01025f
C3015 a_10888_5471# a_10525_5471# 0.00985f
C3016 a_9705_12861# a_10923_12931# 0.00148f
C3017 a_16657_22875# sky130_fd_sc_hd__dfxbp_1_3.Q_N 0.00244f
C3018 a_9556_17271# a_23133_17137# 0.38894f
C3019 a_5895_14763# a_4903_15345# 0
C3020 sky130_fd_sc_hd__inv_4_0.A a_18667_34839# 0
C3021 a_9779_13785# a_10675_14767# 0
C3022 a_14377_5833# a_14491_5723# 0
C3023 a_18625_4938# a_6238_6077# 0.10143f
C3024 a_5975_12927# a_6003_11935# 0
C3025 a_18693_31479# VDPWR 0.00348f
C3026 a_9379_14779# a_9779_13785# 0
C3027 a_9629_14779# a_9491_15377# 0
C3028 a_10975_23147# a_11406_23201# 0.10805f
C3029 uio_in[2] uio_in[1] 0.03102f
C3030 a_10385_4963# a_10160_4571# 0.00559f
C3031 a_18671_29731# sky130_fd_sc_hd__dfxbp_1_6.Q_N 0.12218f
C3032 a_12823_4553# VDPWR 0.18826f
C3033 a_6238_6077# a_14908_5833# 0.0019f
C3034 a_18667_34839# a_18667_34259# 0.10805f
C3035 a_6208_2817# a_14930_2159# 0
C3036 a_16660_2159# a_15119_1793# 0.03325f
C3037 a_18667_33636# VDPWR 0.31458f
C3038 a_11222_5837# a_6238_6077# 0
C3039 a_14940_22875# VDPWR 0
C3040 a_17733_4529# a_18625_5265# 0.00499f
C3041 a_8038_5023# a_6375_5299# 0.0035f
C3042 a_9493_12145# a_4915_10549# 0.00128f
C3043 a_6281_2043# a_8700_2159# 0
C3044 a_18693_24801# a_18667_24771# 0.0027f
C3045 a_9705_12861# a_9587_13813# 0
C3046 a_3199_1791# VDPWR 1.39907f
C3047 a_13284_5459# a_12533_5715# 0.00682f
C3048 VDPWR a_18667_25879# 0.21284f
C3049 a_9779_13785# a_10799_13773# 0
C3050 a_12793_14007# a_11979_13399# 0.00121f
C3051 a_17425_5473# a_16902_5473# 0
C3052 a_23677_14701# a_23731_14309# 0.09132f
C3053 a_4515_11543# a_4597_11543# 0.00641f
C3054 a_3990_1761# a_3938_1787# 0.1439f
C3055 a_18693_31299# a_18667_31684# 0.03733f
C3056 a_10289_4963# a_10160_4571# 0.00792f
C3057 a_18663_27017# a_18667_24771# 0
C3058 sky130_fd_sc_hd__dfxbp_1_4.Q_N a_17605_23241# 0
C3059 a_13161_23139# sky130_fd_sc_hd__dfxbp_1_3.Q_N 0
C3060 a_24234_14385# a_24407_14651# 0.00222f
C3061 a_17544_4895# a_6238_6077# 0
C3062 a_6208_2817# a_7944_1767# 0.00211f
C3063 a_16402_4529# VDPWR 0.18199f
C3064 a_14233_1793# a_13840_1767# 0.02283f
C3065 a_14596_1793# a_6208_2817# 0
C3066 sky130_fd_sc_hd__dfxbp_1_5.CLK sky130_fd_sc_hd__dfxbp_1_7.CLK 0
C3067 a_9715_11297# a_11147_11911# 0.00683f
C3068 a_6238_6077# a_10160_4571# 0
C3069 a_6629_15387# a_4503_16339# 0
C3070 a_18667_33636# sky130_fd_sc_hd__dfxbp_1_9.Q 0.01409f
C3071 a_14825_4547# VDPWR 0.18752f
C3072 a_6208_2817# a_10121_2159# 0
C3073 a_6375_5299# a_7315_5043# 0.13739f
C3074 a_10888_5837# a_12194_5433# 0
C3075 a_15431_5467# VDPWR 1.41244f
C3076 a_8377_5305# a_8794_5415# 0.06611f
C3077 a_10499_4853# a_10385_4597# 0
C3078 a_11439_4597# a_12769_4809# 0.21189f
C3079 a_24407_14651# a_24318_14385# 0
C3080 a_4839_12857# a_6021_13769# 0
C3081 a_18663_27120# sky130_fd_sc_hd__dfxbp_1_7.CLK 0
C3082 a_11406_23201# VDPWR 0.21318f
C3083 a_10235_2049# a_10986_2159# 0.00696f
C3084 a_8729_23143# sky130_fd_sc_hd__dfxbp_1_0.CLK 0
C3085 a_10357_5837# a_10471_5727# 0
C3086 a_9943_22879# a_10477_23245# 0.0027f
C3087 a_5942_1761# a_6208_2817# 0
C3088 a_13284_5459# a_6238_6077# 0
C3089 a_8377_5305# a_8263_5415# 0
C3090 a_17425_5473# a_18625_4938# 0.06919f
C3091 a_9715_11297# a_9771_12117# 0.25132f
C3092 a_5809_14763# a_4903_15345# 0.0039f
C3093 uio_out[4] uio_out[3] 0.03102f
C3094 a_14657_4547# a_14432_4521# 0.00487f
C3095 a_12113_1793# a_12227_2049# 0
C3096 a_9943_22879# a_8561_23241# 0
C3097 a_18667_33636# a_18667_31977# 0
C3098 a_17191_23241# a_17011_22875# 0.00123f
C3099 sky130_fd_sc_hd__dfxbp_1_7.Q a_18697_29053# 0
C3100 a_7863_22875# VDPWR 0.31414f
C3101 sky130_fd_sc_hd__inv_2_0.A a_18667_34470# 0.00379f
C3102 a_23511_14701# a_9556_17271# 0.04167f
C3103 a_9556_17271# sky130_fd_sc_hd__dfxbp_1_0.CLK 0.21701f
C3104 a_16243_2049# a_16129_1793# 0
C3105 a_11411_5471# a_12430_4527# 0
C3106 a_12039_15239# a_11583_15239# 0
C3107 a_13186_4553# a_11439_4597# 0.08907f
C3108 a_8377_5305# VDPWR 0.4515f
C3109 sky130_fd_sc_hd__dfxbp_1_1.Q_N a_12993_23237# 0
C3110 a_17210_4895# VDPWR 0.02205f
C3111 a_6208_2817# a_12655_4553# 0
C3112 a_9223_1793# a_10652_2159# 0.03325f
C3113 sky130_fd_sc_hd__dfxbp_1_6.Q_N sky130_fd_sc_hd__dfxbp_1_9.Q_N 0
C3114 a_6389_13769# a_4849_11293# 0.00488f
C3115 a_6389_13769# a_5851_13769# 0.07901f
C3116 a_9621_13111# a_9379_14779# 0
C3117 a_9713_14529# a_9369_16343# 0
C3118 a_7173_15235# a_4903_15345# 0
C3119 a_14657_4547# a_13709_4553# 0
C3120 a_11195_12931# a_11979_13399# 0
C3121 VDPWR a_8700_2159# 0.02101f
C3122 a_5975_12927# VDPWR 0.23989f
C3123 sky130_fd_sc_hd__dfxbp_1_5.Q_N a_18667_25510# 0.09273f
C3124 a_2706_5051# a_2217_5025# 0.08994f
C3125 a_11411_5471# a_12950_5459# 0.08907f
C3126 a_6429_5409# VDPWR 0.00968f
C3127 a_4839_12857# a_6329_12927# 0.08252f
C3128 a_9371_13111# a_9453_13111# 0.00641f
C3129 a_16583_4529# VDPWR 0.00129f
C3130 a_6021_13769# a_4837_16089# 0.00246f
C3131 a_22274_16171# VDPWR 0.4343f
C3132 a_9705_12861# a_9769_15349# 0.1369f
C3133 a_6717_15235# a_4837_16089# 0
C3134 a_9705_12861# VDPWR 1.04841f
C3135 a_9381_11547# a_9463_11547# 0.00641f
C3136 a_18671_29731# sky130_fd_sc_hd__dfxbp_1_7.Q_N 0
C3137 a_6238_6077# a_24152_14385# 0.01336f
C3138 a_11411_5471# a_12950_5825# 0.03325f
C3139 VDPWR a_4513_14775# 0.54082f
C3140 a_7113_13395# a_4915_10549# 0.2011f
C3141 a_10975_23147# a_10933_22879# 0
C3142 a_14233_1793# a_13969_1793# 0
C3143 a_10923_12931# VDPWR 0
C3144 a_24241_14651# a_24407_14651# 0.00988f
C3145 a_18667_24874# a_19059_24851# 0
C3146 a_18742_16187# a_17254_16187# 0
C3147 a_17096_23241# VDPWR 0.25533f
C3148 a_10717_13773# a_9501_13813# 0
C3149 a_6208_2817# a_12227_2049# 0.00304f
C3150 a_4763_14775# a_4513_14775# 0.02504f
C3151 a_17521_23241# a_17605_23241# 0.00851f
C3152 a_10499_4853# a_10553_4963# 0.03622f
C3153 VDPWR a_18667_33834# 0.19116f
C3154 a_12039_15239# a_9556_17271# 0.04708f
C3155 a_15407_23143# sky130_fd_sc_hd__dfxbp_1_2.Q_N 0
C3156 a_6208_2817# a_14771_4803# 0
C3157 a_8283_2049# a_8337_1793# 0.00386f
C3158 a_11411_5471# a_13473_5459# 0
C3159 a_8377_5305# a_10888_5471# 0
C3160 a_13167_1793# a_12644_1793# 0
C3161 a_13840_1767# a_14065_2159# 0.00559f
C3162 a_12615_14007# a_9556_17271# 0.10822f
C3163 sky130_fd_sc_hd__dfxbp_1_1.Q_N a_10891_23245# 0
C3164 a_9896_1767# a_10289_2159# 0.02301f
C3165 sky130_fd_sc_hd__dfxbp_1_7.Q a_18663_27017# 0
C3166 a_18663_28125# VDPWR 0.21336f
C3167 a_9587_13813# VDPWR 0.003f
C3168 a_6003_11935# VDPWR 0.22391f
C3169 a_14281_5467# a_13473_5459# 0
C3170 a_8283_2049# a_9844_1793# 0
C3171 a_11255_13773# a_9713_14529# 0
C3172 a_9631_11297# a_4915_10549# 0
C3173 a_16402_4529# a_16454_4503# 0.1439f
C3174 a_14179_2049# a_6208_2817# 0.00304f
C3175 a_14940_22875# a_14814_23241# 0.00553f
C3176 sky130_fd_sc_hd__dfxbp_1_9.Q a_18667_33834# 0
C3177 a_17733_4529# a_15711_4547# 0.00125f
C3178 VDPWR a_10933_22879# 0
C3179 a_6281_2043# VDPWR 0.45167f
C3180 sky130_fd_sc_hd__dfxbp_1_9.CLK a_18671_30311# 0.20774f
C3181 a_16454_4503# a_15431_5467# 0
C3182 a_17210_4529# a_16485_5729# 0
C3183 a_18667_25006# a_18693_24801# 0.00772f
C3184 a_16539_5473# VDPWR 0.18676f
C3185 a_6238_6077# a_10525_5471# 0
C3186 a_18667_32188# a_18667_31354# 0.19462f
C3187 a_14100_5467# a_14152_5441# 0.1439f
C3188 a_9223_1793# a_9844_1793# 0.0504f
C3189 a_4837_16089# a_4753_16089# 0.00234f
C3190 sky130_fd_sc_hd__dfxbp_1_2.CLK a_13119_22871# 0
C3191 a_10761_14767# a_9703_16093# 0
C3192 a_10975_23147# a_12483_22871# 0
C3193 a_2289_5307# a_2706_5417# 0.06611f
C3194 a_12736_22983# a_12483_22871# 0
C3195 a_6862_13645# a_4915_10549# 0
C3196 a_9781_10553# a_11728_13649# 0
C3197 a_18667_25006# a_18663_27017# 0
C3198 a_14908_5467# a_16146_5447# 0
C3199 a_14100_5467# a_12533_5715# 0
C3200 a_14545_5833# VDPWR 0.00865f
C3201 sky130_fd_sc_hd__dfxbp_1_1.Q_N a_10109_22879# 0.5114f
C3202 a_23761_14335# ui_in[1] 0.20361f
C3203 a_10975_23147# VDPWR 0.51295f
C3204 a_11810_13649# a_9705_12861# 0
C3205 a_9317_5049# a_15431_5467# 0.05142f
C3206 VDPWR a_12736_22983# 0.19095f
C3207 a_19063_29704# a_18671_29942# 0.00617f
C3208 a_12113_1793# a_6208_2817# 0
C3209 a_9556_17271# a_11979_13399# 0.0349f
C3210 a_16793_4785# a_15431_5467# 0
C3211 a_18671_29942# VDPWR 0.19977f
C3212 a_16297_2159# a_6208_2817# 0.00107f
C3213 a_6281_2043# a_6698_2153# 0.06611f
C3214 a_8794_5415# VDPWR 0.02122f
C3215 a_12129_22871# a_9943_22879# 0
C3216 a_12039_15239# a_9703_16093# 0.04213f
C3217 a_2289_5307# a_2217_5025# 0.25757f
C3218 a_2187_1765# a_5080_2153# 0
C3219 a_3010_2157# a_2187_1765# 0
C3220 a_24234_14385# ui_in[0] 0.28452f
C3221 a_15693_17123# VDPWR 0.41601f
C3222 a_8263_5415# VDPWR 0
C3223 a_14100_5467# a_6238_6077# 0.00306f
C3224 a_23677_14701# a_6238_6077# 0
C3225 a_8377_5305# a_9317_5049# 0.13758f
C3226 a_8645_23241# a_8304_22987# 0
C3227 a_9317_5049# a_17210_4895# 0
C3228 a_15407_23143# a_15365_22875# 0
C3229 a_14541_22875# a_16657_22875# 0
C3230 a_12615_14007# a_12697_14007# 0.00695f
C3231 sky130_fd_sc_hd__dfxbp_1_2.CLK a_12993_23237# 0
C3232 a_16297_2159# a_16033_2159# 0
C3233 a_16454_4503# a_16583_4529# 0.00758f
C3234 a_8561_23241# a_8729_23143# 0.31062f
C3235 a_19063_29704# VDPWR 0
C3236 VDPWR a_12483_22871# 0.07693f
C3237 a_15641_17149# sky130_fd_sc_hd__dfxbp_1_0.CLK 0.02419f
C3238 a_6238_6077# a_16539_5839# 0.00117f
C3239 a_10717_13773# a_11147_11911# 0
C3240 a_4849_11293# a_4597_11543# 0
C3241 a_4847_14525# a_4711_15373# 0
C3242 ui_in[0] a_24318_14385# 0.00255f
C3243 a_7944_1767# a_6335_1787# 0
C3244 a_12281_1793# VDPWR 0.18609f
C3245 a_16793_4785# a_17210_4895# 0.06611f
C3246 a_9769_15349# VDPWR 0.38134f
C3247 a_4119_2153# a_2187_1765# 0
C3248 a_4423_5299# VDPWR 0.45098f
C3249 a_6629_15387# a_4837_16089# 0.27498f
C3250 a_8167_5049# a_8431_5049# 0
C3251 VDPWR a_9034_2159# 0
C3252 a_7173_15235# a_7749_14003# 0.16707f
C3253 sky130_fd_sc_hd__dfxbp_1_0.Q_N sky130_fd_sc_hd__dfxbp_1_1.CLK 0.15244f
C3254 a_11979_13399# a_10841_12931# 0
C3255 a_13473_5459# a_14908_5833# 0.03325f
C3256 a_9160_23197# VDPWR 0.21267f
C3257 a_9369_16343# a_9491_15377# 0.00144f
C3258 a_5942_1761# a_6335_1787# 0.02283f
C3259 a_4763_14775# VDPWR 0.33336f
C3260 a_2259_2047# a_2676_2157# 0.06611f
C3261 a_4847_14525# a_4595_14775# 0
C3262 a_7697_22875# a_9943_22879# 0
C3263 a_17733_4529# a_18839_4938# 0
C3264 a_15119_1793# a_14930_2159# 0
C3265 a_8337_1793# a_8169_1793# 0
C3266 a_11406_23201# sky130_fd_sc_hd__dfxbp_1_2.Q_N 0
C3267 a_6792_5043# a_5363_5043# 0.08907f
C3268 a_14541_22875# a_13161_23139# 0
C3269 sky130_fd_sc_hd__dfxbp_1_9.Q VDPWR 0.27231f
C3270 a_5269_1787# a_6167_1787# 0
C3271 a_18663_28125# a_18671_29203# 0
C3272 a_6208_2817# a_16033_2159# 0
C3273 a_9703_16093# a_11979_13399# 0
C3274 a_18667_25510# sky130_fd_sc_hd__dfxbp_1_7.Q_N 0
C3275 a_12793_14007# a_11147_11911# 0.00264f
C3276 a_12697_14007# a_11979_13399# 0.00223f
C3277 a_16402_4529# a_6238_6077# 0
C3278 a_4849_11293# a_6021_13769# 0
C3279 a_6021_13769# a_5851_13769# 0.00167f
C3280 a_17210_4895# a_16847_4895# 0.00847f
C3281 a_12587_5459# a_10471_5727# 0
C3282 VDPWR a_6698_2153# 0.02101f
C3283 sky130_fd_sc_hd__dfxbp_1_4.CLK a_15838_23197# 0.20705f
C3284 a_14596_1793# a_15119_1793# 0
C3285 a_23731_14309# VDPWR 0.37479f
C3286 a_18667_31449# a_18667_31354# 0.96835f
C3287 a_7113_13395# a_4839_12857# 0.00446f
C3288 a_16243_2049# a_16297_1793# 0.00386f
C3289 a_6238_6077# a_15431_5467# 0.0069f
C3290 a_4329_2043# a_4383_2153# 0.03622f
C3291 a_9713_14529# a_9629_14529# 0.00206f
C3292 a_2313_1791# a_1920_1765# 0.02283f
C3293 a_18667_31977# VDPWR 0.51535f
C3294 a_18663_27545# a_19055_27518# 0
C3295 a_2676_2157# a_2313_2157# 0.00847f
C3296 a_4840_5043# a_2217_5025# 0
C3297 sky130_fd_sc_hd__dfxbp_1_0.Q_N a_10807_23245# 0
C3298 a_17236_5839# a_6238_6077# 0
C3299 sky130_fd_sc_hd__dfxbp_1_5.Q_N a_18689_26867# 0
C3300 a_4746_2153# a_4383_2153# 0.00847f
C3301 a_10888_5471# VDPWR 0.21774f
C3302 ui_in[0] a_24241_14651# 0.06316f
C3303 a_10235_2049# a_11888_1767# 0.00395f
C3304 a_18663_27017# a_18667_25299# 0
C3305 sky130_fd_sc_hd__dfxbp_1_5.CLK a_17096_23241# 0
C3306 a_18742_16187# a_18128_16189# 0.10376f
C3307 sky130_fd_sc_hd__dfxbp_1_1.Q_N a_10508_22879# 0.00188f
C3308 a_8687_22875# sky130_fd_sc_hd__dfxbp_1_0.Q_N 0.00125f
C3309 a_4753_16339# a_4503_16339# 0.02504f
C3310 a_18693_24621# sky130_fd_sc_hd__dfxbp_1_7.CLK 0
C3311 a_9705_12861# a_9715_11297# 0.82006f
C3312 a_11810_13649# VDPWR 0.0014f
C3313 sky130_fd_sc_hd__dfxbp_1_9.Q a_18667_31977# 0.12293f
C3314 a_16679_4895# VDPWR 0
C3315 a_8377_5305# a_6238_6077# 0.00302f
C3316 a_17210_4895# a_6238_6077# 0
C3317 sky130_fd_sc_hd__dfxbp_1_7.Q a_19055_27097# 0
C3318 a_2187_1765# a_4215_2153# 0
C3319 VDPWR a_3010_1791# 0
C3320 a_10923_12931# a_9715_11297# 0.00146f
C3321 a_4847_14525# a_4903_15345# 0.15229f
C3322 a_2706_5051# a_2343_5051# 0.00985f
C3323 a_4849_11293# a_6329_12927# 0.00976f
C3324 a_23761_14335# a_9556_17271# 0.00112f
C3325 a_6329_12927# a_5851_13769# 0
C3326 a_6281_2043# a_7032_1787# 0.00682f
C3327 a_18671_29942# a_18671_29203# 0.03218f
C3328 sky130_fd_sc_hd__dfxbp_1_2.CLK a_10109_22879# 0
C3329 a_14491_5723# a_14908_5833# 0.06611f
C3330 sky130_fd_sc_hd__dfxbp_1_1.Q_N a_10297_22879# 0.142f
C3331 a_6087_14735# a_4903_15345# 0
C3332 a_2259_2047# a_3938_1787# 0
C3333 a_6429_5409# a_6238_6077# 0
C3334 a_7113_13395# a_4837_16089# 0
C3335 a_6629_15387# sky130_fd_sc_hd__dfxbp_1_0.CLK 0.15686f
C3336 a_2145_2157# VDPWR 0
C3337 a_11195_12931# a_11147_11911# 0.00298f
C3338 a_18128_16189# a_17254_16187# 0.10446f
C3339 a_7173_15235# a_8193_13753# 0.04586f
C3340 a_11888_1767# a_11836_1793# 0.1439f
C3341 a_24234_14385# a_23133_17137# 0
C3342 a_17425_5473# a_15431_5467# 0
C3343 a_9381_11547# a_4915_10549# 0.00227f
C3344 VDPWR a_6071_1787# 0.00119f
C3345 a_8038_5023# a_6429_5043# 0
C3346 a_4839_12857# a_6862_13645# 0.00327f
C3347 a_17425_5473# a_17236_5839# 0
C3348 a_16454_4503# VDPWR 0.37087f
C3349 a_9943_22879# a_8304_22987# 0
C3350 a_7863_22875# a_8645_23241# 0
C3351 VDPWR a_5080_1787# 0
C3352 a_3229_5051# a_4309_5043# 0
C3353 VDPWR a_18671_29203# 0.66338f
C3354 a_1868_1791# VDPWR 0.17592f
C3355 a_11411_5471# a_12769_4809# 0
C3356 a_6208_2817# a_10553_4597# 0
C3357 a_18693_31893# a_18667_32188# 0.00851f
C3358 a_23677_14335# VDPWR 0
C3359 a_6717_15235# a_6635_15235# 0.00578f
C3360 a_18667_31684# a_18667_31354# 0.07715f
C3361 a_14152_5441# a_14545_5833# 0.02301f
C3362 a_15239_23241# a_16657_22875# 0
C3363 a_14814_23241# VDPWR 0.25536f
C3364 a_14729_22875# a_13161_23139# 0
C3365 a_9317_5049# VDPWR 2.56669f
C3366 a_14545_5833# a_12533_5715# 0
C3367 a_12295_22871# a_10807_23245# 0
C3368 a_16471_17161# sky130_fd_sc_hd__dfxbp_1_0.CLK 0.02548f
C3369 a_16793_4785# VDPWR 0.46736f
C3370 a_16486_16197# a_17254_16187# 0.1036f
C3371 a_18689_26867# a_18663_27252# 0.03733f
C3372 a_10975_23147# sky130_fd_sc_hd__dfxbp_1_2.Q_N 0
C3373 a_14375_22875# a_15838_23197# 0
C3374 a_10525_5837# a_10471_5727# 0.03622f
C3375 VDPWR a_7032_1787# 0
C3376 sky130_fd_sc_hd__dfxbp_1_2.Q_N a_12736_22983# 0.05782f
C3377 sky130_fd_sc_hd__dfxbp_1_8.Q_N a_18693_34175# 0
C3378 a_14179_2049# a_15119_1793# 0.13739f
C3379 a_4329_2043# a_4746_1787# 0.03016f
C3380 a_6805_15235# VDPWR 0.00152f
C3381 a_12823_4919# VDPWR 0.01321f
C3382 a_4837_16089# a_6862_13645# 0
C3383 a_14065_1793# VDPWR 0
C3384 a_16539_5473# a_6238_6077# 0
C3385 a_18667_24874# a_18667_24771# 0.14145f
C3386 sky130_fd_sc_hd__dfxbp_1_0.Q_N a_10550_22991# 0
C3387 a_9705_12861# a_10993_13773# 0.00253f
C3388 a_3990_1761# a_2187_1765# 0.00211f
C3389 a_6629_15387# a_4625_15373# 0
C3390 a_11175_1793# a_13167_1793# 0
C3391 a_6208_2817# a_9034_1793# 0
C3392 a_10499_4853# a_10471_5727# 0.00177f
C3393 a_6238_6077# a_14545_5833# 0.00115f
C3394 a_12295_22871# sky130_fd_sc_hd__dfxbp_1_3.CLK 0
C3395 a_7697_22875# a_8729_23143# 0.04808f
C3396 sky130_fd_sc_hd__dfxbp_1_5.Q_N a_18663_27252# 0
C3397 a_12823_4553# a_12430_4527# 0.02283f
C3398 a_24234_14385# sky130_fd_sc_hd__dfxbp_1_0.CLK 0.00519f
C3399 sky130_fd_sc_hd__dfxbp_1_5.CLK VDPWR 0.2879f
C3400 a_12823_4553# a_12559_4553# 0
C3401 a_23133_17137# a_24241_14651# 0
C3402 a_10025_1793# a_6208_2817# 0
C3403 VDPWR a_19235_17155# 0.45441f
C3404 a_18671_29438# sky130_fd_sc_hd__dfxbp_1_6.Q_N 0.04247f
C3405 a_13167_1793# a_13840_1767# 0.11878f
C3406 a_10160_4571# a_10385_4597# 0.00487f
C3407 a_14152_5441# VDPWR 0.33918f
C3408 a_7221_1787# a_8283_2049# 0.21187f
C3409 a_16094_5473# a_16275_5839# 0
C3410 a_18663_27756# sky130_fd_sc_hd__dfxbp_1_7.CLK 0
C3411 a_16454_4503# a_16679_4895# 0.00559f
C3412 a_2289_5307# a_2343_5051# 0.00386f
C3413 a_2187_1765# a_4383_1787# 0
C3414 a_16847_4895# VDPWR 0.01197f
C3415 sky130_fd_sc_hd__dfxbp_1_2.Q_N a_12483_22871# 0.142f
C3416 a_16371_5473# a_16485_5729# 0
C3417 a_9715_11297# a_9769_15349# 0.30637f
C3418 a_4213_5409# VDPWR 0
C3419 a_18663_27120# VDPWR 0.19118f
C3420 a_18667_33636# sky130_fd_sc_hd__dfxbp_1_8.Q_N 0.51145f
C3421 a_12533_5715# VDPWR 0.4413f
C3422 a_9715_11297# VDPWR 1.03424f
C3423 a_18693_33581# a_18667_33636# 0.0967f
C3424 a_9556_17271# a_11147_11911# 0.00289f
C3425 a_4755_12857# a_4505_13107# 0.00723f
C3426 a_10385_4963# VDPWR 0
C3427 a_17689_23143# a_18120_23197# 0.10805f
C3428 a_2175_5051# a_2343_5051# 0
C3429 sky130_fd_sc_hd__dfxbp_1_2.Q_N VDPWR 0.60665f
C3430 a_8794_5415# a_6238_6077# 0
C3431 a_12694_22871# a_12568_23237# 0.00553f
C3432 a_12017_1793# a_11175_1793# 0
C3433 a_6208_2817# a_6335_1787# 0
C3434 a_6238_6077# a_8263_5415# 0
C3435 a_14596_1793# a_14233_1793# 0.00985f
C3436 a_18667_32557# VDPWR 0.21288f
C3437 a_16297_2159# a_15119_1793# 0.04534f
C3438 a_11439_4597# a_10916_4597# 0
C3439 sky130_fd_sc_hd__dfxbp_1_2.CLK a_10508_22879# 0
C3440 a_9223_1793# a_7221_1787# 0
C3441 a_10121_2159# a_10289_2159# 0
C3442 a_14930_1793# VDPWR 0
C3443 a_14657_4547# a_14771_4803# 0
C3444 a_14100_5467# a_13473_5459# 0.05057f
C3445 sky130_fd_sc_hd__dfxbp_1_4.CLK a_17222_22875# 0
C3446 a_9371_13111# a_9379_14779# 0
C3447 a_18689_26867# sky130_fd_sc_hd__dfxbp_1_7.Q_N 0.142f
C3448 a_10289_4963# VDPWR 0
C3449 a_16793_4785# a_16679_4895# 0
C3450 sky130_fd_sc_hd__dfxbp_1_2.CLK a_10297_22879# 0
C3451 a_6238_6077# VDPWR 0.6644f
C3452 a_4839_12857# a_4913_13781# 0.44871f
C3453 a_6208_2817# a_10121_1793# 0
C3454 a_9943_22879# a_11406_23201# 0
C3455 sky130_fd_sc_hd__inv_16_0.A VDPWR 2.24965f
C3456 a_13520_4553# a_12769_4809# 0.00682f
C3457 sky130_fd_sc_hd__dfxbp_1_9.Q a_18667_32557# 0.20705f
C3458 a_12323_5825# a_12142_5459# 0
C3459 a_19063_29283# VDPWR 0
C3460 a_15323_23241# VDPWR 0.00628f
C3461 sky130_fd_sc_hd__dfxbp_1_5.Q_N sky130_fd_sc_hd__dfxbp_1_7.Q_N 0
C3462 a_18667_24874# a_19059_25272# 0
C3463 a_4032_5043# a_4084_5017# 0.1439f
C3464 a_9943_22879# a_7863_22875# 0
C3465 a_6629_15387# a_6635_15235# 0.1684f
C3466 a_9317_5049# a_16454_4503# 0
C3467 a_6389_13769# a_6281_11907# 0.00254f
C3468 a_11147_11911# a_10841_12931# 0
C3469 a_20384_16179# a_22274_16171# 0
C3470 a_3990_1761# a_4215_1787# 0.00487f
C3471 ena VGND 0.07038f
C3472 clk VGND 0.04288f
C3473 rst_n VGND 0.04288f
C3474 ui_in[2] VGND 0.04288f
C3475 ui_in[3] VGND 0.04288f
C3476 ui_in[4] VGND 0.04288f
C3477 ui_in[5] VGND 0.04288f
C3478 ui_in[6] VGND 0.04288f
C3479 ui_in[7] VGND 0.04288f
C3480 uio_in[0] VGND 0.04288f
C3481 uio_in[1] VGND 0.04288f
C3482 uio_in[2] VGND 0.04288f
C3483 uio_in[3] VGND 0.04288f
C3484 uio_in[4] VGND 0.04288f
C3485 uio_in[5] VGND 0.04288f
C3486 uio_in[6] VGND 0.04288f
C3487 uio_in[7] VGND 0.04288f
C3488 uo_out[1] VGND 0.04288f
C3489 uo_out[2] VGND 0.04276f
C3490 uo_out[3] VGND 0.04288f
C3491 uo_out[4] VGND 0.04288f
C3492 uo_out[5] VGND 0.04288f
C3493 uo_out[6] VGND 0.04288f
C3494 uo_out[7] VGND 0.04288f
C3495 uio_out[0] VGND 0.04288f
C3496 uio_out[1] VGND 0.04288f
C3497 uio_out[2] VGND 0.04288f
C3498 uio_out[3] VGND 0.04288f
C3499 uio_out[4] VGND 0.04288f
C3500 uio_out[5] VGND 0.04288f
C3501 uio_out[6] VGND 0.04288f
C3502 uio_out[7] VGND 0.04288f
C3503 uio_oe[0] VGND 0.04288f
C3504 uio_oe[1] VGND 0.04288f
C3505 uio_oe[2] VGND 0.04288f
C3506 uio_oe[3] VGND 0.04288f
C3507 uio_oe[4] VGND 0.04288f
C3508 uio_oe[5] VGND 0.04288f
C3509 uio_oe[6] VGND 0.04288f
C3510 uio_oe[7] VGND 0.07038f
C3511 ui_in[1] VGND 8.60028f
C3512 ui_in[0] VGND 9.30665f
C3513 uo_out[0] VGND 2.99304f
C3514 VDPWR VGND 0.27635p
C3515 a_16994_1793# VGND 0
C3516 a_16660_1793# VGND 0.01465f
C3517 a_16297_1793# VGND 0.02017f
C3518 a_16129_1793# VGND 0
C3519 a_16033_1793# VGND 0
C3520 a_14930_1793# VGND 0
C3521 a_14596_1793# VGND 0.01679f
C3522 a_14233_1793# VGND 0.02017f
C3523 a_14065_1793# VGND 0
C3524 a_13969_1793# VGND 0
C3525 a_16994_2159# VGND 0.00217f
C3526 a_16660_2159# VGND 0.1985f
C3527 a_16297_2159# VGND 0.21682f
C3528 a_16129_2159# VGND 0.00234f
C3529 a_16033_2159# VGND 0.00307f
C3530 a_15852_1793# VGND 0.16573f
C3531 a_12978_1793# VGND 0
C3532 a_12644_1793# VGND 0.01679f
C3533 a_12281_1793# VGND 0.02014f
C3534 a_12113_1793# VGND 0
C3535 a_12017_1793# VGND 0
C3536 a_14930_2159# VGND 0.00244f
C3537 a_14596_2159# VGND 0.20226f
C3538 a_14233_2159# VGND 0.21682f
C3539 a_14065_2159# VGND 0.00233f
C3540 a_13969_2159# VGND 0.00307f
C3541 a_13788_1793# VGND 0.16567f
C3542 a_10986_1793# VGND 0
C3543 a_10652_1793# VGND 0.01679f
C3544 a_10289_1793# VGND 0.02017f
C3545 a_10121_1793# VGND 0
C3546 a_10025_1793# VGND 0
C3547 a_12978_2159# VGND 0.00242f
C3548 a_12644_2159# VGND 0.20221f
C3549 a_12281_2159# VGND 0.21675f
C3550 a_12113_2159# VGND 0.00232f
C3551 a_12017_2159# VGND 0.00306f
C3552 a_11836_1793# VGND 0.16493f
C3553 a_9034_1793# VGND 0
C3554 a_8700_1793# VGND 0.01679f
C3555 a_8337_1793# VGND 0.02015f
C3556 a_8169_1793# VGND 0
C3557 a_8073_1793# VGND 0
C3558 a_10986_2159# VGND 0.00244f
C3559 a_10652_2159# VGND 0.20227f
C3560 a_10289_2159# VGND 0.21687f
C3561 a_10121_2159# VGND 0.00233f
C3562 a_10025_2159# VGND 0.00307f
C3563 a_9844_1793# VGND 0.16698f
C3564 a_7032_1787# VGND 0
C3565 a_6698_1787# VGND 0.01676f
C3566 a_6335_1787# VGND 0.02015f
C3567 a_6167_1787# VGND 0
C3568 a_6071_1787# VGND 0
C3569 a_9034_2159# VGND 0.00242f
C3570 a_8700_2159# VGND 0.20221f
C3571 a_8337_2159# VGND 0.21675f
C3572 a_8169_2159# VGND 0.00232f
C3573 a_8073_2159# VGND 0.00307f
C3574 a_7892_1793# VGND 0.16514f
C3575 a_5080_1787# VGND 0
C3576 a_4746_1787# VGND 0.01677f
C3577 a_4383_1787# VGND 0.02013f
C3578 a_4215_1787# VGND 0
C3579 a_4119_1787# VGND 0
C3580 a_7032_2153# VGND 0.00244f
C3581 a_6698_2153# VGND 0.20225f
C3582 a_6335_2153# VGND 0.21685f
C3583 a_6167_2153# VGND 0.00233f
C3584 a_6071_2153# VGND 0.00307f
C3585 a_5890_1787# VGND 0.16691f
C3586 a_3010_1791# VGND 0
C3587 a_2676_1791# VGND 0.01809f
C3588 a_2313_1791# VGND 0.01957f
C3589 a_2145_1791# VGND 0
C3590 a_2049_1791# VGND 0
C3591 a_5080_2153# VGND 0.00242f
C3592 a_4746_2153# VGND 0.20219f
C3593 a_4383_2153# VGND 0.21674f
C3594 a_4215_2153# VGND 0.00231f
C3595 a_4119_2153# VGND 0.00305f
C3596 a_3938_1787# VGND 0.16568f
C3597 a_16243_2049# VGND 1.4551f
C3598 a_15119_1793# VGND 1.29525f
C3599 a_15904_1767# VGND 0.53239f
C3600 a_14179_2049# VGND 1.46693f
C3601 a_13167_1793# VGND 1.24789f
C3602 a_13840_1767# VGND 0.53177f
C3603 a_12227_2049# VGND 1.4658f
C3604 a_11175_1793# VGND 1.26755f
C3605 a_11888_1767# VGND 0.53189f
C3606 a_10235_2049# VGND 1.46646f
C3607 a_9223_1793# VGND 1.24885f
C3608 a_9896_1767# VGND 0.53181f
C3609 a_8283_2049# VGND 1.46581f
C3610 a_7221_1787# VGND 1.27256f
C3611 a_7944_1767# VGND 0.53242f
C3612 a_6281_2043# VGND 1.46581f
C3613 a_5269_1787# VGND 1.24712f
C3614 a_5942_1761# VGND 0.53131f
C3615 a_4329_2043# VGND 1.46563f
C3616 a_3990_1761# VGND 0.53241f
C3617 a_3199_1791# VGND 1.30753f
C3618 a_3010_2157# VGND 0.00242f
C3619 a_2676_2157# VGND 0.20474f
C3620 a_2313_2157# VGND 0.21441f
C3621 a_2145_2157# VGND 0.0024f
C3622 a_2049_2157# VGND 0.00311f
C3623 a_1868_1791# VGND 0.17891f
C3624 a_2259_2047# VGND 1.46655f
C3625 a_1920_1765# VGND 0.54374f
C3626 a_2187_1765# VGND 3.3825f
C3627 a_17544_4529# VGND 0
C3628 a_17210_4529# VGND 0.01738f
C3629 a_16847_4529# VGND 0.01904f
C3630 a_18839_4938# VGND 0
C3631 a_18553_4938# VGND 0
C3632 a_15522_4547# VGND 0
C3633 a_15188_4547# VGND 0.01467f
C3634 a_14825_4547# VGND 0.02052f
C3635 a_14657_4547# VGND 0
C3636 a_14561_4547# VGND 0
C3637 a_17544_4895# VGND 0.00238f
C3638 a_17210_4895# VGND 0.20252f
C3639 a_16847_4895# VGND 0.21482f
C3640 a_16679_4895# VGND 0.00207f
C3641 a_16583_4895# VGND 0.0029f
C3642 a_16402_4529# VGND 0.15964f
C3643 a_16793_4785# VGND 1.46253f
C3644 a_16454_4503# VGND 0.51961f
C3645 a_15711_4547# VGND 1.22622f
C3646 a_13520_4553# VGND 0
C3647 a_13186_4553# VGND 0.01746f
C3648 a_12823_4553# VGND 0.01889f
C3649 a_15522_4913# VGND 0.00221f
C3650 a_15188_4913# VGND 0.19864f
C3651 a_14825_4913# VGND 0.21708f
C3652 a_14657_4913# VGND 0.00233f
C3653 a_14561_4913# VGND 0.00306f
C3654 a_14380_4547# VGND 0.16642f
C3655 a_14771_4803# VGND 1.45148f
C3656 a_14432_4521# VGND 0.53271f
C3657 a_13709_4553# VGND 1.23412f
C3658 a_11250_4597# VGND 0
C3659 a_10916_4597# VGND 0.01491f
C3660 a_10553_4597# VGND 0.01744f
C3661 a_10385_4597# VGND 0
C3662 a_10289_4597# VGND 0
C3663 a_13520_4919# VGND 0.00245f
C3664 a_13186_4919# VGND 0.20276f
C3665 a_12823_4919# VGND 0.21461f
C3666 a_12655_4919# VGND 0.00207f
C3667 a_12559_4919# VGND 0.0029f
C3668 a_12378_4553# VGND 0.16122f
C3669 a_12769_4809# VGND 1.46444f
C3670 a_12430_4527# VGND 0.52093f
C3671 a_11439_4597# VGND 1.30826f
C3672 a_11250_4963# VGND 0.00219f
C3673 a_10916_4963# VGND 0.19899f
C3674 a_10553_4963# VGND 0.21131f
C3675 a_10385_4963# VGND 0.00223f
C3676 a_10289_4963# VGND 0.00325f
C3677 a_10108_4597# VGND 0.18458f
C3678 a_10499_4853# VGND 1.43743f
C3679 a_10160_4571# VGND 0.54628f
C3680 a_9128_5049# VGND 0
C3681 a_8794_5049# VGND 0.01792f
C3682 a_8431_5049# VGND 0.02049f
C3683 a_8263_5049# VGND 0
C3684 a_8167_5049# VGND 0
C3685 a_18846_5265# VGND 0.00346f
C3686 a_18625_5265# VGND 0.00367f
C3687 a_18625_4938# VGND 0.31023f
C3688 a_17733_4529# VGND 0.64799f
C3689 a_18371_4938# VGND 0.36105f
C3690 a_17236_5473# VGND 0
C3691 a_16902_5473# VGND 0.02117f
C3692 a_16539_5473# VGND 0.0211f
C3693 a_16371_5473# VGND 0
C3694 a_16275_5473# VGND 0
C3695 a_17425_5473# VGND 1.04201f
C3696 a_15242_5467# VGND 0
C3697 a_14908_5467# VGND 0.01858f
C3698 a_14545_5467# VGND 0.02292f
C3699 a_14377_5467# VGND 0
C3700 a_14281_5467# VGND 0
C3701 a_17236_5839# VGND 0.00267f
C3702 a_16902_5839# VGND 0.20496f
C3703 a_16539_5839# VGND 0.21767f
C3704 a_16371_5839# VGND 0.00238f
C3705 a_16275_5839# VGND 0.0031f
C3706 a_16094_5473# VGND 0.16598f
C3707 a_13284_5459# VGND 0
C3708 a_12950_5459# VGND 0.02272f
C3709 a_12587_5459# VGND 0.02074f
C3710 a_12419_5459# VGND 0
C3711 a_12323_5459# VGND 0
C3712 a_15242_5833# VGND 0.00246f
C3713 a_14908_5833# VGND 0.20339f
C3714 a_14545_5833# VGND 0.21882f
C3715 a_14377_5833# VGND 0.00261f
C3716 a_14281_5833# VGND 0.00325f
C3717 a_14100_5467# VGND 0.17708f
C3718 a_11222_5471# VGND 0
C3719 a_10888_5471# VGND 0.10793f
C3720 a_10525_5471# VGND 0.10701f
C3721 a_10357_5471# VGND 0
C3722 a_10261_5471# VGND 0
C3723 a_13284_5825# VGND 0.00274f
C3724 a_12950_5825# VGND 0.20604f
C3725 a_12587_5825# VGND 0.21777f
C3726 a_12419_5825# VGND 0.00238f
C3727 a_12323_5825# VGND 0.00309f
C3728 a_12142_5459# VGND 0.16514f
C3729 a_16485_5729# VGND 1.49806f
C3730 a_15431_5467# VGND 1.22901f
C3731 a_16146_5447# VGND 0.53461f
C3732 a_14491_5723# VGND 1.47304f
C3733 a_13473_5459# VGND 1.27472f
C3734 a_14152_5441# VGND 0.55159f
C3735 a_12533_5715# VGND 1.49499f
C3736 a_12194_5433# VGND 0.53402f
C3737 a_11411_5471# VGND 1.25994f
C3738 a_9317_5049# VGND 4.0005f
C3739 a_7126_5043# VGND 0
C3740 a_6792_5043# VGND 0.01675f
C3741 a_6429_5043# VGND 0.02015f
C3742 a_6261_5043# VGND 0
C3743 a_6165_5043# VGND 0
C3744 a_9128_5415# VGND 0.00245f
C3745 a_8794_5415# VGND 0.20264f
C3746 a_8431_5415# VGND 0.21692f
C3747 a_8263_5415# VGND 0.00232f
C3748 a_8167_5415# VGND 0.00307f
C3749 a_7986_5049# VGND 0.164f
C3750 a_5174_5043# VGND 0
C3751 a_4840_5043# VGND 0.01675f
C3752 a_4477_5043# VGND 0.02018f
C3753 a_4309_5043# VGND 0
C3754 a_4213_5043# VGND 0
C3755 a_7126_5409# VGND 0.00244f
C3756 a_6792_5409# VGND 0.20224f
C3757 a_6429_5409# VGND 0.21685f
C3758 a_6261_5409# VGND 0.00234f
C3759 a_6165_5409# VGND 0.00308f
C3760 a_5984_5043# VGND 0.16327f
C3761 a_3040_5051# VGND 0
C3762 a_2706_5051# VGND 0.01704f
C3763 a_2343_5051# VGND 0.02075f
C3764 a_2175_5051# VGND 0
C3765 a_2079_5051# VGND 0
C3766 a_5174_5409# VGND 0.00247f
C3767 a_4840_5409# VGND 0.20252f
C3768 a_4477_5409# VGND 0.21723f
C3769 a_4309_5409# VGND 0.00233f
C3770 a_4213_5409# VGND 0.00308f
C3771 a_4032_5043# VGND 0.16632f
C3772 a_8377_5305# VGND 1.4752f
C3773 a_7315_5043# VGND 1.27412f
C3774 a_8038_5023# VGND 0.53252f
C3775 a_6375_5299# VGND 1.466f
C3776 a_5363_5043# VGND 1.24671f
C3777 a_6036_5017# VGND 0.53163f
C3778 a_4423_5299# VGND 1.4669f
C3779 a_4084_5017# VGND 0.53343f
C3780 a_3229_5051# VGND 1.3407f
C3781 a_3040_5417# VGND 0.00243f
C3782 a_2706_5417# VGND 0.20241f
C3783 a_2343_5417# VGND 0.21713f
C3784 a_2175_5417# VGND 0.0024f
C3785 a_2079_5417# VGND 0.00311f
C3786 a_1898_5051# VGND 0.17876f
C3787 a_2289_5307# VGND 1.46706f
C3788 a_1950_5025# VGND 0.54359f
C3789 a_11222_5837# VGND 0.00261f
C3790 a_10888_5837# VGND 0.23876f
C3791 a_10525_5837# VGND 0.27025f
C3792 a_10357_5837# VGND 0.00294f
C3793 a_10261_5837# VGND 0.00346f
C3794 a_10080_5471# VGND 0.20604f
C3795 a_10471_5727# VGND 1.73088f
C3796 a_10132_5445# VGND 0.65125f
C3797 a_2217_5025# VGND 3.40505f
C3798 a_9589_10581# VGND 0.00699f
C3799 a_4723_10577# VGND 0.00697f
C3800 a_9503_10581# VGND 0.4195f
C3801 a_4637_10577# VGND 0.41935f
C3802 a_9631_11297# VGND 0.00834f
C3803 a_4765_11293# VGND 0.00834f
C3804 a_9631_11547# VGND 0.02839f
C3805 a_9463_11547# VGND 0.00172f
C3806 a_4765_11543# VGND 0.02839f
C3807 a_4597_11543# VGND 0.00172f
C3808 a_9381_11547# VGND 0.51561f
C3809 a_4515_11543# VGND 0.51559f
C3810 a_10955_11939# VGND 0.00568f
C3811 a_6089_11935# VGND 0.00568f
C3812 a_9579_12145# VGND 0.00662f
C3813 a_10869_11939# VGND 0.30868f
C3814 a_9771_12117# VGND 0.97249f
C3815 a_4713_12141# VGND 0.00662f
C3816 a_6003_11935# VGND 0.30868f
C3817 a_4905_12113# VGND 0.97739f
C3818 a_9493_12145# VGND 0.41373f
C3819 a_4627_12141# VGND 0.4141f
C3820 a_10995_12931# VGND 0.00306f
C3821 a_10923_12931# VGND 0.00325f
C3822 a_9621_12861# VGND 0.00847f
C3823 a_6129_12927# VGND 0.00306f
C3824 a_6057_12927# VGND 0.00325f
C3825 a_4755_12857# VGND 0.00847f
C3826 a_9621_13111# VGND 0.02681f
C3827 a_9453_13111# VGND 0.00171f
C3828 a_9371_13111# VGND 0.51196f
C3829 a_10841_12931# VGND 0.30847f
C3830 a_4755_13107# VGND 0.02681f
C3831 a_4587_13107# VGND 0.00171f
C3832 a_4505_13107# VGND 0.51196f
C3833 a_5975_12927# VGND 0.30847f
C3834 a_11810_13649# VGND 0
C3835 a_11195_12931# VGND 0.65373f
C3836 a_11728_13649# VGND 0.28668f
C3837 a_10993_13773# VGND 0.00417f
C3838 a_10887_13773# VGND 0.00482f
C3839 a_10799_13773# VGND 0.00392f
C3840 a_9587_13813# VGND 0.00661f
C3841 a_12865_14007# VGND 0
C3842 a_12793_14007# VGND 0
C3843 a_12697_14007# VGND 0
C3844 a_11979_13399# VGND 0.70622f
C3845 a_11147_11911# VGND 1.75062f
C3846 a_9781_10553# VGND 4.41904f
C3847 a_12615_14007# VGND 0.39608f
C3848 a_11255_13773# VGND 0.58041f
C3849 a_10717_13773# VGND 0.32933f
C3850 a_9779_13785# VGND 1.18115f
C3851 a_6944_13645# VGND 0
C3852 a_6329_12927# VGND 0.65373f
C3853 a_6862_13645# VGND 0.28669f
C3854 a_6127_13769# VGND 0.00417f
C3855 a_6021_13769# VGND 0.00482f
C3856 a_5933_13769# VGND 0.00392f
C3857 a_4721_13809# VGND 0.00661f
C3858 a_7999_14003# VGND 0
C3859 a_7927_14003# VGND 0
C3860 a_7831_14003# VGND 0
C3861 a_7113_13395# VGND 0.70818f
C3862 a_6281_11907# VGND 1.7509f
C3863 a_4915_10549# VGND 4.31319f
C3864 a_7749_14003# VGND 0.39642f
C3865 a_6389_13769# VGND 0.58024f
C3866 a_9501_13813# VGND 0.41423f
C3867 a_5851_13769# VGND 0.32933f
C3868 a_4913_13781# VGND 1.18582f
C3869 a_4635_13809# VGND 0.41597f
C3870 a_24318_14385# VGND 0.11977f
C3871 a_24152_14385# VGND 0.24785f
C3872 a_23677_14335# VGND 0.00194f
C3873 a_23511_14335# VGND 0.27853f
C3874 a_24962_14701# VGND 0.35152f
C3875 a_24774_14701# VGND 0.27668f
C3876 a_24234_14385# VGND 0.09185f
C3877 a_24241_14651# VGND 0.00666f
C3878 a_6208_2817# VGND 12.6203f
C3879 a_6238_6077# VGND 12.5721f
C3880 a_23761_14335# VGND 0.50894f
C3881 a_9629_14529# VGND 0.00834f
C3882 a_4763_14525# VGND 0.00834f
C3883 a_23731_14309# VGND 0.45978f
C3884 a_23677_14701# VGND 0.00793f
C3885 a_23511_14701# VGND 0.03002f
C3886 a_10761_14767# VGND 0.00618f
C3887 a_9629_14779# VGND 0.02779f
C3888 a_9461_14779# VGND 0.00172f
C3889 a_5895_14763# VGND 0.00618f
C3890 a_9379_14779# VGND 0.51319f
C3891 a_9705_12861# VGND 2.64035f
C3892 a_9715_11297# VGND 3.44639f
C3893 a_4763_14775# VGND 0.02779f
C3894 a_4595_14775# VGND 0.00172f
C3895 a_4513_14775# VGND 0.51319f
C3896 a_4839_12857# VGND 2.6442f
C3897 a_4849_11293# VGND 3.44771f
C3898 a_10675_14767# VGND 0.29854f
C3899 a_5809_14763# VGND 0.29858f
C3900 a_11777_15239# VGND 0.00384f
C3901 a_11671_15239# VGND 0.00334f
C3902 a_11583_15239# VGND 0.00151f
C3903 a_12039_15239# VGND 1.2343f
C3904 a_6911_15235# VGND 0.00384f
C3905 a_6805_15235# VGND 0.00334f
C3906 a_6717_15235# VGND 0.00151f
C3907 a_9577_15377# VGND 0.00661f
C3908 a_11501_15239# VGND 0.30157f
C3909 a_10953_14739# VGND 0.68859f
C3910 a_9713_14529# VGND 1.05198f
C3911 a_8193_13753# VGND 3.07271f
C3912 a_9769_15349# VGND 1.66994f
C3913 a_7173_15235# VGND 1.23231f
C3914 a_4711_15373# VGND 0.00661f
C3915 a_6635_15235# VGND 0.30157f
C3916 a_6087_14735# VGND 0.68424f
C3917 a_4847_14525# VGND 1.05927f
C3918 a_4903_15345# VGND 1.67323f
C3919 a_9491_15377# VGND 0.41662f
C3920 a_4625_15373# VGND 0.41665f
C3921 a_9619_16093# VGND 0.00773f
C3922 a_4753_16089# VGND 0.00773f
C3923 a_22274_16171# VGND 0.7476f
C3924 a_21506_16181# VGND 0.67384f
C3925 a_20384_16179# VGND 0.81524f
C3926 a_19510_16177# VGND 0.73239f
C3927 a_18742_16187# VGND 0.66246f
C3928 a_18128_16189# VGND 0.60419f
C3929 a_17254_16187# VGND 0.73256f
C3930 a_16486_16197# VGND 0.67981f
C3931 a_9703_16093# VGND 2.28792f
C3932 a_9619_16343# VGND 0.01843f
C3933 a_9451_16343# VGND 0.00117f
C3934 a_4837_16089# VGND 2.39375f
C3935 a_4753_16339# VGND 0.01843f
C3936 a_4585_16339# VGND 0.00117f
C3937 a_9369_16343# VGND 0.50464f
C3938 a_4503_16339# VGND 0.50495f
C3939 a_23133_17137# VGND 2.24042f
C3940 a_22365_17147# VGND 0.66623f
C3941 a_21491_17145# VGND 0.71701f
C3942 a_20877_17147# VGND 0.58889f
C3943 a_20109_17157# VGND 0.64571f
C3944 a_19235_17155# VGND 0.71158f
C3945 a_18113_17153# VGND 0.78148f
C3946 a_15641_17149# VGND 1.60765f
C3947 a_15693_17123# VGND 0.65426f
C3948 a_17345_17163# VGND 0.65615f
C3949 a_16471_17161# VGND 0.71929f
C3950 a_6629_15387# VGND 2.67988f
C3951 a_9556_17271# VGND 8.73856f
C3952 a_17647_22875# VGND 0.0058f
C3953 a_17222_22875# VGND 0.00795f
C3954 a_17605_23241# VGND 0
C3955 a_15365_22875# VGND 0.0058f
C3956 a_17191_23241# VGND 0
C3957 a_17011_22875# VGND 0.06664f
C3958 a_18120_23197# VGND 0.21543f
C3959 a_17521_23241# VGND 0.30409f
C3960 a_17689_23143# VGND 0.5725f
C3961 a_17096_23241# VGND 0.22722f
C3962 a_17264_22987# VGND 0.27139f
C3963 a_16823_22875# VGND 0.36748f
C3964 sky130_fd_sc_hd__dfxbp_1_4.Q_N VGND 0.69666f
C3965 a_16657_22875# VGND 0.57488f
C3966 sky130_fd_sc_hd__dfxbp_1_4.CLK VGND 0.80935f
C3967 a_14940_22875# VGND 0.00795f
C3968 a_15323_23241# VGND 0
C3969 a_13119_22871# VGND 0.00581f
C3970 a_14909_23241# VGND 0
C3971 a_14729_22875# VGND 0.06662f
C3972 a_15838_23197# VGND 0.20853f
C3973 a_15239_23241# VGND 0.30353f
C3974 a_15407_23143# VGND 0.56668f
C3975 a_14814_23241# VGND 0.22701f
C3976 a_14982_22987# VGND 0.27091f
C3977 a_14541_22875# VGND 0.3673f
C3978 sky130_fd_sc_hd__dfxbp_1_3.Q_N VGND 0.68547f
C3979 a_14375_22875# VGND 0.57353f
C3980 sky130_fd_sc_hd__dfxbp_1_3.CLK VGND 0.7916f
C3981 a_12694_22871# VGND 0.00797f
C3982 a_13077_23237# VGND 0
C3983 a_10933_22879# VGND 0.0058f
C3984 a_12663_23237# VGND 0
C3985 a_12483_22871# VGND 0.0667f
C3986 a_13592_23193# VGND 0.20847f
C3987 a_12993_23237# VGND 0.30357f
C3988 a_13161_23139# VGND 0.56662f
C3989 a_12568_23237# VGND 0.22707f
C3990 a_12736_22983# VGND 0.27094f
C3991 a_12295_22871# VGND 0.36728f
C3992 sky130_fd_sc_hd__dfxbp_1_2.Q_N VGND 0.68341f
C3993 a_12129_22871# VGND 0.57209f
C3994 sky130_fd_sc_hd__dfxbp_1_2.CLK VGND 0.7582f
C3995 a_10508_22879# VGND 0.00795f
C3996 a_10891_23245# VGND 0
C3997 a_8687_22875# VGND 0.0058f
C3998 a_10477_23245# VGND 0
C3999 a_10297_22879# VGND 0.06662f
C4000 a_11406_23201# VGND 0.20801f
C4001 a_10807_23245# VGND 0.30353f
C4002 a_10975_23147# VGND 0.56628f
C4003 a_10382_23245# VGND 0.22725f
C4004 a_10550_22991# VGND 0.27152f
C4005 a_10109_22879# VGND 0.36737f
C4006 sky130_fd_sc_hd__dfxbp_1_1.Q_N VGND 0.68225f
C4007 a_9943_22879# VGND 0.57365f
C4008 sky130_fd_sc_hd__dfxbp_1_1.CLK VGND 0.79274f
C4009 a_8262_22875# VGND 0.00795f
C4010 a_8645_23241# VGND 0
C4011 a_8231_23241# VGND 0
C4012 a_8051_22875# VGND 0.06662f
C4013 a_9160_23197# VGND 0.20845f
C4014 a_8561_23241# VGND 0.30354f
C4015 a_8729_23143# VGND 0.56658f
C4016 a_8136_23241# VGND 0.22701f
C4017 a_8304_22987# VGND 0.27092f
C4018 a_7863_22875# VGND 0.36871f
C4019 sky130_fd_sc_hd__dfxbp_1_0.Q_N VGND 0.68697f
C4020 a_7697_22875# VGND 0.59268f
C4021 sky130_fd_sc_hd__dfxbp_1_0.CLK VGND 15.6228f
C4022 sky130_fd_sc_hd__dfxbp_1_5.CLK VGND 1.40037f
C4023 a_18693_24621# VGND 0.06771f
C4024 a_19059_24851# VGND 0.00818f
C4025 a_18693_24801# VGND 0
C4026 a_18667_25006# VGND 0.22823f
C4027 a_18667_24874# VGND 0.272f
C4028 a_18667_24771# VGND 0.59552f
C4029 a_18667_24676# VGND 0.37151f
C4030 a_19059_25272# VGND 0.0058f
C4031 a_18693_25215# VGND 0
C4032 a_18667_25510# VGND 0.30735f
C4033 a_18667_25299# VGND 0.57527f
C4034 a_18667_25879# VGND 0.21106f
C4035 sky130_fd_sc_hd__dfxbp_1_5.Q_N VGND 0.69959f
C4036 sky130_fd_sc_hd__dfxbp_1_7.CLK VGND 0.81119f
C4037 a_18689_26867# VGND 0.0677f
C4038 a_19055_27097# VGND 0.00818f
C4039 a_18689_27047# VGND 0
C4040 a_18663_27252# VGND 0.22823f
C4041 a_18663_27120# VGND 0.27203f
C4042 a_18663_27017# VGND 0.57798f
C4043 a_18663_26922# VGND 0.37066f
C4044 a_19055_27518# VGND 0.0058f
C4045 a_18689_27461# VGND 0
C4046 a_18663_27756# VGND 0.30733f
C4047 a_18663_27545# VGND 0.57466f
C4048 a_18663_28125# VGND 0.21057f
C4049 sky130_fd_sc_hd__dfxbp_1_7.Q_N VGND 0.6935f
C4050 sky130_fd_sc_hd__dfxbp_1_7.Q VGND 0.77403f
C4051 a_18697_29053# VGND 0.0678f
C4052 a_19063_29283# VGND 0.00821f
C4053 a_18697_29233# VGND 0
C4054 a_18671_29438# VGND 0.2283f
C4055 a_18671_29306# VGND 0.27203f
C4056 a_18671_29203# VGND 0.57659f
C4057 a_18671_29108# VGND 0.37072f
C4058 a_19063_29704# VGND 0.00581f
C4059 a_18697_29647# VGND 0
C4060 a_18671_29942# VGND 0.30737f
C4061 a_18671_29731# VGND 0.5752f
C4062 a_18671_30311# VGND 0.2111f
C4063 sky130_fd_sc_hd__dfxbp_1_6.Q_N VGND 0.69535f
C4064 sky130_fd_sc_hd__dfxbp_1_9.CLK VGND 0.80969f
C4065 a_18693_31299# VGND 0.06771f
C4066 a_19059_31529# VGND 0.00818f
C4067 a_18693_31479# VGND 0
C4068 a_18667_31684# VGND 0.22823f
C4069 a_18667_31552# VGND 0.27199f
C4070 a_18667_31449# VGND 0.57799f
C4071 a_18667_31354# VGND 0.37071f
C4072 a_19059_31950# VGND 0.0058f
C4073 a_18693_31893# VGND 0
C4074 a_18667_32188# VGND 0.30733f
C4075 a_18667_31977# VGND 0.57493f
C4076 a_18667_32557# VGND 0.21114f
C4077 sky130_fd_sc_hd__dfxbp_1_9.Q_N VGND 0.69698f
C4078 sky130_fd_sc_hd__dfxbp_1_9.Q VGND 0.82658f
C4079 a_18693_33581# VGND 0.06772f
C4080 a_19059_33811# VGND 0.00818f
C4081 a_18693_33761# VGND 0
C4082 a_18667_33966# VGND 0.22825f
C4083 a_18667_33834# VGND 0.27203f
C4084 a_18667_33731# VGND 0.58026f
C4085 a_18667_33636# VGND 0.37078f
C4086 a_19059_34232# VGND 0.0058f
C4087 a_18693_34175# VGND 0
C4088 a_18667_34470# VGND 0.30738f
C4089 a_18667_34259# VGND 0.57832f
C4090 a_18667_34839# VGND 0.21444f
C4091 sky130_fd_sc_hd__dfxbp_1_8.Q_N VGND 0.70564f
C4092 sky130_fd_sc_hd__inv_2_0.A VGND 1.24888f
C4093 sky130_fd_sc_hd__inv_4_0.A VGND 1.01027f
C4094 sky130_fd_sc_hd__inv_6_0.A VGND 1.44919f
C4095 sky130_fd_sc_hd__inv_8_0.A VGND 1.65411f
C4096 sky130_fd_sc_hd__inv_12_0.A VGND 2.41535f
C4097 sky130_fd_sc_hd__inv_16_0.A VGND 3.17596f
.ends

