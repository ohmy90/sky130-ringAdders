magic
tech sky130A
magscale 1 2
timestamp 1755029384
<< nwell >>
rect 18428 33348 18749 35264
rect 18436 31042 18757 32958
rect 18444 28828 18765 30744
rect 18426 26628 18747 28544
rect 18434 24414 18755 26330
rect 7508 23105 9424 23426
rect 9722 23113 11638 23434
rect 11922 23095 13838 23416
rect 14136 23103 16052 23424
rect 16442 23111 18358 23432
rect 15443 17064 15881 17385
rect 16229 17102 16659 17423
rect 17095 17104 17533 17425
rect 17873 17094 18301 17415
rect 18989 17096 19423 17417
rect 19855 17098 20297 17419
rect 20625 17088 21065 17409
rect 21327 17086 21771 17407
rect 22111 17088 22553 17409
rect 22969 17078 23411 17399
rect 9296 16307 10016 16628
rect 9394 15563 9930 15884
rect 11436 15453 12156 15774
rect 9306 14743 10026 15064
rect 10578 14953 11114 15274
rect 9404 13999 9940 14320
rect 10652 13987 11372 14308
rect 12550 13971 13178 14292
rect 11622 13613 12158 13934
rect 9298 13075 10018 13396
rect 10776 13145 11312 13466
rect 9396 12331 9932 12652
rect 10772 12125 11308 12446
rect 9308 11511 10028 11832
rect 9406 10767 9942 11088
rect 6074 6018 6426 6339
rect 9980 5386 11528 5707
rect 12042 5374 13588 5695
rect 14000 5382 15546 5703
rect 15994 5388 17542 5709
rect 1798 4966 3346 5287
rect 3932 4958 5480 5279
rect 5884 4958 7432 5279
rect 7886 4964 9434 5285
rect 10008 4512 11556 4833
rect 12278 4468 13826 4789
rect 14280 4462 15828 4783
rect 16302 4444 17850 4765
rect 1768 1706 3316 2027
rect 3838 1702 5386 2023
rect 5790 1702 7338 2023
rect 7792 1708 9340 2029
rect 9744 1708 11292 2029
rect 11736 1708 13284 2029
rect 13688 1708 15236 2029
rect 15752 1708 17300 2029
<< pwell >>
rect 18815 35137 18972 35223
rect 18807 34580 18989 35133
rect 18853 34272 18989 34580
rect 18809 34090 18989 34272
rect 18853 33449 18989 34090
rect 18853 33415 19027 33449
rect 18853 33387 18989 33415
rect 18823 32831 18980 32917
rect 18815 32274 18997 32827
rect 18861 31966 18997 32274
rect 18817 31784 18997 31966
rect 18861 31143 18997 31784
rect 18861 31109 19035 31143
rect 18861 31081 18997 31109
rect 18831 30617 18988 30703
rect 18823 30060 19005 30613
rect 18869 29752 19005 30060
rect 18825 29570 19005 29752
rect 18869 28929 19005 29570
rect 18869 28895 19043 28929
rect 18869 28867 19005 28895
rect 18813 28417 18970 28503
rect 18805 27860 18987 28413
rect 18851 27552 18987 27860
rect 18807 27370 18987 27552
rect 18851 26729 18987 27370
rect 18851 26695 19025 26729
rect 18851 26667 18987 26695
rect 18821 26203 18978 26289
rect 18813 25646 18995 26199
rect 18859 25338 18995 25646
rect 18815 25156 18995 25338
rect 18859 24515 18995 25156
rect 18859 24481 19033 24515
rect 18859 24453 18995 24481
rect 8250 23001 8432 23045
rect 8740 23001 9293 23047
rect 7547 22865 9293 23001
rect 9297 22882 9383 23039
rect 10464 23009 10646 23053
rect 10954 23009 11507 23055
rect 9761 22873 11507 23009
rect 11511 22890 11597 23047
rect 12664 22991 12846 23035
rect 13154 22991 13707 23037
rect 7575 22827 7609 22865
rect 9789 22835 9823 22873
rect 11961 22855 13707 22991
rect 13711 22872 13797 23029
rect 14878 22999 15060 23043
rect 15368 22999 15921 23045
rect 14175 22863 15921 22999
rect 15925 22880 16011 23037
rect 17184 23007 17366 23051
rect 17674 23007 18227 23053
rect 16481 22871 18227 23007
rect 18231 22888 18317 23045
rect 11989 22817 12023 22855
rect 14203 22825 14237 22863
rect 16509 22833 16543 22871
rect 16558 17667 16592 17701
rect 17432 17669 17466 17703
rect 16558 17663 16579 17667
rect 17432 17665 17453 17669
rect 15780 17629 15814 17663
rect 15780 17625 15801 17629
rect 15484 17451 15570 17608
rect 15615 17443 15801 17625
rect 16270 17489 16356 17646
rect 16393 17481 16579 17663
rect 17136 17491 17222 17648
rect 17267 17483 17453 17665
rect 18200 17659 18234 17693
rect 19322 17661 19356 17695
rect 20196 17663 20230 17697
rect 18200 17655 18221 17659
rect 19322 17657 19343 17661
rect 20196 17659 20217 17663
rect 17914 17481 18000 17638
rect 18035 17473 18221 17655
rect 19030 17483 19116 17640
rect 19157 17475 19343 17657
rect 19896 17485 19982 17642
rect 20031 17477 20217 17659
rect 20964 17653 20998 17687
rect 20964 17649 20985 17653
rect 20666 17475 20752 17632
rect 20799 17467 20985 17649
rect 21578 17651 21612 17685
rect 22452 17653 22486 17687
rect 21578 17647 21599 17651
rect 22452 17649 22473 17653
rect 21413 17465 21599 17647
rect 21644 17473 21730 17630
rect 22152 17475 22238 17632
rect 22287 17467 22473 17649
rect 23220 17643 23254 17677
rect 23220 17639 23241 17643
rect 23055 17457 23241 17639
rect 23284 17465 23370 17622
rect 9343 16067 9977 16249
rect 9363 16029 9397 16067
rect 9661 15487 9851 15505
rect 9465 15323 9851 15487
rect 11890 15349 12117 15395
rect 9465 15319 9495 15323
rect 9461 15285 9495 15319
rect 11475 15213 12117 15349
rect 11503 15175 11537 15213
rect 10845 14877 11035 14895
rect 10649 14713 11035 14877
rect 10649 14709 10679 14713
rect 9353 14503 9987 14685
rect 10645 14675 10679 14709
rect 9373 14465 9407 14503
rect 9671 13923 9861 13941
rect 9475 13759 9861 13923
rect 11106 13883 11333 13929
rect 9475 13755 9505 13759
rect 9471 13721 9505 13755
rect 10691 13747 11333 13883
rect 10719 13709 10753 13747
rect 12950 13873 13139 13913
rect 12589 13737 13139 13873
rect 12618 13693 12652 13737
rect 12950 13731 13139 13737
rect 11871 13509 12057 13555
rect 11690 13373 12057 13509
rect 11690 13369 11723 13373
rect 11689 13335 11723 13369
rect 11089 13041 11273 13087
rect 9345 12835 9979 13017
rect 10815 12905 11273 13041
rect 10843 12867 10877 12905
rect 9365 12797 9399 12835
rect 9663 12255 9853 12273
rect 9467 12091 9853 12255
rect 9467 12087 9497 12091
rect 9463 12053 9497 12087
rect 11039 12049 11229 12067
rect 10843 11885 11229 12049
rect 10843 11881 10873 11885
rect 10839 11847 10873 11881
rect 9355 11271 9989 11453
rect 9375 11233 9409 11271
rect 9673 10691 9863 10709
rect 9477 10527 9863 10691
rect 9477 10523 9507 10527
rect 9473 10489 9507 10523
rect 6325 6583 6359 6617
rect 6325 6579 6346 6583
rect 6160 6397 6346 6579
rect 11426 5947 11460 5985
rect 10054 5811 11489 5947
rect 13488 5935 13522 5973
rect 15446 5943 15480 5981
rect 17440 5949 17474 5987
rect 10054 5765 10240 5811
rect 11303 5765 11489 5811
rect 12116 5799 13551 5935
rect 12116 5753 12302 5799
rect 13365 5753 13551 5799
rect 14074 5807 15509 5943
rect 14074 5761 14260 5807
rect 15323 5761 15509 5807
rect 16068 5813 17503 5949
rect 16068 5767 16254 5813
rect 17317 5767 17503 5813
rect 3244 5527 3278 5565
rect 1872 5391 3307 5527
rect 5378 5519 5412 5557
rect 7330 5519 7364 5557
rect 9332 5525 9366 5563
rect 1872 5345 2058 5391
rect 3121 5345 3307 5391
rect 4006 5383 5441 5519
rect 4006 5337 4192 5383
rect 5255 5337 5441 5383
rect 5958 5383 7393 5519
rect 5958 5337 6144 5383
rect 7207 5337 7393 5383
rect 7960 5389 9395 5525
rect 7960 5343 8146 5389
rect 9209 5343 9395 5389
rect 11454 5073 11488 5111
rect 10082 4937 11517 5073
rect 13724 5029 13758 5067
rect 10082 4891 10268 4937
rect 11331 4891 11517 4937
rect 12352 4893 13787 5029
rect 15726 5023 15760 5061
rect 12352 4847 12538 4893
rect 13601 4847 13787 4893
rect 14354 4887 15789 5023
rect 17748 5005 17782 5043
rect 14354 4841 14540 4887
rect 15603 4841 15789 4887
rect 16376 4869 17811 5005
rect 16376 4823 16562 4869
rect 17625 4823 17811 4869
rect 3214 2267 3248 2305
rect 1842 2131 3277 2267
rect 5284 2263 5318 2301
rect 7236 2263 7270 2301
rect 9238 2269 9272 2307
rect 11190 2269 11224 2307
rect 13182 2269 13216 2307
rect 15134 2269 15168 2307
rect 17198 2269 17232 2307
rect 1842 2085 2028 2131
rect 3091 2085 3277 2131
rect 3912 2127 5347 2263
rect 3912 2081 4098 2127
rect 5161 2081 5347 2127
rect 5864 2127 7299 2263
rect 5864 2081 6050 2127
rect 7113 2081 7299 2127
rect 7866 2133 9301 2269
rect 7866 2087 8052 2133
rect 9115 2087 9301 2133
rect 9818 2133 11253 2269
rect 9818 2087 10004 2133
rect 11067 2087 11253 2133
rect 11810 2133 13245 2269
rect 11810 2087 11996 2133
rect 13059 2087 13245 2133
rect 13762 2133 15197 2269
rect 13762 2087 13948 2133
rect 15011 2087 15197 2133
rect 15826 2133 17261 2269
rect 15826 2087 16012 2133
rect 17075 2087 17261 2133
<< ndiff >>
rect 18833 35099 18963 35107
rect 18833 35065 18879 35099
rect 18913 35065 18963 35099
rect 18833 35055 18963 35065
rect 18833 35015 18963 35025
rect 18833 34981 18917 35015
rect 18951 34981 18963 35015
rect 18833 34975 18963 34981
rect 18879 34960 18963 34975
rect 18879 34920 18963 34930
rect 18879 34886 18891 34920
rect 18925 34886 18963 34920
rect 18879 34878 18963 34886
rect 18833 34816 18963 34824
rect 18833 34782 18846 34816
rect 18880 34782 18914 34816
rect 18948 34782 18963 34816
rect 18833 34772 18963 34782
rect 18833 34732 18963 34742
rect 18833 34698 18887 34732
rect 18921 34698 18963 34732
rect 18833 34688 18963 34698
rect 18833 34648 18963 34658
rect 18833 34614 18848 34648
rect 18882 34614 18916 34648
rect 18950 34614 18963 34648
rect 18833 34606 18963 34614
rect 18879 34542 18963 34550
rect 18879 34508 18903 34542
rect 18937 34508 18963 34542
rect 18879 34498 18963 34508
rect 18879 34418 18963 34468
rect 18891 34403 18963 34418
rect 18891 34344 18963 34373
rect 18891 34310 18903 34344
rect 18937 34310 18963 34344
rect 18891 34297 18963 34310
rect 18891 34246 18963 34267
rect 18835 34241 18963 34246
rect 18835 34207 18903 34241
rect 18937 34207 18963 34241
rect 18835 34196 18963 34207
rect 18835 34122 18963 34166
rect 18835 34116 18909 34122
rect 18879 34088 18909 34116
rect 18943 34088 18963 34122
rect 18879 34077 18963 34088
rect 18879 33997 18963 34047
rect 18891 33978 18963 33997
rect 18891 33923 18963 33948
rect 18891 33889 18903 33923
rect 18937 33889 18963 33923
rect 18891 33879 18963 33889
rect 18891 33817 18963 33849
rect 18879 33812 18963 33817
rect 18879 33778 18903 33812
rect 18937 33778 18963 33812
rect 18879 33767 18963 33778
rect 18879 33727 18963 33737
rect 18879 33693 18917 33727
rect 18951 33693 18963 33727
rect 18879 33685 18963 33693
rect 18879 33623 18963 33631
rect 18879 33589 18891 33623
rect 18925 33589 18963 33623
rect 18879 33579 18963 33589
rect 18879 33539 18963 33549
rect 18879 33505 18917 33539
rect 18951 33505 18963 33539
rect 18879 33495 18963 33505
rect 18879 33455 18963 33465
rect 18879 33421 18891 33455
rect 18925 33421 18963 33455
rect 18879 33413 18963 33421
rect 18841 32793 18971 32801
rect 18841 32759 18887 32793
rect 18921 32759 18971 32793
rect 18841 32749 18971 32759
rect 18841 32709 18971 32719
rect 18841 32675 18925 32709
rect 18959 32675 18971 32709
rect 18841 32669 18971 32675
rect 18887 32654 18971 32669
rect 18887 32614 18971 32624
rect 18887 32580 18899 32614
rect 18933 32580 18971 32614
rect 18887 32572 18971 32580
rect 18841 32510 18971 32518
rect 18841 32476 18854 32510
rect 18888 32476 18922 32510
rect 18956 32476 18971 32510
rect 18841 32466 18971 32476
rect 18841 32426 18971 32436
rect 18841 32392 18895 32426
rect 18929 32392 18971 32426
rect 18841 32382 18971 32392
rect 18841 32342 18971 32352
rect 18841 32308 18856 32342
rect 18890 32308 18924 32342
rect 18958 32308 18971 32342
rect 18841 32300 18971 32308
rect 18887 32236 18971 32244
rect 18887 32202 18911 32236
rect 18945 32202 18971 32236
rect 18887 32192 18971 32202
rect 18887 32112 18971 32162
rect 18899 32097 18971 32112
rect 18899 32038 18971 32067
rect 18899 32004 18911 32038
rect 18945 32004 18971 32038
rect 18899 31991 18971 32004
rect 18899 31940 18971 31961
rect 18843 31935 18971 31940
rect 18843 31901 18911 31935
rect 18945 31901 18971 31935
rect 18843 31890 18971 31901
rect 18843 31816 18971 31860
rect 18843 31810 18917 31816
rect 18887 31782 18917 31810
rect 18951 31782 18971 31816
rect 18887 31771 18971 31782
rect 18887 31691 18971 31741
rect 18899 31672 18971 31691
rect 18899 31617 18971 31642
rect 18899 31583 18911 31617
rect 18945 31583 18971 31617
rect 18899 31573 18971 31583
rect 18899 31511 18971 31543
rect 18887 31506 18971 31511
rect 18887 31472 18911 31506
rect 18945 31472 18971 31506
rect 18887 31461 18971 31472
rect 18887 31421 18971 31431
rect 18887 31387 18925 31421
rect 18959 31387 18971 31421
rect 18887 31379 18971 31387
rect 18887 31317 18971 31325
rect 18887 31283 18899 31317
rect 18933 31283 18971 31317
rect 18887 31273 18971 31283
rect 18887 31233 18971 31243
rect 18887 31199 18925 31233
rect 18959 31199 18971 31233
rect 18887 31189 18971 31199
rect 18887 31149 18971 31159
rect 18887 31115 18899 31149
rect 18933 31115 18971 31149
rect 18887 31107 18971 31115
rect 18849 30579 18979 30587
rect 18849 30545 18895 30579
rect 18929 30545 18979 30579
rect 18849 30535 18979 30545
rect 18849 30495 18979 30505
rect 18849 30461 18933 30495
rect 18967 30461 18979 30495
rect 18849 30455 18979 30461
rect 18895 30440 18979 30455
rect 18895 30400 18979 30410
rect 18895 30366 18907 30400
rect 18941 30366 18979 30400
rect 18895 30358 18979 30366
rect 18849 30296 18979 30304
rect 18849 30262 18862 30296
rect 18896 30262 18930 30296
rect 18964 30262 18979 30296
rect 18849 30252 18979 30262
rect 18849 30212 18979 30222
rect 18849 30178 18903 30212
rect 18937 30178 18979 30212
rect 18849 30168 18979 30178
rect 18849 30128 18979 30138
rect 18849 30094 18864 30128
rect 18898 30094 18932 30128
rect 18966 30094 18979 30128
rect 18849 30086 18979 30094
rect 18895 30022 18979 30030
rect 18895 29988 18919 30022
rect 18953 29988 18979 30022
rect 18895 29978 18979 29988
rect 18895 29898 18979 29948
rect 18907 29883 18979 29898
rect 18907 29824 18979 29853
rect 18907 29790 18919 29824
rect 18953 29790 18979 29824
rect 18907 29777 18979 29790
rect 18907 29726 18979 29747
rect 18851 29721 18979 29726
rect 18851 29687 18919 29721
rect 18953 29687 18979 29721
rect 18851 29676 18979 29687
rect 18851 29602 18979 29646
rect 18851 29596 18925 29602
rect 18895 29568 18925 29596
rect 18959 29568 18979 29602
rect 18895 29557 18979 29568
rect 18895 29477 18979 29527
rect 18907 29458 18979 29477
rect 18907 29403 18979 29428
rect 18907 29369 18919 29403
rect 18953 29369 18979 29403
rect 18907 29359 18979 29369
rect 18907 29297 18979 29329
rect 18895 29292 18979 29297
rect 18895 29258 18919 29292
rect 18953 29258 18979 29292
rect 18895 29247 18979 29258
rect 18895 29207 18979 29217
rect 18895 29173 18933 29207
rect 18967 29173 18979 29207
rect 18895 29165 18979 29173
rect 18895 29103 18979 29111
rect 18895 29069 18907 29103
rect 18941 29069 18979 29103
rect 18895 29059 18979 29069
rect 18895 29019 18979 29029
rect 18895 28985 18933 29019
rect 18967 28985 18979 29019
rect 18895 28975 18979 28985
rect 18895 28935 18979 28945
rect 18895 28901 18907 28935
rect 18941 28901 18979 28935
rect 18895 28893 18979 28901
rect 18831 28379 18961 28387
rect 18831 28345 18877 28379
rect 18911 28345 18961 28379
rect 18831 28335 18961 28345
rect 18831 28295 18961 28305
rect 18831 28261 18915 28295
rect 18949 28261 18961 28295
rect 18831 28255 18961 28261
rect 18877 28240 18961 28255
rect 18877 28200 18961 28210
rect 18877 28166 18889 28200
rect 18923 28166 18961 28200
rect 18877 28158 18961 28166
rect 18831 28096 18961 28104
rect 18831 28062 18844 28096
rect 18878 28062 18912 28096
rect 18946 28062 18961 28096
rect 18831 28052 18961 28062
rect 18831 28012 18961 28022
rect 18831 27978 18885 28012
rect 18919 27978 18961 28012
rect 18831 27968 18961 27978
rect 18831 27928 18961 27938
rect 18831 27894 18846 27928
rect 18880 27894 18914 27928
rect 18948 27894 18961 27928
rect 18831 27886 18961 27894
rect 18877 27822 18961 27830
rect 18877 27788 18901 27822
rect 18935 27788 18961 27822
rect 18877 27778 18961 27788
rect 18877 27698 18961 27748
rect 18889 27683 18961 27698
rect 18889 27624 18961 27653
rect 18889 27590 18901 27624
rect 18935 27590 18961 27624
rect 18889 27577 18961 27590
rect 18889 27526 18961 27547
rect 18833 27521 18961 27526
rect 18833 27487 18901 27521
rect 18935 27487 18961 27521
rect 18833 27476 18961 27487
rect 18833 27402 18961 27446
rect 18833 27396 18907 27402
rect 18877 27368 18907 27396
rect 18941 27368 18961 27402
rect 18877 27357 18961 27368
rect 18877 27277 18961 27327
rect 18889 27258 18961 27277
rect 18889 27203 18961 27228
rect 18889 27169 18901 27203
rect 18935 27169 18961 27203
rect 18889 27159 18961 27169
rect 18889 27097 18961 27129
rect 18877 27092 18961 27097
rect 18877 27058 18901 27092
rect 18935 27058 18961 27092
rect 18877 27047 18961 27058
rect 18877 27007 18961 27017
rect 18877 26973 18915 27007
rect 18949 26973 18961 27007
rect 18877 26965 18961 26973
rect 18877 26903 18961 26911
rect 18877 26869 18889 26903
rect 18923 26869 18961 26903
rect 18877 26859 18961 26869
rect 18877 26819 18961 26829
rect 18877 26785 18915 26819
rect 18949 26785 18961 26819
rect 18877 26775 18961 26785
rect 18877 26735 18961 26745
rect 18877 26701 18889 26735
rect 18923 26701 18961 26735
rect 18877 26693 18961 26701
rect 18839 26165 18969 26173
rect 18839 26131 18885 26165
rect 18919 26131 18969 26165
rect 18839 26121 18969 26131
rect 18839 26081 18969 26091
rect 18839 26047 18923 26081
rect 18957 26047 18969 26081
rect 18839 26041 18969 26047
rect 18885 26026 18969 26041
rect 18885 25986 18969 25996
rect 18885 25952 18897 25986
rect 18931 25952 18969 25986
rect 18885 25944 18969 25952
rect 18839 25882 18969 25890
rect 18839 25848 18852 25882
rect 18886 25848 18920 25882
rect 18954 25848 18969 25882
rect 18839 25838 18969 25848
rect 18839 25798 18969 25808
rect 18839 25764 18893 25798
rect 18927 25764 18969 25798
rect 18839 25754 18969 25764
rect 18839 25714 18969 25724
rect 18839 25680 18854 25714
rect 18888 25680 18922 25714
rect 18956 25680 18969 25714
rect 18839 25672 18969 25680
rect 18885 25608 18969 25616
rect 18885 25574 18909 25608
rect 18943 25574 18969 25608
rect 18885 25564 18969 25574
rect 18885 25484 18969 25534
rect 18897 25469 18969 25484
rect 18897 25410 18969 25439
rect 18897 25376 18909 25410
rect 18943 25376 18969 25410
rect 18897 25363 18969 25376
rect 18897 25312 18969 25333
rect 18841 25307 18969 25312
rect 18841 25273 18909 25307
rect 18943 25273 18969 25307
rect 18841 25262 18969 25273
rect 18841 25188 18969 25232
rect 18841 25182 18915 25188
rect 18885 25154 18915 25182
rect 18949 25154 18969 25188
rect 18885 25143 18969 25154
rect 18885 25063 18969 25113
rect 18897 25044 18969 25063
rect 18897 24989 18969 25014
rect 18897 24955 18909 24989
rect 18943 24955 18969 24989
rect 18897 24945 18969 24955
rect 18897 24883 18969 24915
rect 18885 24878 18969 24883
rect 18885 24844 18909 24878
rect 18943 24844 18969 24878
rect 18885 24833 18969 24844
rect 18885 24793 18969 24803
rect 18885 24759 18923 24793
rect 18957 24759 18969 24793
rect 18885 24751 18969 24759
rect 18885 24689 18969 24697
rect 18885 24655 18897 24689
rect 18931 24655 18969 24689
rect 18885 24645 18969 24655
rect 18885 24605 18969 24615
rect 18885 24571 18923 24605
rect 18957 24571 18969 24605
rect 18885 24561 18969 24571
rect 18885 24521 18969 24531
rect 18885 24487 18897 24521
rect 18931 24487 18969 24521
rect 18885 24479 18969 24487
rect 7573 22963 7625 22975
rect 7573 22929 7581 22963
rect 7615 22929 7625 22963
rect 7573 22891 7625 22929
rect 7655 22937 7709 22975
rect 7655 22903 7665 22937
rect 7699 22903 7709 22937
rect 7655 22891 7709 22903
rect 7739 22963 7791 22975
rect 7739 22929 7749 22963
rect 7783 22929 7791 22963
rect 7739 22891 7791 22929
rect 7845 22937 7897 22975
rect 7845 22903 7853 22937
rect 7887 22903 7897 22937
rect 7845 22891 7897 22903
rect 7927 22963 7977 22975
rect 8276 22975 8326 23019
rect 8157 22963 8207 22975
rect 7927 22951 8009 22963
rect 7927 22917 7938 22951
rect 7972 22917 8009 22951
rect 7927 22891 8009 22917
rect 8039 22951 8108 22963
rect 8039 22917 8049 22951
rect 8083 22917 8108 22951
rect 8039 22891 8108 22917
rect 8138 22891 8207 22963
rect 8237 22945 8326 22975
rect 8237 22911 8248 22945
rect 8282 22911 8326 22945
rect 8237 22891 8326 22911
rect 8356 22963 8406 23019
rect 8766 23006 8818 23021
rect 8578 22963 8628 22975
rect 8356 22951 8427 22963
rect 8356 22917 8367 22951
rect 8401 22917 8427 22951
rect 8356 22891 8427 22917
rect 8457 22951 8533 22963
rect 8457 22917 8470 22951
rect 8504 22917 8533 22951
rect 8457 22891 8533 22917
rect 8563 22891 8628 22963
rect 8658 22951 8710 22975
rect 8658 22917 8668 22951
rect 8702 22917 8710 22951
rect 8658 22891 8710 22917
rect 8766 22972 8774 23006
rect 8808 22972 8818 23006
rect 8766 22938 8818 22972
rect 8766 22904 8774 22938
rect 8808 22904 8818 22938
rect 8766 22891 8818 22904
rect 8848 22967 8902 23021
rect 8848 22933 8858 22967
rect 8892 22933 8902 22967
rect 8848 22891 8902 22933
rect 8932 23008 8984 23021
rect 8932 22974 8942 23008
rect 8976 22974 8984 23008
rect 9135 22975 9185 23021
rect 8932 22940 8984 22974
rect 8932 22906 8942 22940
rect 8976 22906 8984 22940
rect 8932 22891 8984 22906
rect 9038 22963 9090 22975
rect 9038 22929 9046 22963
rect 9080 22929 9090 22963
rect 9038 22891 9090 22929
rect 9120 22937 9185 22975
rect 9120 22903 9141 22937
rect 9175 22903 9185 22937
rect 9120 22891 9185 22903
rect 9215 22975 9267 23021
rect 9215 22941 9225 22975
rect 9259 22941 9267 22975
rect 9215 22891 9267 22941
rect 9787 22971 9839 22983
rect 9787 22937 9795 22971
rect 9829 22937 9839 22971
rect 9787 22899 9839 22937
rect 9869 22945 9923 22983
rect 9869 22911 9879 22945
rect 9913 22911 9923 22945
rect 9869 22899 9923 22911
rect 9953 22971 10005 22983
rect 9953 22937 9963 22971
rect 9997 22937 10005 22971
rect 9953 22899 10005 22937
rect 10059 22945 10111 22983
rect 10059 22911 10067 22945
rect 10101 22911 10111 22945
rect 10059 22899 10111 22911
rect 10141 22971 10191 22983
rect 10490 22983 10540 23027
rect 10371 22971 10421 22983
rect 10141 22959 10223 22971
rect 10141 22925 10152 22959
rect 10186 22925 10223 22959
rect 10141 22899 10223 22925
rect 10253 22959 10322 22971
rect 10253 22925 10263 22959
rect 10297 22925 10322 22959
rect 10253 22899 10322 22925
rect 10352 22899 10421 22971
rect 10451 22953 10540 22983
rect 10451 22919 10462 22953
rect 10496 22919 10540 22953
rect 10451 22899 10540 22919
rect 10570 22971 10620 23027
rect 10980 23014 11032 23029
rect 10792 22971 10842 22983
rect 10570 22959 10641 22971
rect 10570 22925 10581 22959
rect 10615 22925 10641 22959
rect 10570 22899 10641 22925
rect 10671 22959 10747 22971
rect 10671 22925 10684 22959
rect 10718 22925 10747 22959
rect 10671 22899 10747 22925
rect 10777 22899 10842 22971
rect 10872 22959 10924 22983
rect 10872 22925 10882 22959
rect 10916 22925 10924 22959
rect 10872 22899 10924 22925
rect 10980 22980 10988 23014
rect 11022 22980 11032 23014
rect 10980 22946 11032 22980
rect 10980 22912 10988 22946
rect 11022 22912 11032 22946
rect 10980 22899 11032 22912
rect 11062 22975 11116 23029
rect 11062 22941 11072 22975
rect 11106 22941 11116 22975
rect 11062 22899 11116 22941
rect 11146 23016 11198 23029
rect 11146 22982 11156 23016
rect 11190 22982 11198 23016
rect 11349 22983 11399 23029
rect 11146 22948 11198 22982
rect 11146 22914 11156 22948
rect 11190 22914 11198 22948
rect 11146 22899 11198 22914
rect 11252 22971 11304 22983
rect 11252 22937 11260 22971
rect 11294 22937 11304 22971
rect 11252 22899 11304 22937
rect 11334 22945 11399 22983
rect 11334 22911 11355 22945
rect 11389 22911 11399 22945
rect 11334 22899 11399 22911
rect 11429 22983 11481 23029
rect 11429 22949 11439 22983
rect 11473 22949 11481 22983
rect 11429 22899 11481 22949
rect 11987 22953 12039 22965
rect 11987 22919 11995 22953
rect 12029 22919 12039 22953
rect 11987 22881 12039 22919
rect 12069 22927 12123 22965
rect 12069 22893 12079 22927
rect 12113 22893 12123 22927
rect 12069 22881 12123 22893
rect 12153 22953 12205 22965
rect 12153 22919 12163 22953
rect 12197 22919 12205 22953
rect 12153 22881 12205 22919
rect 12259 22927 12311 22965
rect 12259 22893 12267 22927
rect 12301 22893 12311 22927
rect 12259 22881 12311 22893
rect 12341 22953 12391 22965
rect 12690 22965 12740 23009
rect 12571 22953 12621 22965
rect 12341 22941 12423 22953
rect 12341 22907 12352 22941
rect 12386 22907 12423 22941
rect 12341 22881 12423 22907
rect 12453 22941 12522 22953
rect 12453 22907 12463 22941
rect 12497 22907 12522 22941
rect 12453 22881 12522 22907
rect 12552 22881 12621 22953
rect 12651 22935 12740 22965
rect 12651 22901 12662 22935
rect 12696 22901 12740 22935
rect 12651 22881 12740 22901
rect 12770 22953 12820 23009
rect 13180 22996 13232 23011
rect 12992 22953 13042 22965
rect 12770 22941 12841 22953
rect 12770 22907 12781 22941
rect 12815 22907 12841 22941
rect 12770 22881 12841 22907
rect 12871 22941 12947 22953
rect 12871 22907 12884 22941
rect 12918 22907 12947 22941
rect 12871 22881 12947 22907
rect 12977 22881 13042 22953
rect 13072 22941 13124 22965
rect 13072 22907 13082 22941
rect 13116 22907 13124 22941
rect 13072 22881 13124 22907
rect 13180 22962 13188 22996
rect 13222 22962 13232 22996
rect 13180 22928 13232 22962
rect 13180 22894 13188 22928
rect 13222 22894 13232 22928
rect 13180 22881 13232 22894
rect 13262 22957 13316 23011
rect 13262 22923 13272 22957
rect 13306 22923 13316 22957
rect 13262 22881 13316 22923
rect 13346 22998 13398 23011
rect 13346 22964 13356 22998
rect 13390 22964 13398 22998
rect 13549 22965 13599 23011
rect 13346 22930 13398 22964
rect 13346 22896 13356 22930
rect 13390 22896 13398 22930
rect 13346 22881 13398 22896
rect 13452 22953 13504 22965
rect 13452 22919 13460 22953
rect 13494 22919 13504 22953
rect 13452 22881 13504 22919
rect 13534 22927 13599 22965
rect 13534 22893 13555 22927
rect 13589 22893 13599 22927
rect 13534 22881 13599 22893
rect 13629 22965 13681 23011
rect 13629 22931 13639 22965
rect 13673 22931 13681 22965
rect 13629 22881 13681 22931
rect 14201 22961 14253 22973
rect 14201 22927 14209 22961
rect 14243 22927 14253 22961
rect 14201 22889 14253 22927
rect 14283 22935 14337 22973
rect 14283 22901 14293 22935
rect 14327 22901 14337 22935
rect 14283 22889 14337 22901
rect 14367 22961 14419 22973
rect 14367 22927 14377 22961
rect 14411 22927 14419 22961
rect 14367 22889 14419 22927
rect 14473 22935 14525 22973
rect 14473 22901 14481 22935
rect 14515 22901 14525 22935
rect 14473 22889 14525 22901
rect 14555 22961 14605 22973
rect 14904 22973 14954 23017
rect 14785 22961 14835 22973
rect 14555 22949 14637 22961
rect 14555 22915 14566 22949
rect 14600 22915 14637 22949
rect 14555 22889 14637 22915
rect 14667 22949 14736 22961
rect 14667 22915 14677 22949
rect 14711 22915 14736 22949
rect 14667 22889 14736 22915
rect 14766 22889 14835 22961
rect 14865 22943 14954 22973
rect 14865 22909 14876 22943
rect 14910 22909 14954 22943
rect 14865 22889 14954 22909
rect 14984 22961 15034 23017
rect 15394 23004 15446 23019
rect 15206 22961 15256 22973
rect 14984 22949 15055 22961
rect 14984 22915 14995 22949
rect 15029 22915 15055 22949
rect 14984 22889 15055 22915
rect 15085 22949 15161 22961
rect 15085 22915 15098 22949
rect 15132 22915 15161 22949
rect 15085 22889 15161 22915
rect 15191 22889 15256 22961
rect 15286 22949 15338 22973
rect 15286 22915 15296 22949
rect 15330 22915 15338 22949
rect 15286 22889 15338 22915
rect 15394 22970 15402 23004
rect 15436 22970 15446 23004
rect 15394 22936 15446 22970
rect 15394 22902 15402 22936
rect 15436 22902 15446 22936
rect 15394 22889 15446 22902
rect 15476 22965 15530 23019
rect 15476 22931 15486 22965
rect 15520 22931 15530 22965
rect 15476 22889 15530 22931
rect 15560 23006 15612 23019
rect 15560 22972 15570 23006
rect 15604 22972 15612 23006
rect 15763 22973 15813 23019
rect 15560 22938 15612 22972
rect 15560 22904 15570 22938
rect 15604 22904 15612 22938
rect 15560 22889 15612 22904
rect 15666 22961 15718 22973
rect 15666 22927 15674 22961
rect 15708 22927 15718 22961
rect 15666 22889 15718 22927
rect 15748 22935 15813 22973
rect 15748 22901 15769 22935
rect 15803 22901 15813 22935
rect 15748 22889 15813 22901
rect 15843 22973 15895 23019
rect 15843 22939 15853 22973
rect 15887 22939 15895 22973
rect 15843 22889 15895 22939
rect 16507 22969 16559 22981
rect 16507 22935 16515 22969
rect 16549 22935 16559 22969
rect 16507 22897 16559 22935
rect 16589 22943 16643 22981
rect 16589 22909 16599 22943
rect 16633 22909 16643 22943
rect 16589 22897 16643 22909
rect 16673 22969 16725 22981
rect 16673 22935 16683 22969
rect 16717 22935 16725 22969
rect 16673 22897 16725 22935
rect 16779 22943 16831 22981
rect 16779 22909 16787 22943
rect 16821 22909 16831 22943
rect 16779 22897 16831 22909
rect 16861 22969 16911 22981
rect 17210 22981 17260 23025
rect 17091 22969 17141 22981
rect 16861 22957 16943 22969
rect 16861 22923 16872 22957
rect 16906 22923 16943 22957
rect 16861 22897 16943 22923
rect 16973 22957 17042 22969
rect 16973 22923 16983 22957
rect 17017 22923 17042 22957
rect 16973 22897 17042 22923
rect 17072 22897 17141 22969
rect 17171 22951 17260 22981
rect 17171 22917 17182 22951
rect 17216 22917 17260 22951
rect 17171 22897 17260 22917
rect 17290 22969 17340 23025
rect 17700 23012 17752 23027
rect 17512 22969 17562 22981
rect 17290 22957 17361 22969
rect 17290 22923 17301 22957
rect 17335 22923 17361 22957
rect 17290 22897 17361 22923
rect 17391 22957 17467 22969
rect 17391 22923 17404 22957
rect 17438 22923 17467 22957
rect 17391 22897 17467 22923
rect 17497 22897 17562 22969
rect 17592 22957 17644 22981
rect 17592 22923 17602 22957
rect 17636 22923 17644 22957
rect 17592 22897 17644 22923
rect 17700 22978 17708 23012
rect 17742 22978 17752 23012
rect 17700 22944 17752 22978
rect 17700 22910 17708 22944
rect 17742 22910 17752 22944
rect 17700 22897 17752 22910
rect 17782 22973 17836 23027
rect 17782 22939 17792 22973
rect 17826 22939 17836 22973
rect 17782 22897 17836 22939
rect 17866 23014 17918 23027
rect 17866 22980 17876 23014
rect 17910 22980 17918 23014
rect 18069 22981 18119 23027
rect 17866 22946 17918 22980
rect 17866 22912 17876 22946
rect 17910 22912 17918 22946
rect 17866 22897 17918 22912
rect 17972 22969 18024 22981
rect 17972 22935 17980 22969
rect 18014 22935 18024 22969
rect 17972 22897 18024 22935
rect 18054 22943 18119 22981
rect 18054 22909 18075 22943
rect 18109 22909 18119 22943
rect 18054 22897 18119 22909
rect 18149 22981 18201 23027
rect 18149 22947 18159 22981
rect 18193 22947 18201 22981
rect 18149 22897 18201 22947
rect 16419 17621 16471 17637
rect 15641 17583 15693 17599
rect 15641 17549 15649 17583
rect 15683 17549 15693 17583
rect 15641 17515 15693 17549
rect 15641 17481 15649 17515
rect 15683 17481 15693 17515
rect 15641 17469 15693 17481
rect 15723 17583 15775 17599
rect 15723 17549 15733 17583
rect 15767 17549 15775 17583
rect 15723 17515 15775 17549
rect 16419 17587 16427 17621
rect 16461 17587 16471 17621
rect 16419 17553 16471 17587
rect 16419 17519 16427 17553
rect 16461 17519 16471 17553
rect 15723 17481 15733 17515
rect 15767 17481 15775 17515
rect 16419 17507 16471 17519
rect 16501 17621 16553 17637
rect 17293 17623 17345 17639
rect 16501 17587 16511 17621
rect 16545 17587 16553 17621
rect 16501 17553 16553 17587
rect 16501 17519 16511 17553
rect 16545 17519 16553 17553
rect 16501 17507 16553 17519
rect 17293 17589 17301 17623
rect 17335 17589 17345 17623
rect 17293 17555 17345 17589
rect 17293 17521 17301 17555
rect 17335 17521 17345 17555
rect 17293 17509 17345 17521
rect 17375 17623 17427 17639
rect 17375 17589 17385 17623
rect 17419 17589 17427 17623
rect 18061 17613 18113 17629
rect 17375 17555 17427 17589
rect 17375 17521 17385 17555
rect 17419 17521 17427 17555
rect 17375 17509 17427 17521
rect 15723 17469 15775 17481
rect 18061 17579 18069 17613
rect 18103 17579 18113 17613
rect 18061 17545 18113 17579
rect 18061 17511 18069 17545
rect 18103 17511 18113 17545
rect 18061 17499 18113 17511
rect 18143 17613 18195 17629
rect 19183 17615 19235 17631
rect 18143 17579 18153 17613
rect 18187 17579 18195 17613
rect 18143 17545 18195 17579
rect 18143 17511 18153 17545
rect 18187 17511 18195 17545
rect 18143 17499 18195 17511
rect 19183 17581 19191 17615
rect 19225 17581 19235 17615
rect 19183 17547 19235 17581
rect 19183 17513 19191 17547
rect 19225 17513 19235 17547
rect 19183 17501 19235 17513
rect 19265 17615 19317 17631
rect 20057 17617 20109 17633
rect 19265 17581 19275 17615
rect 19309 17581 19317 17615
rect 19265 17547 19317 17581
rect 19265 17513 19275 17547
rect 19309 17513 19317 17547
rect 19265 17501 19317 17513
rect 20057 17583 20065 17617
rect 20099 17583 20109 17617
rect 20057 17549 20109 17583
rect 20057 17515 20065 17549
rect 20099 17515 20109 17549
rect 20057 17503 20109 17515
rect 20139 17617 20191 17633
rect 20139 17583 20149 17617
rect 20183 17583 20191 17617
rect 20825 17607 20877 17623
rect 20139 17549 20191 17583
rect 20139 17515 20149 17549
rect 20183 17515 20191 17549
rect 20139 17503 20191 17515
rect 20825 17573 20833 17607
rect 20867 17573 20877 17607
rect 20825 17539 20877 17573
rect 20825 17505 20833 17539
rect 20867 17505 20877 17539
rect 20825 17493 20877 17505
rect 20907 17607 20959 17623
rect 20907 17573 20917 17607
rect 20951 17573 20959 17607
rect 20907 17539 20959 17573
rect 20907 17505 20917 17539
rect 20951 17505 20959 17539
rect 20907 17493 20959 17505
rect 21439 17605 21491 17621
rect 21439 17571 21447 17605
rect 21481 17571 21491 17605
rect 21439 17537 21491 17571
rect 21439 17503 21447 17537
rect 21481 17503 21491 17537
rect 21439 17491 21491 17503
rect 21521 17605 21573 17621
rect 22313 17607 22365 17623
rect 21521 17571 21531 17605
rect 21565 17571 21573 17605
rect 21521 17537 21573 17571
rect 21521 17503 21531 17537
rect 21565 17503 21573 17537
rect 21521 17491 21573 17503
rect 22313 17573 22321 17607
rect 22355 17573 22365 17607
rect 22313 17539 22365 17573
rect 22313 17505 22321 17539
rect 22355 17505 22365 17539
rect 22313 17493 22365 17505
rect 22395 17607 22447 17623
rect 22395 17573 22405 17607
rect 22439 17573 22447 17607
rect 22395 17539 22447 17573
rect 22395 17505 22405 17539
rect 22439 17505 22447 17539
rect 22395 17493 22447 17505
rect 23081 17597 23133 17613
rect 23081 17563 23089 17597
rect 23123 17563 23133 17597
rect 23081 17529 23133 17563
rect 23081 17495 23089 17529
rect 23123 17495 23133 17529
rect 23081 17483 23133 17495
rect 23163 17597 23215 17613
rect 23163 17563 23173 17597
rect 23207 17563 23215 17597
rect 23163 17529 23215 17563
rect 23163 17495 23173 17529
rect 23207 17495 23215 17529
rect 23163 17483 23215 17495
rect 9369 16141 9421 16223
rect 9369 16107 9377 16141
rect 9411 16107 9421 16141
rect 9369 16093 9421 16107
rect 9451 16163 9505 16223
rect 9451 16129 9461 16163
rect 9495 16129 9505 16163
rect 9451 16093 9505 16129
rect 9535 16141 9589 16223
rect 9535 16107 9545 16141
rect 9579 16107 9589 16141
rect 9535 16093 9589 16107
rect 9619 16093 9673 16223
rect 9703 16143 9857 16223
rect 9703 16109 9713 16143
rect 9747 16109 9813 16143
rect 9847 16109 9857 16143
rect 9703 16093 9857 16109
rect 9887 16214 9951 16223
rect 9887 16180 9903 16214
rect 9937 16180 9951 16214
rect 9887 16146 9951 16180
rect 9887 16112 9903 16146
rect 9937 16112 9951 16146
rect 9887 16093 9951 16112
rect 9687 15461 9739 15479
rect 9491 15423 9547 15461
rect 9491 15389 9503 15423
rect 9537 15389 9547 15423
rect 9491 15377 9547 15389
rect 9577 15377 9631 15461
rect 9661 15395 9739 15461
rect 9661 15377 9695 15395
rect 9687 15361 9695 15377
rect 9729 15361 9739 15395
rect 9687 15349 9739 15361
rect 9769 15395 9825 15479
rect 9769 15361 9779 15395
rect 9813 15361 9825 15395
rect 9769 15349 9825 15361
rect 11916 15353 12009 15369
rect 11916 15323 11950 15353
rect 11501 15293 11553 15323
rect 11501 15259 11509 15293
rect 11543 15259 11553 15293
rect 11501 15239 11553 15259
rect 11583 15239 11641 15323
rect 11671 15239 11747 15323
rect 11777 15239 11843 15323
rect 11873 15319 11950 15323
rect 11984 15319 12009 15353
rect 11873 15285 12009 15319
rect 11873 15251 11950 15285
rect 11984 15251 12009 15285
rect 11873 15239 12009 15251
rect 12039 15353 12091 15369
rect 12039 15319 12049 15353
rect 12083 15319 12091 15353
rect 12039 15285 12091 15319
rect 12039 15251 12049 15285
rect 12083 15251 12091 15285
rect 12039 15239 12091 15251
rect 10871 14851 10923 14869
rect 10675 14813 10731 14851
rect 10675 14779 10687 14813
rect 10721 14779 10731 14813
rect 10675 14767 10731 14779
rect 10761 14767 10815 14851
rect 10845 14785 10923 14851
rect 10845 14767 10879 14785
rect 10871 14751 10879 14767
rect 10913 14751 10923 14785
rect 10871 14739 10923 14751
rect 10953 14785 11009 14869
rect 10953 14751 10963 14785
rect 10997 14751 11009 14785
rect 10953 14739 11009 14751
rect 9379 14577 9431 14659
rect 9379 14543 9387 14577
rect 9421 14543 9431 14577
rect 9379 14529 9431 14543
rect 9461 14599 9515 14659
rect 9461 14565 9471 14599
rect 9505 14565 9515 14599
rect 9461 14529 9515 14565
rect 9545 14577 9599 14659
rect 9545 14543 9555 14577
rect 9589 14543 9599 14577
rect 9545 14529 9599 14543
rect 9629 14529 9683 14659
rect 9713 14579 9867 14659
rect 9713 14545 9723 14579
rect 9757 14545 9823 14579
rect 9857 14545 9867 14579
rect 9713 14529 9867 14545
rect 9897 14650 9961 14659
rect 9897 14616 9913 14650
rect 9947 14616 9961 14650
rect 9897 14582 9961 14616
rect 9897 14548 9913 14582
rect 9947 14548 9961 14582
rect 9897 14529 9961 14548
rect 9697 13897 9749 13915
rect 9501 13859 9557 13897
rect 9501 13825 9513 13859
rect 9547 13825 9557 13859
rect 9501 13813 9557 13825
rect 9587 13813 9641 13897
rect 9671 13831 9749 13897
rect 9671 13813 9705 13831
rect 9697 13797 9705 13813
rect 9739 13797 9749 13831
rect 9697 13785 9749 13797
rect 9779 13831 9835 13915
rect 11132 13887 11225 13903
rect 11132 13857 11166 13887
rect 9779 13797 9789 13831
rect 9823 13797 9835 13831
rect 9779 13785 9835 13797
rect 10717 13827 10769 13857
rect 10717 13793 10725 13827
rect 10759 13793 10769 13827
rect 10717 13773 10769 13793
rect 10799 13773 10857 13857
rect 10887 13773 10963 13857
rect 10993 13773 11059 13857
rect 11089 13853 11166 13857
rect 11200 13853 11225 13887
rect 11089 13819 11225 13853
rect 11089 13785 11166 13819
rect 11200 13785 11225 13819
rect 11089 13773 11225 13785
rect 11255 13887 11307 13903
rect 11255 13853 11265 13887
rect 11299 13853 11307 13887
rect 11255 13819 11307 13853
rect 11255 13785 11265 13819
rect 11299 13785 11307 13819
rect 11255 13773 11307 13785
rect 12976 13847 13029 13887
rect 12615 13827 12667 13847
rect 12615 13793 12623 13827
rect 12657 13793 12667 13827
rect 12615 13763 12667 13793
rect 12697 13821 12763 13847
rect 12697 13787 12713 13821
rect 12747 13787 12763 13821
rect 12697 13763 12763 13787
rect 12793 13807 12847 13847
rect 12793 13773 12803 13807
rect 12837 13773 12847 13807
rect 12793 13763 12847 13773
rect 12877 13821 12931 13847
rect 12877 13787 12887 13821
rect 12921 13787 12931 13821
rect 12877 13763 12931 13787
rect 12961 13807 13029 13847
rect 12961 13773 12981 13807
rect 13015 13773 13029 13807
rect 12961 13763 13029 13773
rect 12976 13757 13029 13763
rect 13059 13845 13113 13887
rect 13059 13811 13069 13845
rect 13103 13811 13113 13845
rect 13059 13757 13113 13811
rect 11897 13483 11949 13529
rect 11716 13455 11768 13483
rect 11716 13421 11724 13455
rect 11758 13421 11768 13455
rect 11716 13399 11768 13421
rect 11798 13455 11852 13483
rect 11798 13421 11808 13455
rect 11842 13421 11852 13455
rect 11798 13399 11852 13421
rect 11882 13455 11949 13483
rect 11882 13421 11904 13455
rect 11938 13421 11949 13455
rect 11882 13399 11949 13421
rect 11979 13515 12031 13529
rect 11979 13481 11989 13515
rect 12023 13481 12031 13515
rect 11979 13447 12031 13481
rect 11979 13413 11989 13447
rect 12023 13413 12031 13447
rect 11979 13399 12031 13413
rect 11115 13015 11165 13061
rect 9371 12909 9423 12991
rect 9371 12875 9379 12909
rect 9413 12875 9423 12909
rect 9371 12861 9423 12875
rect 9453 12931 9507 12991
rect 9453 12897 9463 12931
rect 9497 12897 9507 12931
rect 9453 12861 9507 12897
rect 9537 12909 9591 12991
rect 9537 12875 9547 12909
rect 9581 12875 9591 12909
rect 9537 12861 9591 12875
rect 9621 12861 9675 12991
rect 9705 12911 9859 12991
rect 9705 12877 9715 12911
rect 9749 12877 9815 12911
rect 9849 12877 9859 12911
rect 9705 12861 9859 12877
rect 9889 12982 9953 12991
rect 9889 12948 9905 12982
rect 9939 12948 9953 12982
rect 9889 12914 9953 12948
rect 10841 12977 10893 13015
rect 10841 12943 10849 12977
rect 10883 12943 10893 12977
rect 10841 12931 10893 12943
rect 10923 12931 10965 13015
rect 10995 12931 11037 13015
rect 11067 12993 11165 13015
rect 11067 12959 11121 12993
rect 11155 12959 11165 12993
rect 11067 12931 11165 12959
rect 11195 13003 11247 13061
rect 11195 12969 11205 13003
rect 11239 12969 11247 13003
rect 11195 12931 11247 12969
rect 9889 12880 9905 12914
rect 9939 12880 9953 12914
rect 9889 12861 9953 12880
rect 9689 12229 9741 12247
rect 9493 12191 9549 12229
rect 9493 12157 9505 12191
rect 9539 12157 9549 12191
rect 9493 12145 9549 12157
rect 9579 12145 9633 12229
rect 9663 12163 9741 12229
rect 9663 12145 9697 12163
rect 9689 12129 9697 12145
rect 9731 12129 9741 12163
rect 9689 12117 9741 12129
rect 9771 12163 9827 12247
rect 9771 12129 9781 12163
rect 9815 12129 9827 12163
rect 9771 12117 9827 12129
rect 11065 12023 11117 12041
rect 10869 11985 10925 12023
rect 10869 11951 10881 11985
rect 10915 11951 10925 11985
rect 10869 11939 10925 11951
rect 10955 11939 11009 12023
rect 11039 11957 11117 12023
rect 11039 11939 11073 11957
rect 11065 11923 11073 11939
rect 11107 11923 11117 11957
rect 11065 11911 11117 11923
rect 11147 11957 11203 12041
rect 11147 11923 11157 11957
rect 11191 11923 11203 11957
rect 11147 11911 11203 11923
rect 9381 11345 9433 11427
rect 9381 11311 9389 11345
rect 9423 11311 9433 11345
rect 9381 11297 9433 11311
rect 9463 11367 9517 11427
rect 9463 11333 9473 11367
rect 9507 11333 9517 11367
rect 9463 11297 9517 11333
rect 9547 11345 9601 11427
rect 9547 11311 9557 11345
rect 9591 11311 9601 11345
rect 9547 11297 9601 11311
rect 9631 11297 9685 11427
rect 9715 11347 9869 11427
rect 9715 11313 9725 11347
rect 9759 11313 9825 11347
rect 9859 11313 9869 11347
rect 9715 11297 9869 11313
rect 9899 11418 9963 11427
rect 9899 11384 9915 11418
rect 9949 11384 9963 11418
rect 9899 11350 9963 11384
rect 9899 11316 9915 11350
rect 9949 11316 9963 11350
rect 9899 11297 9963 11316
rect 9699 10665 9751 10683
rect 9503 10627 9559 10665
rect 9503 10593 9515 10627
rect 9549 10593 9559 10627
rect 9503 10581 9559 10593
rect 9589 10581 9643 10665
rect 9673 10599 9751 10665
rect 9673 10581 9707 10599
rect 9699 10565 9707 10581
rect 9741 10565 9751 10599
rect 9699 10553 9751 10565
rect 9781 10599 9837 10683
rect 9781 10565 9791 10599
rect 9825 10565 9837 10599
rect 9781 10553 9837 10565
rect 6186 6537 6238 6553
rect 6186 6503 6194 6537
rect 6228 6503 6238 6537
rect 6186 6469 6238 6503
rect 6186 6435 6194 6469
rect 6228 6435 6238 6469
rect 6186 6423 6238 6435
rect 6268 6537 6320 6553
rect 6268 6503 6278 6537
rect 6312 6503 6320 6537
rect 6268 6469 6320 6503
rect 6268 6435 6278 6469
rect 6312 6435 6320 6469
rect 6268 6423 6320 6435
rect 10080 5873 10132 5921
rect 10080 5839 10088 5873
rect 10122 5839 10132 5873
rect 10080 5791 10132 5839
rect 10162 5913 10231 5921
rect 10162 5879 10187 5913
rect 10221 5879 10231 5913
rect 10162 5837 10231 5879
rect 10261 5837 10327 5921
rect 10357 5837 10399 5921
rect 10429 5901 10495 5921
rect 10429 5867 10439 5901
rect 10473 5867 10495 5901
rect 10429 5837 10495 5867
rect 10525 5896 10584 5921
rect 10525 5862 10540 5896
rect 10574 5862 10584 5896
rect 10525 5837 10584 5862
rect 10614 5913 10668 5921
rect 10614 5879 10624 5913
rect 10658 5879 10668 5913
rect 10614 5837 10668 5879
rect 10698 5896 10752 5921
rect 10698 5862 10708 5896
rect 10742 5862 10752 5896
rect 10698 5837 10752 5862
rect 10782 5904 10834 5921
rect 10782 5870 10792 5904
rect 10826 5870 10834 5904
rect 10782 5837 10834 5870
rect 10888 5896 10940 5921
rect 10888 5862 10896 5896
rect 10930 5862 10940 5896
rect 10888 5837 10940 5862
rect 10970 5913 11024 5921
rect 10970 5879 10980 5913
rect 11014 5879 11024 5913
rect 10970 5837 11024 5879
rect 11054 5896 11108 5921
rect 11054 5862 11064 5896
rect 11098 5862 11108 5896
rect 11054 5837 11108 5862
rect 11138 5896 11192 5921
rect 11138 5862 11148 5896
rect 11182 5862 11192 5896
rect 11138 5837 11192 5862
rect 11222 5837 11282 5921
rect 11312 5909 11381 5921
rect 11312 5875 11337 5909
rect 11371 5875 11381 5909
rect 11312 5837 11381 5875
rect 10162 5791 10214 5837
rect 1898 5453 1950 5501
rect 1898 5419 1906 5453
rect 1940 5419 1950 5453
rect 1898 5371 1950 5419
rect 1980 5493 2049 5501
rect 1980 5459 2005 5493
rect 2039 5459 2049 5493
rect 1980 5417 2049 5459
rect 2079 5417 2145 5501
rect 2175 5417 2217 5501
rect 2247 5481 2313 5501
rect 2247 5447 2257 5481
rect 2291 5447 2313 5481
rect 2247 5417 2313 5447
rect 2343 5476 2402 5501
rect 2343 5442 2358 5476
rect 2392 5442 2402 5476
rect 2343 5417 2402 5442
rect 2432 5493 2486 5501
rect 2432 5459 2442 5493
rect 2476 5459 2486 5493
rect 2432 5417 2486 5459
rect 2516 5476 2570 5501
rect 2516 5442 2526 5476
rect 2560 5442 2570 5476
rect 2516 5417 2570 5442
rect 2600 5484 2652 5501
rect 2600 5450 2610 5484
rect 2644 5450 2652 5484
rect 2600 5417 2652 5450
rect 2706 5476 2758 5501
rect 2706 5442 2714 5476
rect 2748 5442 2758 5476
rect 2706 5417 2758 5442
rect 2788 5493 2842 5501
rect 2788 5459 2798 5493
rect 2832 5459 2842 5493
rect 2788 5417 2842 5459
rect 2872 5476 2926 5501
rect 2872 5442 2882 5476
rect 2916 5442 2926 5476
rect 2872 5417 2926 5442
rect 2956 5476 3010 5501
rect 2956 5442 2966 5476
rect 3000 5442 3010 5476
rect 2956 5417 3010 5442
rect 3040 5417 3100 5501
rect 3130 5489 3199 5501
rect 3130 5455 3155 5489
rect 3189 5455 3199 5489
rect 3130 5417 3199 5455
rect 1980 5371 2032 5417
rect 3147 5371 3199 5417
rect 3229 5453 3281 5501
rect 3229 5419 3239 5453
rect 3273 5419 3281 5453
rect 3229 5371 3281 5419
rect 4032 5445 4084 5493
rect 4032 5411 4040 5445
rect 4074 5411 4084 5445
rect 4032 5363 4084 5411
rect 4114 5485 4183 5493
rect 4114 5451 4139 5485
rect 4173 5451 4183 5485
rect 4114 5409 4183 5451
rect 4213 5409 4279 5493
rect 4309 5409 4351 5493
rect 4381 5473 4447 5493
rect 4381 5439 4391 5473
rect 4425 5439 4447 5473
rect 4381 5409 4447 5439
rect 4477 5468 4536 5493
rect 4477 5434 4492 5468
rect 4526 5434 4536 5468
rect 4477 5409 4536 5434
rect 4566 5485 4620 5493
rect 4566 5451 4576 5485
rect 4610 5451 4620 5485
rect 4566 5409 4620 5451
rect 4650 5468 4704 5493
rect 4650 5434 4660 5468
rect 4694 5434 4704 5468
rect 4650 5409 4704 5434
rect 4734 5476 4786 5493
rect 4734 5442 4744 5476
rect 4778 5442 4786 5476
rect 4734 5409 4786 5442
rect 4840 5468 4892 5493
rect 4840 5434 4848 5468
rect 4882 5434 4892 5468
rect 4840 5409 4892 5434
rect 4922 5485 4976 5493
rect 4922 5451 4932 5485
rect 4966 5451 4976 5485
rect 4922 5409 4976 5451
rect 5006 5468 5060 5493
rect 5006 5434 5016 5468
rect 5050 5434 5060 5468
rect 5006 5409 5060 5434
rect 5090 5468 5144 5493
rect 5090 5434 5100 5468
rect 5134 5434 5144 5468
rect 5090 5409 5144 5434
rect 5174 5409 5234 5493
rect 5264 5481 5333 5493
rect 5264 5447 5289 5481
rect 5323 5447 5333 5481
rect 5264 5409 5333 5447
rect 4114 5363 4166 5409
rect 5281 5363 5333 5409
rect 5363 5445 5415 5493
rect 5363 5411 5373 5445
rect 5407 5411 5415 5445
rect 5363 5363 5415 5411
rect 5984 5445 6036 5493
rect 5984 5411 5992 5445
rect 6026 5411 6036 5445
rect 5984 5363 6036 5411
rect 6066 5485 6135 5493
rect 6066 5451 6091 5485
rect 6125 5451 6135 5485
rect 6066 5409 6135 5451
rect 6165 5409 6231 5493
rect 6261 5409 6303 5493
rect 6333 5473 6399 5493
rect 6333 5439 6343 5473
rect 6377 5439 6399 5473
rect 6333 5409 6399 5439
rect 6429 5468 6488 5493
rect 6429 5434 6444 5468
rect 6478 5434 6488 5468
rect 6429 5409 6488 5434
rect 6518 5485 6572 5493
rect 6518 5451 6528 5485
rect 6562 5451 6572 5485
rect 6518 5409 6572 5451
rect 6602 5468 6656 5493
rect 6602 5434 6612 5468
rect 6646 5434 6656 5468
rect 6602 5409 6656 5434
rect 6686 5476 6738 5493
rect 6686 5442 6696 5476
rect 6730 5442 6738 5476
rect 6686 5409 6738 5442
rect 6792 5468 6844 5493
rect 6792 5434 6800 5468
rect 6834 5434 6844 5468
rect 6792 5409 6844 5434
rect 6874 5485 6928 5493
rect 6874 5451 6884 5485
rect 6918 5451 6928 5485
rect 6874 5409 6928 5451
rect 6958 5468 7012 5493
rect 6958 5434 6968 5468
rect 7002 5434 7012 5468
rect 6958 5409 7012 5434
rect 7042 5468 7096 5493
rect 7042 5434 7052 5468
rect 7086 5434 7096 5468
rect 7042 5409 7096 5434
rect 7126 5409 7186 5493
rect 7216 5481 7285 5493
rect 7216 5447 7241 5481
rect 7275 5447 7285 5481
rect 7216 5409 7285 5447
rect 6066 5363 6118 5409
rect 7233 5363 7285 5409
rect 7315 5445 7367 5493
rect 7315 5411 7325 5445
rect 7359 5411 7367 5445
rect 7315 5363 7367 5411
rect 7986 5451 8038 5499
rect 7986 5417 7994 5451
rect 8028 5417 8038 5451
rect 7986 5369 8038 5417
rect 8068 5491 8137 5499
rect 8068 5457 8093 5491
rect 8127 5457 8137 5491
rect 8068 5415 8137 5457
rect 8167 5415 8233 5499
rect 8263 5415 8305 5499
rect 8335 5479 8401 5499
rect 8335 5445 8345 5479
rect 8379 5445 8401 5479
rect 8335 5415 8401 5445
rect 8431 5474 8490 5499
rect 8431 5440 8446 5474
rect 8480 5440 8490 5474
rect 8431 5415 8490 5440
rect 8520 5491 8574 5499
rect 8520 5457 8530 5491
rect 8564 5457 8574 5491
rect 8520 5415 8574 5457
rect 8604 5474 8658 5499
rect 8604 5440 8614 5474
rect 8648 5440 8658 5474
rect 8604 5415 8658 5440
rect 8688 5482 8740 5499
rect 8688 5448 8698 5482
rect 8732 5448 8740 5482
rect 8688 5415 8740 5448
rect 8794 5474 8846 5499
rect 8794 5440 8802 5474
rect 8836 5440 8846 5474
rect 8794 5415 8846 5440
rect 8876 5491 8930 5499
rect 8876 5457 8886 5491
rect 8920 5457 8930 5491
rect 8876 5415 8930 5457
rect 8960 5474 9014 5499
rect 8960 5440 8970 5474
rect 9004 5440 9014 5474
rect 8960 5415 9014 5440
rect 9044 5474 9098 5499
rect 9044 5440 9054 5474
rect 9088 5440 9098 5474
rect 9044 5415 9098 5440
rect 9128 5415 9188 5499
rect 9218 5487 9287 5499
rect 9218 5453 9243 5487
rect 9277 5453 9287 5487
rect 9218 5415 9287 5453
rect 8068 5369 8120 5415
rect 9235 5369 9287 5415
rect 9317 5451 9369 5499
rect 11329 5791 11381 5837
rect 11411 5873 11463 5921
rect 11411 5839 11421 5873
rect 11455 5839 11463 5873
rect 11411 5791 11463 5839
rect 12142 5861 12194 5909
rect 12142 5827 12150 5861
rect 12184 5827 12194 5861
rect 12142 5779 12194 5827
rect 12224 5901 12293 5909
rect 12224 5867 12249 5901
rect 12283 5867 12293 5901
rect 12224 5825 12293 5867
rect 12323 5825 12389 5909
rect 12419 5825 12461 5909
rect 12491 5889 12557 5909
rect 12491 5855 12501 5889
rect 12535 5855 12557 5889
rect 12491 5825 12557 5855
rect 12587 5884 12646 5909
rect 12587 5850 12602 5884
rect 12636 5850 12646 5884
rect 12587 5825 12646 5850
rect 12676 5901 12730 5909
rect 12676 5867 12686 5901
rect 12720 5867 12730 5901
rect 12676 5825 12730 5867
rect 12760 5884 12814 5909
rect 12760 5850 12770 5884
rect 12804 5850 12814 5884
rect 12760 5825 12814 5850
rect 12844 5892 12896 5909
rect 12844 5858 12854 5892
rect 12888 5858 12896 5892
rect 12844 5825 12896 5858
rect 12950 5884 13002 5909
rect 12950 5850 12958 5884
rect 12992 5850 13002 5884
rect 12950 5825 13002 5850
rect 13032 5901 13086 5909
rect 13032 5867 13042 5901
rect 13076 5867 13086 5901
rect 13032 5825 13086 5867
rect 13116 5884 13170 5909
rect 13116 5850 13126 5884
rect 13160 5850 13170 5884
rect 13116 5825 13170 5850
rect 13200 5884 13254 5909
rect 13200 5850 13210 5884
rect 13244 5850 13254 5884
rect 13200 5825 13254 5850
rect 13284 5825 13344 5909
rect 13374 5897 13443 5909
rect 13374 5863 13399 5897
rect 13433 5863 13443 5897
rect 13374 5825 13443 5863
rect 12224 5779 12276 5825
rect 9317 5417 9327 5451
rect 9361 5417 9369 5451
rect 13391 5779 13443 5825
rect 13473 5861 13525 5909
rect 13473 5827 13483 5861
rect 13517 5827 13525 5861
rect 13473 5779 13525 5827
rect 14100 5869 14152 5917
rect 14100 5835 14108 5869
rect 14142 5835 14152 5869
rect 14100 5787 14152 5835
rect 14182 5909 14251 5917
rect 14182 5875 14207 5909
rect 14241 5875 14251 5909
rect 14182 5833 14251 5875
rect 14281 5833 14347 5917
rect 14377 5833 14419 5917
rect 14449 5897 14515 5917
rect 14449 5863 14459 5897
rect 14493 5863 14515 5897
rect 14449 5833 14515 5863
rect 14545 5892 14604 5917
rect 14545 5858 14560 5892
rect 14594 5858 14604 5892
rect 14545 5833 14604 5858
rect 14634 5909 14688 5917
rect 14634 5875 14644 5909
rect 14678 5875 14688 5909
rect 14634 5833 14688 5875
rect 14718 5892 14772 5917
rect 14718 5858 14728 5892
rect 14762 5858 14772 5892
rect 14718 5833 14772 5858
rect 14802 5900 14854 5917
rect 14802 5866 14812 5900
rect 14846 5866 14854 5900
rect 14802 5833 14854 5866
rect 14908 5892 14960 5917
rect 14908 5858 14916 5892
rect 14950 5858 14960 5892
rect 14908 5833 14960 5858
rect 14990 5909 15044 5917
rect 14990 5875 15000 5909
rect 15034 5875 15044 5909
rect 14990 5833 15044 5875
rect 15074 5892 15128 5917
rect 15074 5858 15084 5892
rect 15118 5858 15128 5892
rect 15074 5833 15128 5858
rect 15158 5892 15212 5917
rect 15158 5858 15168 5892
rect 15202 5858 15212 5892
rect 15158 5833 15212 5858
rect 15242 5833 15302 5917
rect 15332 5905 15401 5917
rect 15332 5871 15357 5905
rect 15391 5871 15401 5905
rect 15332 5833 15401 5871
rect 14182 5787 14234 5833
rect 15349 5787 15401 5833
rect 15431 5869 15483 5917
rect 15431 5835 15441 5869
rect 15475 5835 15483 5869
rect 15431 5787 15483 5835
rect 16094 5875 16146 5923
rect 16094 5841 16102 5875
rect 16136 5841 16146 5875
rect 16094 5793 16146 5841
rect 16176 5915 16245 5923
rect 16176 5881 16201 5915
rect 16235 5881 16245 5915
rect 16176 5839 16245 5881
rect 16275 5839 16341 5923
rect 16371 5839 16413 5923
rect 16443 5903 16509 5923
rect 16443 5869 16453 5903
rect 16487 5869 16509 5903
rect 16443 5839 16509 5869
rect 16539 5898 16598 5923
rect 16539 5864 16554 5898
rect 16588 5864 16598 5898
rect 16539 5839 16598 5864
rect 16628 5915 16682 5923
rect 16628 5881 16638 5915
rect 16672 5881 16682 5915
rect 16628 5839 16682 5881
rect 16712 5898 16766 5923
rect 16712 5864 16722 5898
rect 16756 5864 16766 5898
rect 16712 5839 16766 5864
rect 16796 5906 16848 5923
rect 16796 5872 16806 5906
rect 16840 5872 16848 5906
rect 16796 5839 16848 5872
rect 16902 5898 16954 5923
rect 16902 5864 16910 5898
rect 16944 5864 16954 5898
rect 16902 5839 16954 5864
rect 16984 5915 17038 5923
rect 16984 5881 16994 5915
rect 17028 5881 17038 5915
rect 16984 5839 17038 5881
rect 17068 5898 17122 5923
rect 17068 5864 17078 5898
rect 17112 5864 17122 5898
rect 17068 5839 17122 5864
rect 17152 5898 17206 5923
rect 17152 5864 17162 5898
rect 17196 5864 17206 5898
rect 17152 5839 17206 5864
rect 17236 5839 17296 5923
rect 17326 5911 17395 5923
rect 17326 5877 17351 5911
rect 17385 5877 17395 5911
rect 17326 5839 17395 5877
rect 16176 5793 16228 5839
rect 17343 5793 17395 5839
rect 17425 5875 17477 5923
rect 17425 5841 17435 5875
rect 17469 5841 17477 5875
rect 17425 5793 17477 5841
rect 9317 5369 9369 5417
rect 10108 4999 10160 5047
rect 10108 4965 10116 4999
rect 10150 4965 10160 4999
rect 10108 4917 10160 4965
rect 10190 5039 10259 5047
rect 10190 5005 10215 5039
rect 10249 5005 10259 5039
rect 10190 4963 10259 5005
rect 10289 4963 10355 5047
rect 10385 4963 10427 5047
rect 10457 5027 10523 5047
rect 10457 4993 10467 5027
rect 10501 4993 10523 5027
rect 10457 4963 10523 4993
rect 10553 5022 10612 5047
rect 10553 4988 10568 5022
rect 10602 4988 10612 5022
rect 10553 4963 10612 4988
rect 10642 5039 10696 5047
rect 10642 5005 10652 5039
rect 10686 5005 10696 5039
rect 10642 4963 10696 5005
rect 10726 5022 10780 5047
rect 10726 4988 10736 5022
rect 10770 4988 10780 5022
rect 10726 4963 10780 4988
rect 10810 5030 10862 5047
rect 10810 4996 10820 5030
rect 10854 4996 10862 5030
rect 10810 4963 10862 4996
rect 10916 5022 10968 5047
rect 10916 4988 10924 5022
rect 10958 4988 10968 5022
rect 10916 4963 10968 4988
rect 10998 5039 11052 5047
rect 10998 5005 11008 5039
rect 11042 5005 11052 5039
rect 10998 4963 11052 5005
rect 11082 5022 11136 5047
rect 11082 4988 11092 5022
rect 11126 4988 11136 5022
rect 11082 4963 11136 4988
rect 11166 5022 11220 5047
rect 11166 4988 11176 5022
rect 11210 4988 11220 5022
rect 11166 4963 11220 4988
rect 11250 4963 11310 5047
rect 11340 5035 11409 5047
rect 11340 5001 11365 5035
rect 11399 5001 11409 5035
rect 11340 4963 11409 5001
rect 10190 4917 10242 4963
rect 11357 4917 11409 4963
rect 11439 4999 11491 5047
rect 11439 4965 11449 4999
rect 11483 4965 11491 4999
rect 11439 4917 11491 4965
rect 12378 4955 12430 5003
rect 12378 4921 12386 4955
rect 12420 4921 12430 4955
rect 12378 4873 12430 4921
rect 12460 4995 12529 5003
rect 12460 4961 12485 4995
rect 12519 4961 12529 4995
rect 12460 4919 12529 4961
rect 12559 4919 12625 5003
rect 12655 4919 12697 5003
rect 12727 4983 12793 5003
rect 12727 4949 12737 4983
rect 12771 4949 12793 4983
rect 12727 4919 12793 4949
rect 12823 4978 12882 5003
rect 12823 4944 12838 4978
rect 12872 4944 12882 4978
rect 12823 4919 12882 4944
rect 12912 4995 12966 5003
rect 12912 4961 12922 4995
rect 12956 4961 12966 4995
rect 12912 4919 12966 4961
rect 12996 4978 13050 5003
rect 12996 4944 13006 4978
rect 13040 4944 13050 4978
rect 12996 4919 13050 4944
rect 13080 4986 13132 5003
rect 13080 4952 13090 4986
rect 13124 4952 13132 4986
rect 13080 4919 13132 4952
rect 13186 4978 13238 5003
rect 13186 4944 13194 4978
rect 13228 4944 13238 4978
rect 13186 4919 13238 4944
rect 13268 4995 13322 5003
rect 13268 4961 13278 4995
rect 13312 4961 13322 4995
rect 13268 4919 13322 4961
rect 13352 4978 13406 5003
rect 13352 4944 13362 4978
rect 13396 4944 13406 4978
rect 13352 4919 13406 4944
rect 13436 4978 13490 5003
rect 13436 4944 13446 4978
rect 13480 4944 13490 4978
rect 13436 4919 13490 4944
rect 13520 4919 13580 5003
rect 13610 4991 13679 5003
rect 13610 4957 13635 4991
rect 13669 4957 13679 4991
rect 13610 4919 13679 4957
rect 12460 4873 12512 4919
rect 13627 4873 13679 4919
rect 13709 4955 13761 5003
rect 13709 4921 13719 4955
rect 13753 4921 13761 4955
rect 13709 4873 13761 4921
rect 14380 4949 14432 4997
rect 14380 4915 14388 4949
rect 14422 4915 14432 4949
rect 14380 4867 14432 4915
rect 14462 4989 14531 4997
rect 14462 4955 14487 4989
rect 14521 4955 14531 4989
rect 14462 4913 14531 4955
rect 14561 4913 14627 4997
rect 14657 4913 14699 4997
rect 14729 4977 14795 4997
rect 14729 4943 14739 4977
rect 14773 4943 14795 4977
rect 14729 4913 14795 4943
rect 14825 4972 14884 4997
rect 14825 4938 14840 4972
rect 14874 4938 14884 4972
rect 14825 4913 14884 4938
rect 14914 4989 14968 4997
rect 14914 4955 14924 4989
rect 14958 4955 14968 4989
rect 14914 4913 14968 4955
rect 14998 4972 15052 4997
rect 14998 4938 15008 4972
rect 15042 4938 15052 4972
rect 14998 4913 15052 4938
rect 15082 4980 15134 4997
rect 15082 4946 15092 4980
rect 15126 4946 15134 4980
rect 15082 4913 15134 4946
rect 15188 4972 15240 4997
rect 15188 4938 15196 4972
rect 15230 4938 15240 4972
rect 15188 4913 15240 4938
rect 15270 4989 15324 4997
rect 15270 4955 15280 4989
rect 15314 4955 15324 4989
rect 15270 4913 15324 4955
rect 15354 4972 15408 4997
rect 15354 4938 15364 4972
rect 15398 4938 15408 4972
rect 15354 4913 15408 4938
rect 15438 4972 15492 4997
rect 15438 4938 15448 4972
rect 15482 4938 15492 4972
rect 15438 4913 15492 4938
rect 15522 4913 15582 4997
rect 15612 4985 15681 4997
rect 15612 4951 15637 4985
rect 15671 4951 15681 4985
rect 15612 4913 15681 4951
rect 14462 4867 14514 4913
rect 15629 4867 15681 4913
rect 15711 4949 15763 4997
rect 15711 4915 15721 4949
rect 15755 4915 15763 4949
rect 15711 4867 15763 4915
rect 16402 4931 16454 4979
rect 16402 4897 16410 4931
rect 16444 4897 16454 4931
rect 16402 4849 16454 4897
rect 16484 4971 16553 4979
rect 16484 4937 16509 4971
rect 16543 4937 16553 4971
rect 16484 4895 16553 4937
rect 16583 4895 16649 4979
rect 16679 4895 16721 4979
rect 16751 4959 16817 4979
rect 16751 4925 16761 4959
rect 16795 4925 16817 4959
rect 16751 4895 16817 4925
rect 16847 4954 16906 4979
rect 16847 4920 16862 4954
rect 16896 4920 16906 4954
rect 16847 4895 16906 4920
rect 16936 4971 16990 4979
rect 16936 4937 16946 4971
rect 16980 4937 16990 4971
rect 16936 4895 16990 4937
rect 17020 4954 17074 4979
rect 17020 4920 17030 4954
rect 17064 4920 17074 4954
rect 17020 4895 17074 4920
rect 17104 4962 17156 4979
rect 17104 4928 17114 4962
rect 17148 4928 17156 4962
rect 17104 4895 17156 4928
rect 17210 4954 17262 4979
rect 17210 4920 17218 4954
rect 17252 4920 17262 4954
rect 17210 4895 17262 4920
rect 17292 4971 17346 4979
rect 17292 4937 17302 4971
rect 17336 4937 17346 4971
rect 17292 4895 17346 4937
rect 17376 4954 17430 4979
rect 17376 4920 17386 4954
rect 17420 4920 17430 4954
rect 17376 4895 17430 4920
rect 17460 4954 17514 4979
rect 17460 4920 17470 4954
rect 17504 4920 17514 4954
rect 17460 4895 17514 4920
rect 17544 4895 17604 4979
rect 17634 4967 17703 4979
rect 17634 4933 17659 4967
rect 17693 4933 17703 4967
rect 17634 4895 17703 4933
rect 16484 4849 16536 4895
rect 17651 4849 17703 4895
rect 17733 4931 17785 4979
rect 17733 4897 17743 4931
rect 17777 4897 17785 4931
rect 17733 4849 17785 4897
rect 1868 2193 1920 2241
rect 1868 2159 1876 2193
rect 1910 2159 1920 2193
rect 1868 2111 1920 2159
rect 1950 2233 2019 2241
rect 1950 2199 1975 2233
rect 2009 2199 2019 2233
rect 1950 2157 2019 2199
rect 2049 2157 2115 2241
rect 2145 2157 2187 2241
rect 2217 2221 2283 2241
rect 2217 2187 2227 2221
rect 2261 2187 2283 2221
rect 2217 2157 2283 2187
rect 2313 2216 2372 2241
rect 2313 2182 2328 2216
rect 2362 2182 2372 2216
rect 2313 2157 2372 2182
rect 2402 2233 2456 2241
rect 2402 2199 2412 2233
rect 2446 2199 2456 2233
rect 2402 2157 2456 2199
rect 2486 2216 2540 2241
rect 2486 2182 2496 2216
rect 2530 2182 2540 2216
rect 2486 2157 2540 2182
rect 2570 2224 2622 2241
rect 2570 2190 2580 2224
rect 2614 2190 2622 2224
rect 2570 2157 2622 2190
rect 2676 2216 2728 2241
rect 2676 2182 2684 2216
rect 2718 2182 2728 2216
rect 2676 2157 2728 2182
rect 2758 2233 2812 2241
rect 2758 2199 2768 2233
rect 2802 2199 2812 2233
rect 2758 2157 2812 2199
rect 2842 2216 2896 2241
rect 2842 2182 2852 2216
rect 2886 2182 2896 2216
rect 2842 2157 2896 2182
rect 2926 2216 2980 2241
rect 2926 2182 2936 2216
rect 2970 2182 2980 2216
rect 2926 2157 2980 2182
rect 3010 2157 3070 2241
rect 3100 2229 3169 2241
rect 3100 2195 3125 2229
rect 3159 2195 3169 2229
rect 3100 2157 3169 2195
rect 1950 2111 2002 2157
rect 3117 2111 3169 2157
rect 3199 2193 3251 2241
rect 3199 2159 3209 2193
rect 3243 2159 3251 2193
rect 3199 2111 3251 2159
rect 3938 2189 3990 2237
rect 3938 2155 3946 2189
rect 3980 2155 3990 2189
rect 3938 2107 3990 2155
rect 4020 2229 4089 2237
rect 4020 2195 4045 2229
rect 4079 2195 4089 2229
rect 4020 2153 4089 2195
rect 4119 2153 4185 2237
rect 4215 2153 4257 2237
rect 4287 2217 4353 2237
rect 4287 2183 4297 2217
rect 4331 2183 4353 2217
rect 4287 2153 4353 2183
rect 4383 2212 4442 2237
rect 4383 2178 4398 2212
rect 4432 2178 4442 2212
rect 4383 2153 4442 2178
rect 4472 2229 4526 2237
rect 4472 2195 4482 2229
rect 4516 2195 4526 2229
rect 4472 2153 4526 2195
rect 4556 2212 4610 2237
rect 4556 2178 4566 2212
rect 4600 2178 4610 2212
rect 4556 2153 4610 2178
rect 4640 2220 4692 2237
rect 4640 2186 4650 2220
rect 4684 2186 4692 2220
rect 4640 2153 4692 2186
rect 4746 2212 4798 2237
rect 4746 2178 4754 2212
rect 4788 2178 4798 2212
rect 4746 2153 4798 2178
rect 4828 2229 4882 2237
rect 4828 2195 4838 2229
rect 4872 2195 4882 2229
rect 4828 2153 4882 2195
rect 4912 2212 4966 2237
rect 4912 2178 4922 2212
rect 4956 2178 4966 2212
rect 4912 2153 4966 2178
rect 4996 2212 5050 2237
rect 4996 2178 5006 2212
rect 5040 2178 5050 2212
rect 4996 2153 5050 2178
rect 5080 2153 5140 2237
rect 5170 2225 5239 2237
rect 5170 2191 5195 2225
rect 5229 2191 5239 2225
rect 5170 2153 5239 2191
rect 4020 2107 4072 2153
rect 5187 2107 5239 2153
rect 5269 2189 5321 2237
rect 5269 2155 5279 2189
rect 5313 2155 5321 2189
rect 5269 2107 5321 2155
rect 5890 2189 5942 2237
rect 5890 2155 5898 2189
rect 5932 2155 5942 2189
rect 5890 2107 5942 2155
rect 5972 2229 6041 2237
rect 5972 2195 5997 2229
rect 6031 2195 6041 2229
rect 5972 2153 6041 2195
rect 6071 2153 6137 2237
rect 6167 2153 6209 2237
rect 6239 2217 6305 2237
rect 6239 2183 6249 2217
rect 6283 2183 6305 2217
rect 6239 2153 6305 2183
rect 6335 2212 6394 2237
rect 6335 2178 6350 2212
rect 6384 2178 6394 2212
rect 6335 2153 6394 2178
rect 6424 2229 6478 2237
rect 6424 2195 6434 2229
rect 6468 2195 6478 2229
rect 6424 2153 6478 2195
rect 6508 2212 6562 2237
rect 6508 2178 6518 2212
rect 6552 2178 6562 2212
rect 6508 2153 6562 2178
rect 6592 2220 6644 2237
rect 6592 2186 6602 2220
rect 6636 2186 6644 2220
rect 6592 2153 6644 2186
rect 6698 2212 6750 2237
rect 6698 2178 6706 2212
rect 6740 2178 6750 2212
rect 6698 2153 6750 2178
rect 6780 2229 6834 2237
rect 6780 2195 6790 2229
rect 6824 2195 6834 2229
rect 6780 2153 6834 2195
rect 6864 2212 6918 2237
rect 6864 2178 6874 2212
rect 6908 2178 6918 2212
rect 6864 2153 6918 2178
rect 6948 2212 7002 2237
rect 6948 2178 6958 2212
rect 6992 2178 7002 2212
rect 6948 2153 7002 2178
rect 7032 2153 7092 2237
rect 7122 2225 7191 2237
rect 7122 2191 7147 2225
rect 7181 2191 7191 2225
rect 7122 2153 7191 2191
rect 5972 2107 6024 2153
rect 7139 2107 7191 2153
rect 7221 2189 7273 2237
rect 7221 2155 7231 2189
rect 7265 2155 7273 2189
rect 7221 2107 7273 2155
rect 7892 2195 7944 2243
rect 7892 2161 7900 2195
rect 7934 2161 7944 2195
rect 7892 2113 7944 2161
rect 7974 2235 8043 2243
rect 7974 2201 7999 2235
rect 8033 2201 8043 2235
rect 7974 2159 8043 2201
rect 8073 2159 8139 2243
rect 8169 2159 8211 2243
rect 8241 2223 8307 2243
rect 8241 2189 8251 2223
rect 8285 2189 8307 2223
rect 8241 2159 8307 2189
rect 8337 2218 8396 2243
rect 8337 2184 8352 2218
rect 8386 2184 8396 2218
rect 8337 2159 8396 2184
rect 8426 2235 8480 2243
rect 8426 2201 8436 2235
rect 8470 2201 8480 2235
rect 8426 2159 8480 2201
rect 8510 2218 8564 2243
rect 8510 2184 8520 2218
rect 8554 2184 8564 2218
rect 8510 2159 8564 2184
rect 8594 2226 8646 2243
rect 8594 2192 8604 2226
rect 8638 2192 8646 2226
rect 8594 2159 8646 2192
rect 8700 2218 8752 2243
rect 8700 2184 8708 2218
rect 8742 2184 8752 2218
rect 8700 2159 8752 2184
rect 8782 2235 8836 2243
rect 8782 2201 8792 2235
rect 8826 2201 8836 2235
rect 8782 2159 8836 2201
rect 8866 2218 8920 2243
rect 8866 2184 8876 2218
rect 8910 2184 8920 2218
rect 8866 2159 8920 2184
rect 8950 2218 9004 2243
rect 8950 2184 8960 2218
rect 8994 2184 9004 2218
rect 8950 2159 9004 2184
rect 9034 2159 9094 2243
rect 9124 2231 9193 2243
rect 9124 2197 9149 2231
rect 9183 2197 9193 2231
rect 9124 2159 9193 2197
rect 7974 2113 8026 2159
rect 9141 2113 9193 2159
rect 9223 2195 9275 2243
rect 9223 2161 9233 2195
rect 9267 2161 9275 2195
rect 9223 2113 9275 2161
rect 9844 2195 9896 2243
rect 9844 2161 9852 2195
rect 9886 2161 9896 2195
rect 9844 2113 9896 2161
rect 9926 2235 9995 2243
rect 9926 2201 9951 2235
rect 9985 2201 9995 2235
rect 9926 2159 9995 2201
rect 10025 2159 10091 2243
rect 10121 2159 10163 2243
rect 10193 2223 10259 2243
rect 10193 2189 10203 2223
rect 10237 2189 10259 2223
rect 10193 2159 10259 2189
rect 10289 2218 10348 2243
rect 10289 2184 10304 2218
rect 10338 2184 10348 2218
rect 10289 2159 10348 2184
rect 10378 2235 10432 2243
rect 10378 2201 10388 2235
rect 10422 2201 10432 2235
rect 10378 2159 10432 2201
rect 10462 2218 10516 2243
rect 10462 2184 10472 2218
rect 10506 2184 10516 2218
rect 10462 2159 10516 2184
rect 10546 2226 10598 2243
rect 10546 2192 10556 2226
rect 10590 2192 10598 2226
rect 10546 2159 10598 2192
rect 10652 2218 10704 2243
rect 10652 2184 10660 2218
rect 10694 2184 10704 2218
rect 10652 2159 10704 2184
rect 10734 2235 10788 2243
rect 10734 2201 10744 2235
rect 10778 2201 10788 2235
rect 10734 2159 10788 2201
rect 10818 2218 10872 2243
rect 10818 2184 10828 2218
rect 10862 2184 10872 2218
rect 10818 2159 10872 2184
rect 10902 2218 10956 2243
rect 10902 2184 10912 2218
rect 10946 2184 10956 2218
rect 10902 2159 10956 2184
rect 10986 2159 11046 2243
rect 11076 2231 11145 2243
rect 11076 2197 11101 2231
rect 11135 2197 11145 2231
rect 11076 2159 11145 2197
rect 9926 2113 9978 2159
rect 11093 2113 11145 2159
rect 11175 2195 11227 2243
rect 11175 2161 11185 2195
rect 11219 2161 11227 2195
rect 11175 2113 11227 2161
rect 11836 2195 11888 2243
rect 11836 2161 11844 2195
rect 11878 2161 11888 2195
rect 11836 2113 11888 2161
rect 11918 2235 11987 2243
rect 11918 2201 11943 2235
rect 11977 2201 11987 2235
rect 11918 2159 11987 2201
rect 12017 2159 12083 2243
rect 12113 2159 12155 2243
rect 12185 2223 12251 2243
rect 12185 2189 12195 2223
rect 12229 2189 12251 2223
rect 12185 2159 12251 2189
rect 12281 2218 12340 2243
rect 12281 2184 12296 2218
rect 12330 2184 12340 2218
rect 12281 2159 12340 2184
rect 12370 2235 12424 2243
rect 12370 2201 12380 2235
rect 12414 2201 12424 2235
rect 12370 2159 12424 2201
rect 12454 2218 12508 2243
rect 12454 2184 12464 2218
rect 12498 2184 12508 2218
rect 12454 2159 12508 2184
rect 12538 2226 12590 2243
rect 12538 2192 12548 2226
rect 12582 2192 12590 2226
rect 12538 2159 12590 2192
rect 12644 2218 12696 2243
rect 12644 2184 12652 2218
rect 12686 2184 12696 2218
rect 12644 2159 12696 2184
rect 12726 2235 12780 2243
rect 12726 2201 12736 2235
rect 12770 2201 12780 2235
rect 12726 2159 12780 2201
rect 12810 2218 12864 2243
rect 12810 2184 12820 2218
rect 12854 2184 12864 2218
rect 12810 2159 12864 2184
rect 12894 2218 12948 2243
rect 12894 2184 12904 2218
rect 12938 2184 12948 2218
rect 12894 2159 12948 2184
rect 12978 2159 13038 2243
rect 13068 2231 13137 2243
rect 13068 2197 13093 2231
rect 13127 2197 13137 2231
rect 13068 2159 13137 2197
rect 11918 2113 11970 2159
rect 13085 2113 13137 2159
rect 13167 2195 13219 2243
rect 13167 2161 13177 2195
rect 13211 2161 13219 2195
rect 13167 2113 13219 2161
rect 13788 2195 13840 2243
rect 13788 2161 13796 2195
rect 13830 2161 13840 2195
rect 13788 2113 13840 2161
rect 13870 2235 13939 2243
rect 13870 2201 13895 2235
rect 13929 2201 13939 2235
rect 13870 2159 13939 2201
rect 13969 2159 14035 2243
rect 14065 2159 14107 2243
rect 14137 2223 14203 2243
rect 14137 2189 14147 2223
rect 14181 2189 14203 2223
rect 14137 2159 14203 2189
rect 14233 2218 14292 2243
rect 14233 2184 14248 2218
rect 14282 2184 14292 2218
rect 14233 2159 14292 2184
rect 14322 2235 14376 2243
rect 14322 2201 14332 2235
rect 14366 2201 14376 2235
rect 14322 2159 14376 2201
rect 14406 2218 14460 2243
rect 14406 2184 14416 2218
rect 14450 2184 14460 2218
rect 14406 2159 14460 2184
rect 14490 2226 14542 2243
rect 14490 2192 14500 2226
rect 14534 2192 14542 2226
rect 14490 2159 14542 2192
rect 14596 2218 14648 2243
rect 14596 2184 14604 2218
rect 14638 2184 14648 2218
rect 14596 2159 14648 2184
rect 14678 2235 14732 2243
rect 14678 2201 14688 2235
rect 14722 2201 14732 2235
rect 14678 2159 14732 2201
rect 14762 2218 14816 2243
rect 14762 2184 14772 2218
rect 14806 2184 14816 2218
rect 14762 2159 14816 2184
rect 14846 2218 14900 2243
rect 14846 2184 14856 2218
rect 14890 2184 14900 2218
rect 14846 2159 14900 2184
rect 14930 2159 14990 2243
rect 15020 2231 15089 2243
rect 15020 2197 15045 2231
rect 15079 2197 15089 2231
rect 15020 2159 15089 2197
rect 13870 2113 13922 2159
rect 15037 2113 15089 2159
rect 15119 2195 15171 2243
rect 15119 2161 15129 2195
rect 15163 2161 15171 2195
rect 15119 2113 15171 2161
rect 15852 2195 15904 2243
rect 15852 2161 15860 2195
rect 15894 2161 15904 2195
rect 15852 2113 15904 2161
rect 15934 2235 16003 2243
rect 15934 2201 15959 2235
rect 15993 2201 16003 2235
rect 15934 2159 16003 2201
rect 16033 2159 16099 2243
rect 16129 2159 16171 2243
rect 16201 2223 16267 2243
rect 16201 2189 16211 2223
rect 16245 2189 16267 2223
rect 16201 2159 16267 2189
rect 16297 2218 16356 2243
rect 16297 2184 16312 2218
rect 16346 2184 16356 2218
rect 16297 2159 16356 2184
rect 16386 2235 16440 2243
rect 16386 2201 16396 2235
rect 16430 2201 16440 2235
rect 16386 2159 16440 2201
rect 16470 2218 16524 2243
rect 16470 2184 16480 2218
rect 16514 2184 16524 2218
rect 16470 2159 16524 2184
rect 16554 2226 16606 2243
rect 16554 2192 16564 2226
rect 16598 2192 16606 2226
rect 16554 2159 16606 2192
rect 16660 2218 16712 2243
rect 16660 2184 16668 2218
rect 16702 2184 16712 2218
rect 16660 2159 16712 2184
rect 16742 2235 16796 2243
rect 16742 2201 16752 2235
rect 16786 2201 16796 2235
rect 16742 2159 16796 2201
rect 16826 2218 16880 2243
rect 16826 2184 16836 2218
rect 16870 2184 16880 2218
rect 16826 2159 16880 2184
rect 16910 2218 16964 2243
rect 16910 2184 16920 2218
rect 16954 2184 16964 2218
rect 16910 2159 16964 2184
rect 16994 2159 17054 2243
rect 17084 2231 17153 2243
rect 17084 2197 17109 2231
rect 17143 2197 17153 2231
rect 17084 2159 17153 2197
rect 15934 2113 15986 2159
rect 17101 2113 17153 2159
rect 17183 2195 17235 2243
rect 17183 2161 17193 2195
rect 17227 2161 17235 2195
rect 17183 2113 17235 2161
<< pdiff >>
rect 18513 35099 18713 35107
rect 18513 35065 18525 35099
rect 18559 35065 18596 35099
rect 18630 35065 18667 35099
rect 18701 35065 18713 35099
rect 18513 35055 18713 35065
rect 18513 35015 18713 35025
rect 18513 34981 18525 35015
rect 18559 34981 18593 35015
rect 18627 34981 18661 35015
rect 18695 34981 18713 35015
rect 18513 34973 18713 34981
rect 18513 34958 18641 34973
rect 18513 34918 18641 34928
rect 18513 34884 18525 34918
rect 18559 34884 18593 34918
rect 18627 34884 18641 34918
rect 18513 34876 18641 34884
rect 18513 34814 18713 34822
rect 18513 34780 18531 34814
rect 18565 34780 18599 34814
rect 18633 34780 18667 34814
rect 18701 34780 18713 34814
rect 18513 34770 18713 34780
rect 18513 34730 18713 34740
rect 18513 34696 18555 34730
rect 18589 34696 18635 34730
rect 18669 34696 18713 34730
rect 18513 34686 18713 34696
rect 18513 34644 18713 34656
rect 18513 34610 18525 34644
rect 18559 34610 18596 34644
rect 18630 34610 18667 34644
rect 18701 34610 18713 34644
rect 18513 34602 18713 34610
rect 18513 34520 18597 34528
rect 18513 34486 18533 34520
rect 18567 34486 18597 34520
rect 18513 34475 18597 34486
rect 18513 34361 18597 34445
rect 18513 34321 18597 34331
rect 18513 34287 18543 34321
rect 18577 34287 18597 34321
rect 18513 34277 18597 34287
rect 18513 34232 18597 34247
rect 18513 34226 18663 34232
rect 18513 34192 18533 34226
rect 18567 34192 18663 34226
rect 18513 34182 18663 34192
rect 18513 34142 18663 34152
rect 18513 34108 18525 34142
rect 18559 34108 18593 34142
rect 18627 34108 18663 34142
rect 18513 34065 18663 34108
rect 18513 34050 18597 34065
rect 18513 33947 18597 34020
rect 18513 33903 18597 33917
rect 18513 33869 18538 33903
rect 18572 33869 18597 33903
rect 18513 33852 18597 33869
rect 18513 33811 18597 33822
rect 18513 33777 18533 33811
rect 18567 33777 18597 33811
rect 18513 33767 18597 33777
rect 18513 33727 18597 33737
rect 18513 33693 18525 33727
rect 18559 33693 18597 33727
rect 18513 33685 18597 33693
rect 18519 33623 18647 33631
rect 18519 33589 18533 33623
rect 18567 33589 18601 33623
rect 18635 33589 18647 33623
rect 18519 33579 18647 33589
rect 18519 33539 18647 33549
rect 18519 33505 18549 33539
rect 18583 33505 18647 33539
rect 18519 33495 18647 33505
rect 18519 33455 18647 33465
rect 18519 33421 18533 33455
rect 18567 33421 18601 33455
rect 18635 33421 18647 33455
rect 18519 33413 18647 33421
rect 18521 32793 18721 32801
rect 18521 32759 18533 32793
rect 18567 32759 18604 32793
rect 18638 32759 18675 32793
rect 18709 32759 18721 32793
rect 18521 32749 18721 32759
rect 18521 32709 18721 32719
rect 18521 32675 18533 32709
rect 18567 32675 18601 32709
rect 18635 32675 18669 32709
rect 18703 32675 18721 32709
rect 18521 32667 18721 32675
rect 18521 32652 18649 32667
rect 18521 32612 18649 32622
rect 18521 32578 18533 32612
rect 18567 32578 18601 32612
rect 18635 32578 18649 32612
rect 18521 32570 18649 32578
rect 18521 32508 18721 32516
rect 18521 32474 18539 32508
rect 18573 32474 18607 32508
rect 18641 32474 18675 32508
rect 18709 32474 18721 32508
rect 18521 32464 18721 32474
rect 18521 32424 18721 32434
rect 18521 32390 18563 32424
rect 18597 32390 18643 32424
rect 18677 32390 18721 32424
rect 18521 32380 18721 32390
rect 18521 32338 18721 32350
rect 18521 32304 18533 32338
rect 18567 32304 18604 32338
rect 18638 32304 18675 32338
rect 18709 32304 18721 32338
rect 18521 32296 18721 32304
rect 18521 32214 18605 32222
rect 18521 32180 18541 32214
rect 18575 32180 18605 32214
rect 18521 32169 18605 32180
rect 18521 32055 18605 32139
rect 18521 32015 18605 32025
rect 18521 31981 18551 32015
rect 18585 31981 18605 32015
rect 18521 31971 18605 31981
rect 18521 31926 18605 31941
rect 18521 31920 18671 31926
rect 18521 31886 18541 31920
rect 18575 31886 18671 31920
rect 18521 31876 18671 31886
rect 18521 31836 18671 31846
rect 18521 31802 18533 31836
rect 18567 31802 18601 31836
rect 18635 31802 18671 31836
rect 18521 31759 18671 31802
rect 18521 31744 18605 31759
rect 18521 31641 18605 31714
rect 18521 31597 18605 31611
rect 18521 31563 18546 31597
rect 18580 31563 18605 31597
rect 18521 31546 18605 31563
rect 18521 31505 18605 31516
rect 18521 31471 18541 31505
rect 18575 31471 18605 31505
rect 18521 31461 18605 31471
rect 18521 31421 18605 31431
rect 18521 31387 18533 31421
rect 18567 31387 18605 31421
rect 18521 31379 18605 31387
rect 18527 31317 18655 31325
rect 18527 31283 18541 31317
rect 18575 31283 18609 31317
rect 18643 31283 18655 31317
rect 18527 31273 18655 31283
rect 18527 31233 18655 31243
rect 18527 31199 18557 31233
rect 18591 31199 18655 31233
rect 18527 31189 18655 31199
rect 18527 31149 18655 31159
rect 18527 31115 18541 31149
rect 18575 31115 18609 31149
rect 18643 31115 18655 31149
rect 18527 31107 18655 31115
rect 18529 30579 18729 30587
rect 18529 30545 18541 30579
rect 18575 30545 18612 30579
rect 18646 30545 18683 30579
rect 18717 30545 18729 30579
rect 18529 30535 18729 30545
rect 18529 30495 18729 30505
rect 18529 30461 18541 30495
rect 18575 30461 18609 30495
rect 18643 30461 18677 30495
rect 18711 30461 18729 30495
rect 18529 30453 18729 30461
rect 18529 30438 18657 30453
rect 18529 30398 18657 30408
rect 18529 30364 18541 30398
rect 18575 30364 18609 30398
rect 18643 30364 18657 30398
rect 18529 30356 18657 30364
rect 18529 30294 18729 30302
rect 18529 30260 18547 30294
rect 18581 30260 18615 30294
rect 18649 30260 18683 30294
rect 18717 30260 18729 30294
rect 18529 30250 18729 30260
rect 18529 30210 18729 30220
rect 18529 30176 18571 30210
rect 18605 30176 18651 30210
rect 18685 30176 18729 30210
rect 18529 30166 18729 30176
rect 18529 30124 18729 30136
rect 18529 30090 18541 30124
rect 18575 30090 18612 30124
rect 18646 30090 18683 30124
rect 18717 30090 18729 30124
rect 18529 30082 18729 30090
rect 18529 30000 18613 30008
rect 18529 29966 18549 30000
rect 18583 29966 18613 30000
rect 18529 29955 18613 29966
rect 18529 29841 18613 29925
rect 18529 29801 18613 29811
rect 18529 29767 18559 29801
rect 18593 29767 18613 29801
rect 18529 29757 18613 29767
rect 18529 29712 18613 29727
rect 18529 29706 18679 29712
rect 18529 29672 18549 29706
rect 18583 29672 18679 29706
rect 18529 29662 18679 29672
rect 18529 29622 18679 29632
rect 18529 29588 18541 29622
rect 18575 29588 18609 29622
rect 18643 29588 18679 29622
rect 18529 29545 18679 29588
rect 18529 29530 18613 29545
rect 18529 29427 18613 29500
rect 18529 29383 18613 29397
rect 18529 29349 18554 29383
rect 18588 29349 18613 29383
rect 18529 29332 18613 29349
rect 18529 29291 18613 29302
rect 18529 29257 18549 29291
rect 18583 29257 18613 29291
rect 18529 29247 18613 29257
rect 18529 29207 18613 29217
rect 18529 29173 18541 29207
rect 18575 29173 18613 29207
rect 18529 29165 18613 29173
rect 18535 29103 18663 29111
rect 18535 29069 18549 29103
rect 18583 29069 18617 29103
rect 18651 29069 18663 29103
rect 18535 29059 18663 29069
rect 18535 29019 18663 29029
rect 18535 28985 18565 29019
rect 18599 28985 18663 29019
rect 18535 28975 18663 28985
rect 18535 28935 18663 28945
rect 18535 28901 18549 28935
rect 18583 28901 18617 28935
rect 18651 28901 18663 28935
rect 18535 28893 18663 28901
rect 18511 28379 18711 28387
rect 18511 28345 18523 28379
rect 18557 28345 18594 28379
rect 18628 28345 18665 28379
rect 18699 28345 18711 28379
rect 18511 28335 18711 28345
rect 18511 28295 18711 28305
rect 18511 28261 18523 28295
rect 18557 28261 18591 28295
rect 18625 28261 18659 28295
rect 18693 28261 18711 28295
rect 18511 28253 18711 28261
rect 18511 28238 18639 28253
rect 18511 28198 18639 28208
rect 18511 28164 18523 28198
rect 18557 28164 18591 28198
rect 18625 28164 18639 28198
rect 18511 28156 18639 28164
rect 18511 28094 18711 28102
rect 18511 28060 18529 28094
rect 18563 28060 18597 28094
rect 18631 28060 18665 28094
rect 18699 28060 18711 28094
rect 18511 28050 18711 28060
rect 18511 28010 18711 28020
rect 18511 27976 18553 28010
rect 18587 27976 18633 28010
rect 18667 27976 18711 28010
rect 18511 27966 18711 27976
rect 18511 27924 18711 27936
rect 18511 27890 18523 27924
rect 18557 27890 18594 27924
rect 18628 27890 18665 27924
rect 18699 27890 18711 27924
rect 18511 27882 18711 27890
rect 18511 27800 18595 27808
rect 18511 27766 18531 27800
rect 18565 27766 18595 27800
rect 18511 27755 18595 27766
rect 18511 27641 18595 27725
rect 18511 27601 18595 27611
rect 18511 27567 18541 27601
rect 18575 27567 18595 27601
rect 18511 27557 18595 27567
rect 18511 27512 18595 27527
rect 18511 27506 18661 27512
rect 18511 27472 18531 27506
rect 18565 27472 18661 27506
rect 18511 27462 18661 27472
rect 18511 27422 18661 27432
rect 18511 27388 18523 27422
rect 18557 27388 18591 27422
rect 18625 27388 18661 27422
rect 18511 27345 18661 27388
rect 18511 27330 18595 27345
rect 18511 27227 18595 27300
rect 18511 27183 18595 27197
rect 18511 27149 18536 27183
rect 18570 27149 18595 27183
rect 18511 27132 18595 27149
rect 18511 27091 18595 27102
rect 18511 27057 18531 27091
rect 18565 27057 18595 27091
rect 18511 27047 18595 27057
rect 18511 27007 18595 27017
rect 18511 26973 18523 27007
rect 18557 26973 18595 27007
rect 18511 26965 18595 26973
rect 18517 26903 18645 26911
rect 18517 26869 18531 26903
rect 18565 26869 18599 26903
rect 18633 26869 18645 26903
rect 18517 26859 18645 26869
rect 18517 26819 18645 26829
rect 18517 26785 18547 26819
rect 18581 26785 18645 26819
rect 18517 26775 18645 26785
rect 18517 26735 18645 26745
rect 18517 26701 18531 26735
rect 18565 26701 18599 26735
rect 18633 26701 18645 26735
rect 18517 26693 18645 26701
rect 18519 26165 18719 26173
rect 18519 26131 18531 26165
rect 18565 26131 18602 26165
rect 18636 26131 18673 26165
rect 18707 26131 18719 26165
rect 18519 26121 18719 26131
rect 18519 26081 18719 26091
rect 18519 26047 18531 26081
rect 18565 26047 18599 26081
rect 18633 26047 18667 26081
rect 18701 26047 18719 26081
rect 18519 26039 18719 26047
rect 18519 26024 18647 26039
rect 18519 25984 18647 25994
rect 18519 25950 18531 25984
rect 18565 25950 18599 25984
rect 18633 25950 18647 25984
rect 18519 25942 18647 25950
rect 18519 25880 18719 25888
rect 18519 25846 18537 25880
rect 18571 25846 18605 25880
rect 18639 25846 18673 25880
rect 18707 25846 18719 25880
rect 18519 25836 18719 25846
rect 18519 25796 18719 25806
rect 18519 25762 18561 25796
rect 18595 25762 18641 25796
rect 18675 25762 18719 25796
rect 18519 25752 18719 25762
rect 18519 25710 18719 25722
rect 18519 25676 18531 25710
rect 18565 25676 18602 25710
rect 18636 25676 18673 25710
rect 18707 25676 18719 25710
rect 18519 25668 18719 25676
rect 18519 25586 18603 25594
rect 18519 25552 18539 25586
rect 18573 25552 18603 25586
rect 18519 25541 18603 25552
rect 18519 25427 18603 25511
rect 18519 25387 18603 25397
rect 18519 25353 18549 25387
rect 18583 25353 18603 25387
rect 18519 25343 18603 25353
rect 18519 25298 18603 25313
rect 18519 25292 18669 25298
rect 18519 25258 18539 25292
rect 18573 25258 18669 25292
rect 18519 25248 18669 25258
rect 18519 25208 18669 25218
rect 18519 25174 18531 25208
rect 18565 25174 18599 25208
rect 18633 25174 18669 25208
rect 18519 25131 18669 25174
rect 18519 25116 18603 25131
rect 18519 25013 18603 25086
rect 18519 24969 18603 24983
rect 18519 24935 18544 24969
rect 18578 24935 18603 24969
rect 18519 24918 18603 24935
rect 18519 24877 18603 24888
rect 18519 24843 18539 24877
rect 18573 24843 18603 24877
rect 18519 24833 18603 24843
rect 18519 24793 18603 24803
rect 18519 24759 18531 24793
rect 18565 24759 18603 24793
rect 18519 24751 18603 24759
rect 18525 24689 18653 24697
rect 18525 24655 18539 24689
rect 18573 24655 18607 24689
rect 18641 24655 18653 24689
rect 18525 24645 18653 24655
rect 18525 24605 18653 24615
rect 18525 24571 18555 24605
rect 18589 24571 18653 24605
rect 18525 24561 18653 24571
rect 18525 24521 18653 24531
rect 18525 24487 18539 24521
rect 18573 24487 18607 24521
rect 18641 24487 18653 24521
rect 18525 24479 18653 24487
rect 7573 23321 7625 23335
rect 7573 23287 7581 23321
rect 7615 23287 7625 23321
rect 7573 23253 7625 23287
rect 7573 23219 7581 23253
rect 7615 23219 7625 23253
rect 7573 23207 7625 23219
rect 7655 23305 7709 23335
rect 7655 23271 7665 23305
rect 7699 23271 7709 23305
rect 7655 23207 7709 23271
rect 7739 23321 7791 23335
rect 7739 23287 7749 23321
rect 7783 23287 7791 23321
rect 7739 23253 7791 23287
rect 7845 23329 7897 23341
rect 7845 23295 7853 23329
rect 7887 23295 7897 23329
rect 7845 23257 7897 23295
rect 7927 23321 7982 23341
rect 7927 23287 7937 23321
rect 7971 23287 7982 23321
rect 7927 23257 7982 23287
rect 8012 23316 8077 23341
rect 8012 23282 8029 23316
rect 8063 23282 8077 23316
rect 8012 23257 8077 23282
rect 8107 23257 8180 23341
rect 8210 23329 8312 23341
rect 8210 23295 8268 23329
rect 8302 23295 8312 23329
rect 8210 23261 8312 23295
rect 8210 23257 8268 23261
rect 7739 23219 7749 23253
rect 7783 23219 7791 23253
rect 7739 23207 7791 23219
rect 8225 23227 8268 23257
rect 8302 23227 8312 23261
rect 8225 23191 8312 23227
rect 8342 23321 8407 23341
rect 8342 23287 8352 23321
rect 8386 23287 8407 23321
rect 8342 23257 8407 23287
rect 8437 23311 8491 23341
rect 8437 23277 8447 23311
rect 8481 23277 8491 23311
rect 8437 23257 8491 23277
rect 8521 23257 8605 23341
rect 8635 23321 8688 23341
rect 8635 23287 8646 23321
rect 8680 23287 8688 23321
rect 8635 23257 8688 23287
rect 8762 23329 8816 23341
rect 8762 23295 8770 23329
rect 8804 23295 8816 23329
rect 8762 23258 8816 23295
rect 8342 23191 8392 23257
rect 8762 23224 8770 23258
rect 8804 23224 8816 23258
rect 8762 23187 8816 23224
rect 8762 23153 8770 23187
rect 8804 23153 8816 23187
rect 8762 23141 8816 23153
rect 8846 23299 8900 23341
rect 8846 23265 8856 23299
rect 8890 23265 8900 23299
rect 8846 23219 8900 23265
rect 8846 23185 8856 23219
rect 8890 23185 8900 23219
rect 8846 23141 8900 23185
rect 8930 23323 8982 23341
rect 8930 23289 8940 23323
rect 8974 23289 8982 23323
rect 8930 23255 8982 23289
rect 8930 23221 8940 23255
rect 8974 23221 8982 23255
rect 8930 23187 8982 23221
rect 9036 23329 9088 23341
rect 9036 23295 9044 23329
rect 9078 23295 9088 23329
rect 9036 23261 9088 23295
rect 9036 23227 9044 23261
rect 9078 23227 9088 23261
rect 9036 23213 9088 23227
rect 9118 23329 9185 23341
rect 9118 23295 9141 23329
rect 9175 23295 9185 23329
rect 9118 23261 9185 23295
rect 9118 23227 9141 23261
rect 9175 23227 9185 23261
rect 9118 23213 9185 23227
rect 8930 23153 8940 23187
rect 8974 23153 8982 23187
rect 8930 23141 8982 23153
rect 9133 23193 9185 23213
rect 9133 23159 9141 23193
rect 9175 23159 9185 23193
rect 9133 23141 9185 23159
rect 9215 23329 9267 23341
rect 9215 23295 9225 23329
rect 9259 23295 9267 23329
rect 9787 23329 9839 23343
rect 9215 23258 9267 23295
rect 9215 23224 9225 23258
rect 9259 23224 9267 23258
rect 9215 23187 9267 23224
rect 9215 23153 9225 23187
rect 9259 23153 9267 23187
rect 9215 23141 9267 23153
rect 9787 23295 9795 23329
rect 9829 23295 9839 23329
rect 9787 23261 9839 23295
rect 9787 23227 9795 23261
rect 9829 23227 9839 23261
rect 9787 23215 9839 23227
rect 9869 23313 9923 23343
rect 9869 23279 9879 23313
rect 9913 23279 9923 23313
rect 9869 23215 9923 23279
rect 9953 23329 10005 23343
rect 9953 23295 9963 23329
rect 9997 23295 10005 23329
rect 9953 23261 10005 23295
rect 10059 23337 10111 23349
rect 10059 23303 10067 23337
rect 10101 23303 10111 23337
rect 10059 23265 10111 23303
rect 10141 23329 10196 23349
rect 10141 23295 10151 23329
rect 10185 23295 10196 23329
rect 10141 23265 10196 23295
rect 10226 23324 10291 23349
rect 10226 23290 10243 23324
rect 10277 23290 10291 23324
rect 10226 23265 10291 23290
rect 10321 23265 10394 23349
rect 10424 23337 10526 23349
rect 10424 23303 10482 23337
rect 10516 23303 10526 23337
rect 10424 23269 10526 23303
rect 10424 23265 10482 23269
rect 9953 23227 9963 23261
rect 9997 23227 10005 23261
rect 9953 23215 10005 23227
rect 10439 23235 10482 23265
rect 10516 23235 10526 23269
rect 10439 23199 10526 23235
rect 10556 23329 10621 23349
rect 10556 23295 10566 23329
rect 10600 23295 10621 23329
rect 10556 23265 10621 23295
rect 10651 23319 10705 23349
rect 10651 23285 10661 23319
rect 10695 23285 10705 23319
rect 10651 23265 10705 23285
rect 10735 23265 10819 23349
rect 10849 23329 10902 23349
rect 10849 23295 10860 23329
rect 10894 23295 10902 23329
rect 10849 23265 10902 23295
rect 10976 23337 11030 23349
rect 10976 23303 10984 23337
rect 11018 23303 11030 23337
rect 10976 23266 11030 23303
rect 10556 23199 10606 23265
rect 10976 23232 10984 23266
rect 11018 23232 11030 23266
rect 10976 23195 11030 23232
rect 10976 23161 10984 23195
rect 11018 23161 11030 23195
rect 10976 23149 11030 23161
rect 11060 23307 11114 23349
rect 11060 23273 11070 23307
rect 11104 23273 11114 23307
rect 11060 23227 11114 23273
rect 11060 23193 11070 23227
rect 11104 23193 11114 23227
rect 11060 23149 11114 23193
rect 11144 23331 11196 23349
rect 11144 23297 11154 23331
rect 11188 23297 11196 23331
rect 11144 23263 11196 23297
rect 11144 23229 11154 23263
rect 11188 23229 11196 23263
rect 11144 23195 11196 23229
rect 11250 23337 11302 23349
rect 11250 23303 11258 23337
rect 11292 23303 11302 23337
rect 11250 23269 11302 23303
rect 11250 23235 11258 23269
rect 11292 23235 11302 23269
rect 11250 23221 11302 23235
rect 11332 23337 11399 23349
rect 11332 23303 11355 23337
rect 11389 23303 11399 23337
rect 11332 23269 11399 23303
rect 11332 23235 11355 23269
rect 11389 23235 11399 23269
rect 11332 23221 11399 23235
rect 11144 23161 11154 23195
rect 11188 23161 11196 23195
rect 11144 23149 11196 23161
rect 11347 23201 11399 23221
rect 11347 23167 11355 23201
rect 11389 23167 11399 23201
rect 11347 23149 11399 23167
rect 11429 23337 11481 23349
rect 11429 23303 11439 23337
rect 11473 23303 11481 23337
rect 11429 23266 11481 23303
rect 11429 23232 11439 23266
rect 11473 23232 11481 23266
rect 11429 23195 11481 23232
rect 11429 23161 11439 23195
rect 11473 23161 11481 23195
rect 11429 23149 11481 23161
rect 11987 23311 12039 23325
rect 11987 23277 11995 23311
rect 12029 23277 12039 23311
rect 11987 23243 12039 23277
rect 11987 23209 11995 23243
rect 12029 23209 12039 23243
rect 11987 23197 12039 23209
rect 12069 23295 12123 23325
rect 12069 23261 12079 23295
rect 12113 23261 12123 23295
rect 12069 23197 12123 23261
rect 12153 23311 12205 23325
rect 12153 23277 12163 23311
rect 12197 23277 12205 23311
rect 12153 23243 12205 23277
rect 12259 23319 12311 23331
rect 12259 23285 12267 23319
rect 12301 23285 12311 23319
rect 12259 23247 12311 23285
rect 12341 23311 12396 23331
rect 12341 23277 12351 23311
rect 12385 23277 12396 23311
rect 12341 23247 12396 23277
rect 12426 23306 12491 23331
rect 12426 23272 12443 23306
rect 12477 23272 12491 23306
rect 12426 23247 12491 23272
rect 12521 23247 12594 23331
rect 12624 23319 12726 23331
rect 12624 23285 12682 23319
rect 12716 23285 12726 23319
rect 12624 23251 12726 23285
rect 12624 23247 12682 23251
rect 12153 23209 12163 23243
rect 12197 23209 12205 23243
rect 12153 23197 12205 23209
rect 12639 23217 12682 23247
rect 12716 23217 12726 23251
rect 12639 23181 12726 23217
rect 12756 23311 12821 23331
rect 12756 23277 12766 23311
rect 12800 23277 12821 23311
rect 12756 23247 12821 23277
rect 12851 23301 12905 23331
rect 12851 23267 12861 23301
rect 12895 23267 12905 23301
rect 12851 23247 12905 23267
rect 12935 23247 13019 23331
rect 13049 23311 13102 23331
rect 13049 23277 13060 23311
rect 13094 23277 13102 23311
rect 13049 23247 13102 23277
rect 13176 23319 13230 23331
rect 13176 23285 13184 23319
rect 13218 23285 13230 23319
rect 13176 23248 13230 23285
rect 12756 23181 12806 23247
rect 13176 23214 13184 23248
rect 13218 23214 13230 23248
rect 13176 23177 13230 23214
rect 13176 23143 13184 23177
rect 13218 23143 13230 23177
rect 13176 23131 13230 23143
rect 13260 23289 13314 23331
rect 13260 23255 13270 23289
rect 13304 23255 13314 23289
rect 13260 23209 13314 23255
rect 13260 23175 13270 23209
rect 13304 23175 13314 23209
rect 13260 23131 13314 23175
rect 13344 23313 13396 23331
rect 13344 23279 13354 23313
rect 13388 23279 13396 23313
rect 13344 23245 13396 23279
rect 13344 23211 13354 23245
rect 13388 23211 13396 23245
rect 13344 23177 13396 23211
rect 13450 23319 13502 23331
rect 13450 23285 13458 23319
rect 13492 23285 13502 23319
rect 13450 23251 13502 23285
rect 13450 23217 13458 23251
rect 13492 23217 13502 23251
rect 13450 23203 13502 23217
rect 13532 23319 13599 23331
rect 13532 23285 13555 23319
rect 13589 23285 13599 23319
rect 13532 23251 13599 23285
rect 13532 23217 13555 23251
rect 13589 23217 13599 23251
rect 13532 23203 13599 23217
rect 13344 23143 13354 23177
rect 13388 23143 13396 23177
rect 13344 23131 13396 23143
rect 13547 23183 13599 23203
rect 13547 23149 13555 23183
rect 13589 23149 13599 23183
rect 13547 23131 13599 23149
rect 13629 23319 13681 23331
rect 13629 23285 13639 23319
rect 13673 23285 13681 23319
rect 14201 23319 14253 23333
rect 13629 23248 13681 23285
rect 13629 23214 13639 23248
rect 13673 23214 13681 23248
rect 13629 23177 13681 23214
rect 13629 23143 13639 23177
rect 13673 23143 13681 23177
rect 13629 23131 13681 23143
rect 14201 23285 14209 23319
rect 14243 23285 14253 23319
rect 14201 23251 14253 23285
rect 14201 23217 14209 23251
rect 14243 23217 14253 23251
rect 14201 23205 14253 23217
rect 14283 23303 14337 23333
rect 14283 23269 14293 23303
rect 14327 23269 14337 23303
rect 14283 23205 14337 23269
rect 14367 23319 14419 23333
rect 14367 23285 14377 23319
rect 14411 23285 14419 23319
rect 14367 23251 14419 23285
rect 14473 23327 14525 23339
rect 14473 23293 14481 23327
rect 14515 23293 14525 23327
rect 14473 23255 14525 23293
rect 14555 23319 14610 23339
rect 14555 23285 14565 23319
rect 14599 23285 14610 23319
rect 14555 23255 14610 23285
rect 14640 23314 14705 23339
rect 14640 23280 14657 23314
rect 14691 23280 14705 23314
rect 14640 23255 14705 23280
rect 14735 23255 14808 23339
rect 14838 23327 14940 23339
rect 14838 23293 14896 23327
rect 14930 23293 14940 23327
rect 14838 23259 14940 23293
rect 14838 23255 14896 23259
rect 14367 23217 14377 23251
rect 14411 23217 14419 23251
rect 14367 23205 14419 23217
rect 14853 23225 14896 23255
rect 14930 23225 14940 23259
rect 14853 23189 14940 23225
rect 14970 23319 15035 23339
rect 14970 23285 14980 23319
rect 15014 23285 15035 23319
rect 14970 23255 15035 23285
rect 15065 23309 15119 23339
rect 15065 23275 15075 23309
rect 15109 23275 15119 23309
rect 15065 23255 15119 23275
rect 15149 23255 15233 23339
rect 15263 23319 15316 23339
rect 15263 23285 15274 23319
rect 15308 23285 15316 23319
rect 15263 23255 15316 23285
rect 15390 23327 15444 23339
rect 15390 23293 15398 23327
rect 15432 23293 15444 23327
rect 15390 23256 15444 23293
rect 14970 23189 15020 23255
rect 15390 23222 15398 23256
rect 15432 23222 15444 23256
rect 15390 23185 15444 23222
rect 15390 23151 15398 23185
rect 15432 23151 15444 23185
rect 15390 23139 15444 23151
rect 15474 23297 15528 23339
rect 15474 23263 15484 23297
rect 15518 23263 15528 23297
rect 15474 23217 15528 23263
rect 15474 23183 15484 23217
rect 15518 23183 15528 23217
rect 15474 23139 15528 23183
rect 15558 23321 15610 23339
rect 15558 23287 15568 23321
rect 15602 23287 15610 23321
rect 15558 23253 15610 23287
rect 15558 23219 15568 23253
rect 15602 23219 15610 23253
rect 15558 23185 15610 23219
rect 15664 23327 15716 23339
rect 15664 23293 15672 23327
rect 15706 23293 15716 23327
rect 15664 23259 15716 23293
rect 15664 23225 15672 23259
rect 15706 23225 15716 23259
rect 15664 23211 15716 23225
rect 15746 23327 15813 23339
rect 15746 23293 15769 23327
rect 15803 23293 15813 23327
rect 15746 23259 15813 23293
rect 15746 23225 15769 23259
rect 15803 23225 15813 23259
rect 15746 23211 15813 23225
rect 15558 23151 15568 23185
rect 15602 23151 15610 23185
rect 15558 23139 15610 23151
rect 15761 23191 15813 23211
rect 15761 23157 15769 23191
rect 15803 23157 15813 23191
rect 15761 23139 15813 23157
rect 15843 23327 15895 23339
rect 15843 23293 15853 23327
rect 15887 23293 15895 23327
rect 16507 23327 16559 23341
rect 15843 23256 15895 23293
rect 15843 23222 15853 23256
rect 15887 23222 15895 23256
rect 15843 23185 15895 23222
rect 15843 23151 15853 23185
rect 15887 23151 15895 23185
rect 15843 23139 15895 23151
rect 16507 23293 16515 23327
rect 16549 23293 16559 23327
rect 16507 23259 16559 23293
rect 16507 23225 16515 23259
rect 16549 23225 16559 23259
rect 16507 23213 16559 23225
rect 16589 23311 16643 23341
rect 16589 23277 16599 23311
rect 16633 23277 16643 23311
rect 16589 23213 16643 23277
rect 16673 23327 16725 23341
rect 16673 23293 16683 23327
rect 16717 23293 16725 23327
rect 16673 23259 16725 23293
rect 16779 23335 16831 23347
rect 16779 23301 16787 23335
rect 16821 23301 16831 23335
rect 16779 23263 16831 23301
rect 16861 23327 16916 23347
rect 16861 23293 16871 23327
rect 16905 23293 16916 23327
rect 16861 23263 16916 23293
rect 16946 23322 17011 23347
rect 16946 23288 16963 23322
rect 16997 23288 17011 23322
rect 16946 23263 17011 23288
rect 17041 23263 17114 23347
rect 17144 23335 17246 23347
rect 17144 23301 17202 23335
rect 17236 23301 17246 23335
rect 17144 23267 17246 23301
rect 17144 23263 17202 23267
rect 16673 23225 16683 23259
rect 16717 23225 16725 23259
rect 16673 23213 16725 23225
rect 17159 23233 17202 23263
rect 17236 23233 17246 23267
rect 17159 23197 17246 23233
rect 17276 23327 17341 23347
rect 17276 23293 17286 23327
rect 17320 23293 17341 23327
rect 17276 23263 17341 23293
rect 17371 23317 17425 23347
rect 17371 23283 17381 23317
rect 17415 23283 17425 23317
rect 17371 23263 17425 23283
rect 17455 23263 17539 23347
rect 17569 23327 17622 23347
rect 17569 23293 17580 23327
rect 17614 23293 17622 23327
rect 17569 23263 17622 23293
rect 17696 23335 17750 23347
rect 17696 23301 17704 23335
rect 17738 23301 17750 23335
rect 17696 23264 17750 23301
rect 17276 23197 17326 23263
rect 17696 23230 17704 23264
rect 17738 23230 17750 23264
rect 17696 23193 17750 23230
rect 17696 23159 17704 23193
rect 17738 23159 17750 23193
rect 17696 23147 17750 23159
rect 17780 23305 17834 23347
rect 17780 23271 17790 23305
rect 17824 23271 17834 23305
rect 17780 23225 17834 23271
rect 17780 23191 17790 23225
rect 17824 23191 17834 23225
rect 17780 23147 17834 23191
rect 17864 23329 17916 23347
rect 17864 23295 17874 23329
rect 17908 23295 17916 23329
rect 17864 23261 17916 23295
rect 17864 23227 17874 23261
rect 17908 23227 17916 23261
rect 17864 23193 17916 23227
rect 17970 23335 18022 23347
rect 17970 23301 17978 23335
rect 18012 23301 18022 23335
rect 17970 23267 18022 23301
rect 17970 23233 17978 23267
rect 18012 23233 18022 23267
rect 17970 23219 18022 23233
rect 18052 23335 18119 23347
rect 18052 23301 18075 23335
rect 18109 23301 18119 23335
rect 18052 23267 18119 23301
rect 18052 23233 18075 23267
rect 18109 23233 18119 23267
rect 18052 23219 18119 23233
rect 17864 23159 17874 23193
rect 17908 23159 17916 23193
rect 17864 23147 17916 23159
rect 18067 23199 18119 23219
rect 18067 23165 18075 23199
rect 18109 23165 18119 23199
rect 18067 23147 18119 23165
rect 18149 23335 18201 23347
rect 18149 23301 18159 23335
rect 18193 23301 18201 23335
rect 18149 23264 18201 23301
rect 18149 23230 18159 23264
rect 18193 23230 18201 23264
rect 18149 23193 18201 23230
rect 18149 23159 18159 23193
rect 18193 23159 18201 23193
rect 18149 23147 18201 23159
rect 15641 17331 15693 17349
rect 15641 17297 15649 17331
rect 15683 17297 15693 17331
rect 15641 17263 15693 17297
rect 15641 17229 15649 17263
rect 15683 17229 15693 17263
rect 15641 17195 15693 17229
rect 15641 17161 15649 17195
rect 15683 17161 15693 17195
rect 15641 17149 15693 17161
rect 15723 17331 15775 17349
rect 15723 17297 15733 17331
rect 15767 17297 15775 17331
rect 15723 17263 15775 17297
rect 15723 17229 15733 17263
rect 15767 17229 15775 17263
rect 15723 17195 15775 17229
rect 16419 17369 16471 17387
rect 16419 17335 16427 17369
rect 16461 17335 16471 17369
rect 16419 17301 16471 17335
rect 16419 17267 16427 17301
rect 16461 17267 16471 17301
rect 16419 17233 16471 17267
rect 15723 17161 15733 17195
rect 15767 17161 15775 17195
rect 16419 17199 16427 17233
rect 16461 17199 16471 17233
rect 16419 17187 16471 17199
rect 16501 17369 16553 17387
rect 16501 17335 16511 17369
rect 16545 17335 16553 17369
rect 16501 17301 16553 17335
rect 16501 17267 16511 17301
rect 16545 17267 16553 17301
rect 16501 17233 16553 17267
rect 16501 17199 16511 17233
rect 16545 17199 16553 17233
rect 17293 17371 17345 17389
rect 17293 17337 17301 17371
rect 17335 17337 17345 17371
rect 17293 17303 17345 17337
rect 17293 17269 17301 17303
rect 17335 17269 17345 17303
rect 17293 17235 17345 17269
rect 16501 17187 16553 17199
rect 17293 17201 17301 17235
rect 17335 17201 17345 17235
rect 17293 17189 17345 17201
rect 17375 17371 17427 17389
rect 17375 17337 17385 17371
rect 17419 17337 17427 17371
rect 17375 17303 17427 17337
rect 17375 17269 17385 17303
rect 17419 17269 17427 17303
rect 17375 17235 17427 17269
rect 17375 17201 17385 17235
rect 17419 17201 17427 17235
rect 17375 17189 17427 17201
rect 18061 17361 18113 17379
rect 18061 17327 18069 17361
rect 18103 17327 18113 17361
rect 18061 17293 18113 17327
rect 18061 17259 18069 17293
rect 18103 17259 18113 17293
rect 18061 17225 18113 17259
rect 18061 17191 18069 17225
rect 18103 17191 18113 17225
rect 18061 17179 18113 17191
rect 18143 17361 18195 17379
rect 18143 17327 18153 17361
rect 18187 17327 18195 17361
rect 18143 17293 18195 17327
rect 18143 17259 18153 17293
rect 18187 17259 18195 17293
rect 18143 17225 18195 17259
rect 18143 17191 18153 17225
rect 18187 17191 18195 17225
rect 19183 17363 19235 17381
rect 19183 17329 19191 17363
rect 19225 17329 19235 17363
rect 19183 17295 19235 17329
rect 19183 17261 19191 17295
rect 19225 17261 19235 17295
rect 19183 17227 19235 17261
rect 18143 17179 18195 17191
rect 19183 17193 19191 17227
rect 19225 17193 19235 17227
rect 19183 17181 19235 17193
rect 19265 17363 19317 17381
rect 19265 17329 19275 17363
rect 19309 17329 19317 17363
rect 19265 17295 19317 17329
rect 19265 17261 19275 17295
rect 19309 17261 19317 17295
rect 19265 17227 19317 17261
rect 19265 17193 19275 17227
rect 19309 17193 19317 17227
rect 20057 17365 20109 17383
rect 20057 17331 20065 17365
rect 20099 17331 20109 17365
rect 20057 17297 20109 17331
rect 20057 17263 20065 17297
rect 20099 17263 20109 17297
rect 20057 17229 20109 17263
rect 19265 17181 19317 17193
rect 20057 17195 20065 17229
rect 20099 17195 20109 17229
rect 20057 17183 20109 17195
rect 20139 17365 20191 17383
rect 20139 17331 20149 17365
rect 20183 17331 20191 17365
rect 20139 17297 20191 17331
rect 20139 17263 20149 17297
rect 20183 17263 20191 17297
rect 20139 17229 20191 17263
rect 20139 17195 20149 17229
rect 20183 17195 20191 17229
rect 20139 17183 20191 17195
rect 20825 17355 20877 17373
rect 20825 17321 20833 17355
rect 20867 17321 20877 17355
rect 20825 17287 20877 17321
rect 20825 17253 20833 17287
rect 20867 17253 20877 17287
rect 20825 17219 20877 17253
rect 20825 17185 20833 17219
rect 20867 17185 20877 17219
rect 15723 17149 15775 17161
rect 20825 17173 20877 17185
rect 20907 17355 20959 17373
rect 20907 17321 20917 17355
rect 20951 17321 20959 17355
rect 20907 17287 20959 17321
rect 20907 17253 20917 17287
rect 20951 17253 20959 17287
rect 20907 17219 20959 17253
rect 20907 17185 20917 17219
rect 20951 17185 20959 17219
rect 20907 17173 20959 17185
rect 21439 17353 21491 17371
rect 21439 17319 21447 17353
rect 21481 17319 21491 17353
rect 21439 17285 21491 17319
rect 21439 17251 21447 17285
rect 21481 17251 21491 17285
rect 21439 17217 21491 17251
rect 21439 17183 21447 17217
rect 21481 17183 21491 17217
rect 21439 17171 21491 17183
rect 21521 17353 21573 17371
rect 21521 17319 21531 17353
rect 21565 17319 21573 17353
rect 21521 17285 21573 17319
rect 21521 17251 21531 17285
rect 21565 17251 21573 17285
rect 21521 17217 21573 17251
rect 21521 17183 21531 17217
rect 21565 17183 21573 17217
rect 22313 17355 22365 17373
rect 22313 17321 22321 17355
rect 22355 17321 22365 17355
rect 22313 17287 22365 17321
rect 22313 17253 22321 17287
rect 22355 17253 22365 17287
rect 22313 17219 22365 17253
rect 21521 17171 21573 17183
rect 22313 17185 22321 17219
rect 22355 17185 22365 17219
rect 22313 17173 22365 17185
rect 22395 17355 22447 17373
rect 22395 17321 22405 17355
rect 22439 17321 22447 17355
rect 22395 17287 22447 17321
rect 22395 17253 22405 17287
rect 22439 17253 22447 17287
rect 22395 17219 22447 17253
rect 22395 17185 22405 17219
rect 22439 17185 22447 17219
rect 22395 17173 22447 17185
rect 23081 17345 23133 17363
rect 23081 17311 23089 17345
rect 23123 17311 23133 17345
rect 23081 17277 23133 17311
rect 23081 17243 23089 17277
rect 23123 17243 23133 17277
rect 23081 17209 23133 17243
rect 23081 17175 23089 17209
rect 23123 17175 23133 17209
rect 23081 17163 23133 17175
rect 23163 17345 23215 17363
rect 23163 17311 23173 17345
rect 23207 17311 23215 17345
rect 23163 17277 23215 17311
rect 23163 17243 23173 17277
rect 23207 17243 23215 17277
rect 23163 17209 23215 17243
rect 23163 17175 23173 17209
rect 23207 17175 23215 17209
rect 23163 17163 23215 17175
rect 9369 16531 9421 16543
rect 9369 16497 9377 16531
rect 9411 16497 9421 16531
rect 9369 16463 9421 16497
rect 9369 16429 9377 16463
rect 9411 16429 9421 16463
rect 9369 16343 9421 16429
rect 9451 16343 9505 16543
rect 9535 16521 9589 16543
rect 9535 16487 9545 16521
rect 9579 16487 9589 16521
rect 9535 16453 9589 16487
rect 9535 16419 9545 16453
rect 9579 16419 9589 16453
rect 9535 16343 9589 16419
rect 9619 16521 9673 16543
rect 9619 16487 9629 16521
rect 9663 16487 9673 16521
rect 9619 16453 9673 16487
rect 9619 16419 9629 16453
rect 9663 16419 9673 16453
rect 9619 16343 9673 16419
rect 9703 16521 9755 16543
rect 9703 16487 9713 16521
rect 9747 16487 9755 16521
rect 9703 16343 9755 16487
rect 9809 16521 9861 16543
rect 9809 16487 9817 16521
rect 9851 16487 9861 16521
rect 9809 16453 9861 16487
rect 9809 16419 9817 16453
rect 9851 16419 9861 16453
rect 9809 16343 9861 16419
rect 9891 16523 9951 16543
rect 9891 16489 9901 16523
rect 9935 16489 9951 16523
rect 9891 16455 9951 16489
rect 9891 16421 9901 16455
rect 9935 16421 9951 16455
rect 9891 16387 9951 16421
rect 9891 16353 9901 16387
rect 9935 16353 9951 16387
rect 9891 16343 9951 16353
rect 9687 15787 9739 15799
rect 9687 15757 9695 15787
rect 9491 15745 9547 15757
rect 9491 15711 9503 15745
rect 9537 15711 9547 15745
rect 9491 15673 9547 15711
rect 9577 15745 9631 15757
rect 9577 15711 9587 15745
rect 9621 15711 9631 15745
rect 9577 15673 9631 15711
rect 9661 15753 9695 15757
rect 9729 15753 9739 15787
rect 9661 15719 9739 15753
rect 9661 15685 9695 15719
rect 9729 15685 9739 15719
rect 9661 15673 9739 15685
rect 9677 15599 9739 15673
rect 9769 15787 9864 15799
rect 9769 15753 9799 15787
rect 9833 15753 9864 15787
rect 9769 15719 9864 15753
rect 9769 15685 9799 15719
rect 9833 15685 9864 15719
rect 9769 15599 9864 15685
rect 11501 15677 11553 15689
rect 11501 15643 11509 15677
rect 11543 15643 11553 15677
rect 11501 15605 11553 15643
rect 11583 15669 11653 15689
rect 11583 15635 11601 15669
rect 11635 15635 11653 15669
rect 11583 15605 11653 15635
rect 11683 15677 11757 15689
rect 11683 15643 11703 15677
rect 11737 15643 11757 15677
rect 11683 15605 11757 15643
rect 11787 15669 11843 15689
rect 11787 15635 11798 15669
rect 11832 15635 11843 15669
rect 11787 15605 11843 15635
rect 11873 15677 12009 15689
rect 11873 15643 11949 15677
rect 11983 15643 12009 15677
rect 11873 15609 12009 15643
rect 11873 15605 11949 15609
rect 11892 15575 11949 15605
rect 11983 15575 12009 15609
rect 11892 15489 12009 15575
rect 12039 15677 12091 15689
rect 12039 15643 12049 15677
rect 12083 15643 12091 15677
rect 12039 15609 12091 15643
rect 12039 15575 12049 15609
rect 12083 15575 12091 15609
rect 12039 15541 12091 15575
rect 12039 15507 12049 15541
rect 12083 15507 12091 15541
rect 12039 15489 12091 15507
rect 10871 15177 10923 15189
rect 10871 15147 10879 15177
rect 10675 15135 10731 15147
rect 10675 15101 10687 15135
rect 10721 15101 10731 15135
rect 10675 15063 10731 15101
rect 10761 15135 10815 15147
rect 10761 15101 10771 15135
rect 10805 15101 10815 15135
rect 10761 15063 10815 15101
rect 10845 15143 10879 15147
rect 10913 15143 10923 15177
rect 10845 15109 10923 15143
rect 10845 15075 10879 15109
rect 10913 15075 10923 15109
rect 10845 15063 10923 15075
rect 9379 14967 9431 14979
rect 9379 14933 9387 14967
rect 9421 14933 9431 14967
rect 9379 14899 9431 14933
rect 9379 14865 9387 14899
rect 9421 14865 9431 14899
rect 9379 14779 9431 14865
rect 9461 14779 9515 14979
rect 9545 14957 9599 14979
rect 9545 14923 9555 14957
rect 9589 14923 9599 14957
rect 9545 14889 9599 14923
rect 9545 14855 9555 14889
rect 9589 14855 9599 14889
rect 9545 14779 9599 14855
rect 9629 14957 9683 14979
rect 9629 14923 9639 14957
rect 9673 14923 9683 14957
rect 9629 14889 9683 14923
rect 9629 14855 9639 14889
rect 9673 14855 9683 14889
rect 9629 14779 9683 14855
rect 9713 14957 9765 14979
rect 9713 14923 9723 14957
rect 9757 14923 9765 14957
rect 9713 14779 9765 14923
rect 9819 14957 9871 14979
rect 9819 14923 9827 14957
rect 9861 14923 9871 14957
rect 9819 14889 9871 14923
rect 9819 14855 9827 14889
rect 9861 14855 9871 14889
rect 9819 14779 9871 14855
rect 9901 14959 9961 14979
rect 9901 14925 9911 14959
rect 9945 14925 9961 14959
rect 9901 14891 9961 14925
rect 9901 14857 9911 14891
rect 9945 14857 9961 14891
rect 9901 14823 9961 14857
rect 10861 14989 10923 15063
rect 10953 15177 11048 15189
rect 10953 15143 10983 15177
rect 11017 15143 11048 15177
rect 10953 15109 11048 15143
rect 10953 15075 10983 15109
rect 11017 15075 11048 15109
rect 10953 14989 11048 15075
rect 9901 14789 9911 14823
rect 9945 14789 9961 14823
rect 9901 14779 9961 14789
rect 9697 14223 9749 14235
rect 9697 14193 9705 14223
rect 9501 14181 9557 14193
rect 9501 14147 9513 14181
rect 9547 14147 9557 14181
rect 9501 14109 9557 14147
rect 9587 14181 9641 14193
rect 9587 14147 9597 14181
rect 9631 14147 9641 14181
rect 9587 14109 9641 14147
rect 9671 14189 9705 14193
rect 9739 14189 9749 14223
rect 9671 14155 9749 14189
rect 9671 14121 9705 14155
rect 9739 14121 9749 14155
rect 9671 14109 9749 14121
rect 9687 14035 9749 14109
rect 9779 14223 9874 14235
rect 9779 14189 9809 14223
rect 9843 14189 9874 14223
rect 9779 14155 9874 14189
rect 9779 14121 9809 14155
rect 9843 14121 9874 14155
rect 10717 14211 10769 14223
rect 10717 14177 10725 14211
rect 10759 14177 10769 14211
rect 10717 14139 10769 14177
rect 10799 14203 10869 14223
rect 10799 14169 10817 14203
rect 10851 14169 10869 14203
rect 10799 14139 10869 14169
rect 10899 14211 10973 14223
rect 10899 14177 10919 14211
rect 10953 14177 10973 14211
rect 10899 14139 10973 14177
rect 11003 14203 11059 14223
rect 11003 14169 11014 14203
rect 11048 14169 11059 14203
rect 11003 14139 11059 14169
rect 11089 14211 11225 14223
rect 11089 14177 11165 14211
rect 11199 14177 11225 14211
rect 11089 14143 11225 14177
rect 11089 14139 11165 14143
rect 9779 14035 9874 14121
rect 11108 14109 11165 14139
rect 11199 14109 11225 14143
rect 11108 14023 11225 14109
rect 11255 14211 11307 14223
rect 11255 14177 11265 14211
rect 11299 14177 11307 14211
rect 12976 14195 13029 14207
rect 11255 14143 11307 14177
rect 11255 14109 11265 14143
rect 11299 14109 11307 14143
rect 12976 14161 12984 14195
rect 13018 14161 13029 14195
rect 11255 14075 11307 14109
rect 12976 14127 13029 14161
rect 12976 14093 12984 14127
rect 13018 14093 13029 14127
rect 12976 14091 13029 14093
rect 11255 14041 11265 14075
rect 11299 14041 11307 14075
rect 11255 14023 11307 14041
rect 12615 14064 12667 14091
rect 12615 14030 12623 14064
rect 12657 14030 12667 14064
rect 12615 14007 12667 14030
rect 12697 14007 12763 14091
rect 12793 14007 12835 14091
rect 12865 14007 12931 14091
rect 12961 14007 13029 14091
rect 13059 14164 13113 14207
rect 13059 14130 13069 14164
rect 13103 14130 13113 14164
rect 13059 14096 13113 14130
rect 13059 14062 13069 14096
rect 13103 14062 13113 14096
rect 13059 14007 13113 14062
rect 11897 13821 11949 13849
rect 11897 13787 11905 13821
rect 11939 13787 11949 13821
rect 11897 13753 11949 13787
rect 11897 13733 11905 13753
rect 11728 13701 11780 13733
rect 11728 13667 11736 13701
rect 11770 13667 11780 13701
rect 11728 13649 11780 13667
rect 11810 13649 11852 13733
rect 11882 13719 11905 13733
rect 11939 13719 11949 13753
rect 11882 13649 11949 13719
rect 11979 13837 12047 13849
rect 11979 13803 12005 13837
rect 12039 13803 12047 13837
rect 11979 13769 12047 13803
rect 11979 13735 12005 13769
rect 12039 13735 12047 13769
rect 11979 13649 12047 13735
rect 9371 13299 9423 13311
rect 9371 13265 9379 13299
rect 9413 13265 9423 13299
rect 9371 13231 9423 13265
rect 9371 13197 9379 13231
rect 9413 13197 9423 13231
rect 9371 13111 9423 13197
rect 9453 13111 9507 13311
rect 9537 13289 9591 13311
rect 9537 13255 9547 13289
rect 9581 13255 9591 13289
rect 9537 13221 9591 13255
rect 9537 13187 9547 13221
rect 9581 13187 9591 13221
rect 9537 13111 9591 13187
rect 9621 13289 9675 13311
rect 9621 13255 9631 13289
rect 9665 13255 9675 13289
rect 9621 13221 9675 13255
rect 9621 13187 9631 13221
rect 9665 13187 9675 13221
rect 9621 13111 9675 13187
rect 9705 13289 9757 13311
rect 9705 13255 9715 13289
rect 9749 13255 9757 13289
rect 9705 13111 9757 13255
rect 9811 13289 9863 13311
rect 9811 13255 9819 13289
rect 9853 13255 9863 13289
rect 9811 13221 9863 13255
rect 9811 13187 9819 13221
rect 9853 13187 9863 13221
rect 9811 13111 9863 13187
rect 9893 13291 9953 13311
rect 11113 13369 11165 13381
rect 11113 13335 11121 13369
rect 11155 13335 11165 13369
rect 11113 13322 11165 13335
rect 9893 13257 9903 13291
rect 9937 13257 9953 13291
rect 11115 13268 11165 13322
rect 9893 13223 9953 13257
rect 9893 13189 9903 13223
rect 9937 13189 9953 13223
rect 9893 13155 9953 13189
rect 10841 13230 10893 13268
rect 10841 13196 10849 13230
rect 10883 13196 10893 13230
rect 10841 13184 10893 13196
rect 10923 13260 10977 13268
rect 10923 13226 10933 13260
rect 10967 13226 10977 13260
rect 10923 13184 10977 13226
rect 11007 13241 11070 13268
rect 11007 13207 11026 13241
rect 11060 13207 11070 13241
rect 11007 13184 11070 13207
rect 11100 13184 11165 13268
rect 9893 13121 9903 13155
rect 9937 13121 9953 13155
rect 9893 13111 9953 13121
rect 11115 13181 11165 13184
rect 11195 13355 11247 13381
rect 11195 13321 11205 13355
rect 11239 13321 11247 13355
rect 11195 13287 11247 13321
rect 11195 13253 11205 13287
rect 11239 13253 11247 13287
rect 11195 13181 11247 13253
rect 9689 12555 9741 12567
rect 9689 12525 9697 12555
rect 9493 12513 9549 12525
rect 9493 12479 9505 12513
rect 9539 12479 9549 12513
rect 9493 12441 9549 12479
rect 9579 12513 9633 12525
rect 9579 12479 9589 12513
rect 9623 12479 9633 12513
rect 9579 12441 9633 12479
rect 9663 12521 9697 12525
rect 9731 12521 9741 12555
rect 9663 12487 9741 12521
rect 9663 12453 9697 12487
rect 9731 12453 9741 12487
rect 9663 12441 9741 12453
rect 9679 12367 9741 12441
rect 9771 12555 9866 12567
rect 9771 12521 9801 12555
rect 9835 12521 9866 12555
rect 9771 12487 9866 12521
rect 9771 12453 9801 12487
rect 9835 12453 9866 12487
rect 9771 12367 9866 12453
rect 11065 12349 11117 12361
rect 11065 12319 11073 12349
rect 10869 12307 10925 12319
rect 10869 12273 10881 12307
rect 10915 12273 10925 12307
rect 10869 12235 10925 12273
rect 10955 12307 11009 12319
rect 10955 12273 10965 12307
rect 10999 12273 11009 12307
rect 10955 12235 11009 12273
rect 11039 12315 11073 12319
rect 11107 12315 11117 12349
rect 11039 12281 11117 12315
rect 11039 12247 11073 12281
rect 11107 12247 11117 12281
rect 11039 12235 11117 12247
rect 11055 12161 11117 12235
rect 11147 12349 11242 12361
rect 11147 12315 11177 12349
rect 11211 12315 11242 12349
rect 11147 12281 11242 12315
rect 11147 12247 11177 12281
rect 11211 12247 11242 12281
rect 11147 12161 11242 12247
rect 9381 11735 9433 11747
rect 9381 11701 9389 11735
rect 9423 11701 9433 11735
rect 9381 11667 9433 11701
rect 9381 11633 9389 11667
rect 9423 11633 9433 11667
rect 9381 11547 9433 11633
rect 9463 11547 9517 11747
rect 9547 11725 9601 11747
rect 9547 11691 9557 11725
rect 9591 11691 9601 11725
rect 9547 11657 9601 11691
rect 9547 11623 9557 11657
rect 9591 11623 9601 11657
rect 9547 11547 9601 11623
rect 9631 11725 9685 11747
rect 9631 11691 9641 11725
rect 9675 11691 9685 11725
rect 9631 11657 9685 11691
rect 9631 11623 9641 11657
rect 9675 11623 9685 11657
rect 9631 11547 9685 11623
rect 9715 11725 9767 11747
rect 9715 11691 9725 11725
rect 9759 11691 9767 11725
rect 9715 11547 9767 11691
rect 9821 11725 9873 11747
rect 9821 11691 9829 11725
rect 9863 11691 9873 11725
rect 9821 11657 9873 11691
rect 9821 11623 9829 11657
rect 9863 11623 9873 11657
rect 9821 11547 9873 11623
rect 9903 11727 9963 11747
rect 9903 11693 9913 11727
rect 9947 11693 9963 11727
rect 9903 11659 9963 11693
rect 9903 11625 9913 11659
rect 9947 11625 9963 11659
rect 9903 11591 9963 11625
rect 9903 11557 9913 11591
rect 9947 11557 9963 11591
rect 9903 11547 9963 11557
rect 9699 10991 9751 11003
rect 9699 10961 9707 10991
rect 9503 10949 9559 10961
rect 9503 10915 9515 10949
rect 9549 10915 9559 10949
rect 9503 10877 9559 10915
rect 9589 10949 9643 10961
rect 9589 10915 9599 10949
rect 9633 10915 9643 10949
rect 9589 10877 9643 10915
rect 9673 10957 9707 10961
rect 9741 10957 9751 10991
rect 9673 10923 9751 10957
rect 9673 10889 9707 10923
rect 9741 10889 9751 10923
rect 9673 10877 9751 10889
rect 9689 10803 9751 10877
rect 9781 10991 9876 11003
rect 9781 10957 9811 10991
rect 9845 10957 9876 10991
rect 9781 10923 9876 10957
rect 9781 10889 9811 10923
rect 9845 10889 9876 10923
rect 9781 10803 9876 10889
rect 6186 6285 6238 6303
rect 6186 6251 6194 6285
rect 6228 6251 6238 6285
rect 6186 6217 6238 6251
rect 6186 6183 6194 6217
rect 6228 6183 6238 6217
rect 6186 6149 6238 6183
rect 6186 6115 6194 6149
rect 6228 6115 6238 6149
rect 6186 6103 6238 6115
rect 6268 6285 6320 6303
rect 6268 6251 6278 6285
rect 6312 6251 6320 6285
rect 6268 6217 6320 6251
rect 6268 6183 6278 6217
rect 6312 6183 6320 6217
rect 6268 6149 6320 6183
rect 6268 6115 6278 6149
rect 6312 6115 6320 6149
rect 6268 6103 6320 6115
rect 10080 5633 10132 5671
rect 10080 5599 10088 5633
rect 10122 5599 10132 5633
rect 10080 5543 10132 5599
rect 1898 5213 1950 5251
rect 1898 5179 1906 5213
rect 1940 5179 1950 5213
rect 1898 5123 1950 5179
rect 1898 5089 1906 5123
rect 1940 5089 1950 5123
rect 1898 5051 1950 5089
rect 1980 5135 2032 5251
rect 10080 5509 10088 5543
rect 10122 5509 10132 5543
rect 3147 5135 3199 5251
rect 1980 5093 2049 5135
rect 1980 5059 1990 5093
rect 2024 5059 2049 5093
rect 1980 5051 2049 5059
rect 2079 5051 2145 5135
rect 2175 5051 2217 5135
rect 2247 5105 2313 5135
rect 2247 5071 2257 5105
rect 2291 5071 2313 5105
rect 2247 5051 2313 5071
rect 2343 5110 2402 5135
rect 2343 5076 2358 5110
rect 2392 5076 2402 5110
rect 2343 5051 2402 5076
rect 2432 5093 2486 5135
rect 2432 5059 2442 5093
rect 2476 5059 2486 5093
rect 2432 5051 2486 5059
rect 2516 5110 2570 5135
rect 2516 5076 2526 5110
rect 2560 5076 2570 5110
rect 2516 5051 2570 5076
rect 2600 5097 2652 5135
rect 2600 5063 2610 5097
rect 2644 5063 2652 5097
rect 2600 5051 2652 5063
rect 2706 5110 2758 5135
rect 2706 5076 2714 5110
rect 2748 5076 2758 5110
rect 2706 5051 2758 5076
rect 2788 5093 2842 5135
rect 2788 5059 2798 5093
rect 2832 5059 2842 5093
rect 2788 5051 2842 5059
rect 2872 5110 2926 5135
rect 2872 5076 2882 5110
rect 2916 5076 2926 5110
rect 2872 5051 2926 5076
rect 2956 5110 3010 5135
rect 2956 5076 2966 5110
rect 3000 5076 3010 5110
rect 2956 5051 3010 5076
rect 3040 5051 3100 5135
rect 3130 5101 3199 5135
rect 3130 5067 3155 5101
rect 3189 5067 3199 5101
rect 3130 5051 3199 5067
rect 3229 5210 3281 5251
rect 3229 5176 3239 5210
rect 3273 5176 3281 5210
rect 3229 5116 3281 5176
rect 3229 5082 3239 5116
rect 3273 5082 3281 5116
rect 3229 5051 3281 5082
rect 4032 5205 4084 5243
rect 4032 5171 4040 5205
rect 4074 5171 4084 5205
rect 4032 5115 4084 5171
rect 4032 5081 4040 5115
rect 4074 5081 4084 5115
rect 4032 5043 4084 5081
rect 4114 5127 4166 5243
rect 5281 5127 5333 5243
rect 4114 5085 4183 5127
rect 4114 5051 4124 5085
rect 4158 5051 4183 5085
rect 4114 5043 4183 5051
rect 4213 5043 4279 5127
rect 4309 5043 4351 5127
rect 4381 5097 4447 5127
rect 4381 5063 4391 5097
rect 4425 5063 4447 5097
rect 4381 5043 4447 5063
rect 4477 5102 4536 5127
rect 4477 5068 4492 5102
rect 4526 5068 4536 5102
rect 4477 5043 4536 5068
rect 4566 5085 4620 5127
rect 4566 5051 4576 5085
rect 4610 5051 4620 5085
rect 4566 5043 4620 5051
rect 4650 5102 4704 5127
rect 4650 5068 4660 5102
rect 4694 5068 4704 5102
rect 4650 5043 4704 5068
rect 4734 5089 4786 5127
rect 4734 5055 4744 5089
rect 4778 5055 4786 5089
rect 4734 5043 4786 5055
rect 4840 5102 4892 5127
rect 4840 5068 4848 5102
rect 4882 5068 4892 5102
rect 4840 5043 4892 5068
rect 4922 5085 4976 5127
rect 4922 5051 4932 5085
rect 4966 5051 4976 5085
rect 4922 5043 4976 5051
rect 5006 5102 5060 5127
rect 5006 5068 5016 5102
rect 5050 5068 5060 5102
rect 5006 5043 5060 5068
rect 5090 5102 5144 5127
rect 5090 5068 5100 5102
rect 5134 5068 5144 5102
rect 5090 5043 5144 5068
rect 5174 5043 5234 5127
rect 5264 5093 5333 5127
rect 5264 5059 5289 5093
rect 5323 5059 5333 5093
rect 5264 5043 5333 5059
rect 5363 5202 5415 5243
rect 5363 5168 5373 5202
rect 5407 5168 5415 5202
rect 5363 5108 5415 5168
rect 5363 5074 5373 5108
rect 5407 5074 5415 5108
rect 5363 5043 5415 5074
rect 5984 5205 6036 5243
rect 5984 5171 5992 5205
rect 6026 5171 6036 5205
rect 5984 5115 6036 5171
rect 5984 5081 5992 5115
rect 6026 5081 6036 5115
rect 5984 5043 6036 5081
rect 6066 5127 6118 5243
rect 7233 5127 7285 5243
rect 6066 5085 6135 5127
rect 6066 5051 6076 5085
rect 6110 5051 6135 5085
rect 6066 5043 6135 5051
rect 6165 5043 6231 5127
rect 6261 5043 6303 5127
rect 6333 5097 6399 5127
rect 6333 5063 6343 5097
rect 6377 5063 6399 5097
rect 6333 5043 6399 5063
rect 6429 5102 6488 5127
rect 6429 5068 6444 5102
rect 6478 5068 6488 5102
rect 6429 5043 6488 5068
rect 6518 5085 6572 5127
rect 6518 5051 6528 5085
rect 6562 5051 6572 5085
rect 6518 5043 6572 5051
rect 6602 5102 6656 5127
rect 6602 5068 6612 5102
rect 6646 5068 6656 5102
rect 6602 5043 6656 5068
rect 6686 5089 6738 5127
rect 6686 5055 6696 5089
rect 6730 5055 6738 5089
rect 6686 5043 6738 5055
rect 6792 5102 6844 5127
rect 6792 5068 6800 5102
rect 6834 5068 6844 5102
rect 6792 5043 6844 5068
rect 6874 5085 6928 5127
rect 6874 5051 6884 5085
rect 6918 5051 6928 5085
rect 6874 5043 6928 5051
rect 6958 5102 7012 5127
rect 6958 5068 6968 5102
rect 7002 5068 7012 5102
rect 6958 5043 7012 5068
rect 7042 5102 7096 5127
rect 7042 5068 7052 5102
rect 7086 5068 7096 5102
rect 7042 5043 7096 5068
rect 7126 5043 7186 5127
rect 7216 5093 7285 5127
rect 7216 5059 7241 5093
rect 7275 5059 7285 5093
rect 7216 5043 7285 5059
rect 7315 5202 7367 5243
rect 7315 5168 7325 5202
rect 7359 5168 7367 5202
rect 7315 5108 7367 5168
rect 7315 5074 7325 5108
rect 7359 5074 7367 5108
rect 7315 5043 7367 5074
rect 7986 5211 8038 5249
rect 7986 5177 7994 5211
rect 8028 5177 8038 5211
rect 7986 5121 8038 5177
rect 7986 5087 7994 5121
rect 8028 5087 8038 5121
rect 7986 5049 8038 5087
rect 8068 5133 8120 5249
rect 10080 5471 10132 5509
rect 10162 5555 10214 5671
rect 11329 5555 11381 5671
rect 10162 5513 10231 5555
rect 10162 5479 10172 5513
rect 10206 5479 10231 5513
rect 10162 5471 10231 5479
rect 10261 5471 10327 5555
rect 10357 5471 10399 5555
rect 10429 5525 10495 5555
rect 10429 5491 10439 5525
rect 10473 5491 10495 5525
rect 10429 5471 10495 5491
rect 10525 5530 10584 5555
rect 10525 5496 10540 5530
rect 10574 5496 10584 5530
rect 10525 5471 10584 5496
rect 10614 5513 10668 5555
rect 10614 5479 10624 5513
rect 10658 5479 10668 5513
rect 10614 5471 10668 5479
rect 10698 5530 10752 5555
rect 10698 5496 10708 5530
rect 10742 5496 10752 5530
rect 10698 5471 10752 5496
rect 10782 5517 10834 5555
rect 10782 5483 10792 5517
rect 10826 5483 10834 5517
rect 10782 5471 10834 5483
rect 10888 5530 10940 5555
rect 10888 5496 10896 5530
rect 10930 5496 10940 5530
rect 10888 5471 10940 5496
rect 10970 5513 11024 5555
rect 10970 5479 10980 5513
rect 11014 5479 11024 5513
rect 10970 5471 11024 5479
rect 11054 5530 11108 5555
rect 11054 5496 11064 5530
rect 11098 5496 11108 5530
rect 11054 5471 11108 5496
rect 11138 5530 11192 5555
rect 11138 5496 11148 5530
rect 11182 5496 11192 5530
rect 11138 5471 11192 5496
rect 11222 5471 11282 5555
rect 11312 5521 11381 5555
rect 11312 5487 11337 5521
rect 11371 5487 11381 5521
rect 11312 5471 11381 5487
rect 11411 5630 11463 5671
rect 11411 5596 11421 5630
rect 11455 5596 11463 5630
rect 11411 5536 11463 5596
rect 11411 5502 11421 5536
rect 11455 5502 11463 5536
rect 11411 5471 11463 5502
rect 12142 5621 12194 5659
rect 12142 5587 12150 5621
rect 12184 5587 12194 5621
rect 12142 5531 12194 5587
rect 12142 5497 12150 5531
rect 12184 5497 12194 5531
rect 12142 5459 12194 5497
rect 12224 5543 12276 5659
rect 13391 5543 13443 5659
rect 12224 5501 12293 5543
rect 12224 5467 12234 5501
rect 12268 5467 12293 5501
rect 12224 5459 12293 5467
rect 12323 5459 12389 5543
rect 12419 5459 12461 5543
rect 12491 5513 12557 5543
rect 12491 5479 12501 5513
rect 12535 5479 12557 5513
rect 12491 5459 12557 5479
rect 12587 5518 12646 5543
rect 12587 5484 12602 5518
rect 12636 5484 12646 5518
rect 12587 5459 12646 5484
rect 12676 5501 12730 5543
rect 12676 5467 12686 5501
rect 12720 5467 12730 5501
rect 12676 5459 12730 5467
rect 12760 5518 12814 5543
rect 12760 5484 12770 5518
rect 12804 5484 12814 5518
rect 12760 5459 12814 5484
rect 12844 5505 12896 5543
rect 12844 5471 12854 5505
rect 12888 5471 12896 5505
rect 12844 5459 12896 5471
rect 12950 5518 13002 5543
rect 12950 5484 12958 5518
rect 12992 5484 13002 5518
rect 12950 5459 13002 5484
rect 13032 5501 13086 5543
rect 13032 5467 13042 5501
rect 13076 5467 13086 5501
rect 13032 5459 13086 5467
rect 13116 5518 13170 5543
rect 13116 5484 13126 5518
rect 13160 5484 13170 5518
rect 13116 5459 13170 5484
rect 13200 5518 13254 5543
rect 13200 5484 13210 5518
rect 13244 5484 13254 5518
rect 13200 5459 13254 5484
rect 13284 5459 13344 5543
rect 13374 5509 13443 5543
rect 13374 5475 13399 5509
rect 13433 5475 13443 5509
rect 13374 5459 13443 5475
rect 13473 5618 13525 5659
rect 13473 5584 13483 5618
rect 13517 5584 13525 5618
rect 13473 5524 13525 5584
rect 13473 5490 13483 5524
rect 13517 5490 13525 5524
rect 13473 5459 13525 5490
rect 14100 5629 14152 5667
rect 14100 5595 14108 5629
rect 14142 5595 14152 5629
rect 14100 5539 14152 5595
rect 14100 5505 14108 5539
rect 14142 5505 14152 5539
rect 14100 5467 14152 5505
rect 14182 5551 14234 5667
rect 15349 5551 15401 5667
rect 14182 5509 14251 5551
rect 14182 5475 14192 5509
rect 14226 5475 14251 5509
rect 14182 5467 14251 5475
rect 14281 5467 14347 5551
rect 14377 5467 14419 5551
rect 14449 5521 14515 5551
rect 14449 5487 14459 5521
rect 14493 5487 14515 5521
rect 14449 5467 14515 5487
rect 14545 5526 14604 5551
rect 14545 5492 14560 5526
rect 14594 5492 14604 5526
rect 14545 5467 14604 5492
rect 14634 5509 14688 5551
rect 14634 5475 14644 5509
rect 14678 5475 14688 5509
rect 14634 5467 14688 5475
rect 14718 5526 14772 5551
rect 14718 5492 14728 5526
rect 14762 5492 14772 5526
rect 14718 5467 14772 5492
rect 14802 5513 14854 5551
rect 14802 5479 14812 5513
rect 14846 5479 14854 5513
rect 14802 5467 14854 5479
rect 14908 5526 14960 5551
rect 14908 5492 14916 5526
rect 14950 5492 14960 5526
rect 14908 5467 14960 5492
rect 14990 5509 15044 5551
rect 14990 5475 15000 5509
rect 15034 5475 15044 5509
rect 14990 5467 15044 5475
rect 15074 5526 15128 5551
rect 15074 5492 15084 5526
rect 15118 5492 15128 5526
rect 15074 5467 15128 5492
rect 15158 5526 15212 5551
rect 15158 5492 15168 5526
rect 15202 5492 15212 5526
rect 15158 5467 15212 5492
rect 15242 5467 15302 5551
rect 15332 5517 15401 5551
rect 15332 5483 15357 5517
rect 15391 5483 15401 5517
rect 15332 5467 15401 5483
rect 15431 5626 15483 5667
rect 15431 5592 15441 5626
rect 15475 5592 15483 5626
rect 15431 5532 15483 5592
rect 15431 5498 15441 5532
rect 15475 5498 15483 5532
rect 15431 5467 15483 5498
rect 16094 5635 16146 5673
rect 16094 5601 16102 5635
rect 16136 5601 16146 5635
rect 16094 5545 16146 5601
rect 16094 5511 16102 5545
rect 16136 5511 16146 5545
rect 16094 5473 16146 5511
rect 16176 5557 16228 5673
rect 17343 5557 17395 5673
rect 16176 5515 16245 5557
rect 16176 5481 16186 5515
rect 16220 5481 16245 5515
rect 16176 5473 16245 5481
rect 16275 5473 16341 5557
rect 16371 5473 16413 5557
rect 16443 5527 16509 5557
rect 16443 5493 16453 5527
rect 16487 5493 16509 5527
rect 16443 5473 16509 5493
rect 16539 5532 16598 5557
rect 16539 5498 16554 5532
rect 16588 5498 16598 5532
rect 16539 5473 16598 5498
rect 16628 5515 16682 5557
rect 16628 5481 16638 5515
rect 16672 5481 16682 5515
rect 16628 5473 16682 5481
rect 16712 5532 16766 5557
rect 16712 5498 16722 5532
rect 16756 5498 16766 5532
rect 16712 5473 16766 5498
rect 16796 5519 16848 5557
rect 16796 5485 16806 5519
rect 16840 5485 16848 5519
rect 16796 5473 16848 5485
rect 16902 5532 16954 5557
rect 16902 5498 16910 5532
rect 16944 5498 16954 5532
rect 16902 5473 16954 5498
rect 16984 5515 17038 5557
rect 16984 5481 16994 5515
rect 17028 5481 17038 5515
rect 16984 5473 17038 5481
rect 17068 5532 17122 5557
rect 17068 5498 17078 5532
rect 17112 5498 17122 5532
rect 17068 5473 17122 5498
rect 17152 5532 17206 5557
rect 17152 5498 17162 5532
rect 17196 5498 17206 5532
rect 17152 5473 17206 5498
rect 17236 5473 17296 5557
rect 17326 5523 17395 5557
rect 17326 5489 17351 5523
rect 17385 5489 17395 5523
rect 17326 5473 17395 5489
rect 17425 5632 17477 5673
rect 17425 5598 17435 5632
rect 17469 5598 17477 5632
rect 17425 5538 17477 5598
rect 17425 5504 17435 5538
rect 17469 5504 17477 5538
rect 17425 5473 17477 5504
rect 9235 5133 9287 5249
rect 8068 5091 8137 5133
rect 8068 5057 8078 5091
rect 8112 5057 8137 5091
rect 8068 5049 8137 5057
rect 8167 5049 8233 5133
rect 8263 5049 8305 5133
rect 8335 5103 8401 5133
rect 8335 5069 8345 5103
rect 8379 5069 8401 5103
rect 8335 5049 8401 5069
rect 8431 5108 8490 5133
rect 8431 5074 8446 5108
rect 8480 5074 8490 5108
rect 8431 5049 8490 5074
rect 8520 5091 8574 5133
rect 8520 5057 8530 5091
rect 8564 5057 8574 5091
rect 8520 5049 8574 5057
rect 8604 5108 8658 5133
rect 8604 5074 8614 5108
rect 8648 5074 8658 5108
rect 8604 5049 8658 5074
rect 8688 5095 8740 5133
rect 8688 5061 8698 5095
rect 8732 5061 8740 5095
rect 8688 5049 8740 5061
rect 8794 5108 8846 5133
rect 8794 5074 8802 5108
rect 8836 5074 8846 5108
rect 8794 5049 8846 5074
rect 8876 5091 8930 5133
rect 8876 5057 8886 5091
rect 8920 5057 8930 5091
rect 8876 5049 8930 5057
rect 8960 5108 9014 5133
rect 8960 5074 8970 5108
rect 9004 5074 9014 5108
rect 8960 5049 9014 5074
rect 9044 5108 9098 5133
rect 9044 5074 9054 5108
rect 9088 5074 9098 5108
rect 9044 5049 9098 5074
rect 9128 5049 9188 5133
rect 9218 5099 9287 5133
rect 9218 5065 9243 5099
rect 9277 5065 9287 5099
rect 9218 5049 9287 5065
rect 9317 5208 9369 5249
rect 9317 5174 9327 5208
rect 9361 5174 9369 5208
rect 9317 5114 9369 5174
rect 9317 5080 9327 5114
rect 9361 5080 9369 5114
rect 9317 5049 9369 5080
rect 10108 4759 10160 4797
rect 10108 4725 10116 4759
rect 10150 4725 10160 4759
rect 10108 4669 10160 4725
rect 10108 4635 10116 4669
rect 10150 4635 10160 4669
rect 10108 4597 10160 4635
rect 10190 4681 10242 4797
rect 11357 4681 11409 4797
rect 10190 4639 10259 4681
rect 10190 4605 10200 4639
rect 10234 4605 10259 4639
rect 10190 4597 10259 4605
rect 10289 4597 10355 4681
rect 10385 4597 10427 4681
rect 10457 4651 10523 4681
rect 10457 4617 10467 4651
rect 10501 4617 10523 4651
rect 10457 4597 10523 4617
rect 10553 4656 10612 4681
rect 10553 4622 10568 4656
rect 10602 4622 10612 4656
rect 10553 4597 10612 4622
rect 10642 4639 10696 4681
rect 10642 4605 10652 4639
rect 10686 4605 10696 4639
rect 10642 4597 10696 4605
rect 10726 4656 10780 4681
rect 10726 4622 10736 4656
rect 10770 4622 10780 4656
rect 10726 4597 10780 4622
rect 10810 4643 10862 4681
rect 10810 4609 10820 4643
rect 10854 4609 10862 4643
rect 10810 4597 10862 4609
rect 10916 4656 10968 4681
rect 10916 4622 10924 4656
rect 10958 4622 10968 4656
rect 10916 4597 10968 4622
rect 10998 4639 11052 4681
rect 10998 4605 11008 4639
rect 11042 4605 11052 4639
rect 10998 4597 11052 4605
rect 11082 4656 11136 4681
rect 11082 4622 11092 4656
rect 11126 4622 11136 4656
rect 11082 4597 11136 4622
rect 11166 4656 11220 4681
rect 11166 4622 11176 4656
rect 11210 4622 11220 4656
rect 11166 4597 11220 4622
rect 11250 4597 11310 4681
rect 11340 4647 11409 4681
rect 11340 4613 11365 4647
rect 11399 4613 11409 4647
rect 11340 4597 11409 4613
rect 11439 4756 11491 4797
rect 11439 4722 11449 4756
rect 11483 4722 11491 4756
rect 11439 4662 11491 4722
rect 11439 4628 11449 4662
rect 11483 4628 11491 4662
rect 11439 4597 11491 4628
rect 12378 4715 12430 4753
rect 12378 4681 12386 4715
rect 12420 4681 12430 4715
rect 12378 4625 12430 4681
rect 12378 4591 12386 4625
rect 12420 4591 12430 4625
rect 12378 4553 12430 4591
rect 12460 4637 12512 4753
rect 13627 4637 13679 4753
rect 12460 4595 12529 4637
rect 12460 4561 12470 4595
rect 12504 4561 12529 4595
rect 12460 4553 12529 4561
rect 12559 4553 12625 4637
rect 12655 4553 12697 4637
rect 12727 4607 12793 4637
rect 12727 4573 12737 4607
rect 12771 4573 12793 4607
rect 12727 4553 12793 4573
rect 12823 4612 12882 4637
rect 12823 4578 12838 4612
rect 12872 4578 12882 4612
rect 12823 4553 12882 4578
rect 12912 4595 12966 4637
rect 12912 4561 12922 4595
rect 12956 4561 12966 4595
rect 12912 4553 12966 4561
rect 12996 4612 13050 4637
rect 12996 4578 13006 4612
rect 13040 4578 13050 4612
rect 12996 4553 13050 4578
rect 13080 4599 13132 4637
rect 13080 4565 13090 4599
rect 13124 4565 13132 4599
rect 13080 4553 13132 4565
rect 13186 4612 13238 4637
rect 13186 4578 13194 4612
rect 13228 4578 13238 4612
rect 13186 4553 13238 4578
rect 13268 4595 13322 4637
rect 13268 4561 13278 4595
rect 13312 4561 13322 4595
rect 13268 4553 13322 4561
rect 13352 4612 13406 4637
rect 13352 4578 13362 4612
rect 13396 4578 13406 4612
rect 13352 4553 13406 4578
rect 13436 4612 13490 4637
rect 13436 4578 13446 4612
rect 13480 4578 13490 4612
rect 13436 4553 13490 4578
rect 13520 4553 13580 4637
rect 13610 4603 13679 4637
rect 13610 4569 13635 4603
rect 13669 4569 13679 4603
rect 13610 4553 13679 4569
rect 13709 4712 13761 4753
rect 13709 4678 13719 4712
rect 13753 4678 13761 4712
rect 13709 4618 13761 4678
rect 13709 4584 13719 4618
rect 13753 4584 13761 4618
rect 13709 4553 13761 4584
rect 14380 4709 14432 4747
rect 14380 4675 14388 4709
rect 14422 4675 14432 4709
rect 14380 4619 14432 4675
rect 14380 4585 14388 4619
rect 14422 4585 14432 4619
rect 14380 4547 14432 4585
rect 14462 4631 14514 4747
rect 15629 4631 15681 4747
rect 14462 4589 14531 4631
rect 14462 4555 14472 4589
rect 14506 4555 14531 4589
rect 14462 4547 14531 4555
rect 14561 4547 14627 4631
rect 14657 4547 14699 4631
rect 14729 4601 14795 4631
rect 14729 4567 14739 4601
rect 14773 4567 14795 4601
rect 14729 4547 14795 4567
rect 14825 4606 14884 4631
rect 14825 4572 14840 4606
rect 14874 4572 14884 4606
rect 14825 4547 14884 4572
rect 14914 4589 14968 4631
rect 14914 4555 14924 4589
rect 14958 4555 14968 4589
rect 14914 4547 14968 4555
rect 14998 4606 15052 4631
rect 14998 4572 15008 4606
rect 15042 4572 15052 4606
rect 14998 4547 15052 4572
rect 15082 4593 15134 4631
rect 15082 4559 15092 4593
rect 15126 4559 15134 4593
rect 15082 4547 15134 4559
rect 15188 4606 15240 4631
rect 15188 4572 15196 4606
rect 15230 4572 15240 4606
rect 15188 4547 15240 4572
rect 15270 4589 15324 4631
rect 15270 4555 15280 4589
rect 15314 4555 15324 4589
rect 15270 4547 15324 4555
rect 15354 4606 15408 4631
rect 15354 4572 15364 4606
rect 15398 4572 15408 4606
rect 15354 4547 15408 4572
rect 15438 4606 15492 4631
rect 15438 4572 15448 4606
rect 15482 4572 15492 4606
rect 15438 4547 15492 4572
rect 15522 4547 15582 4631
rect 15612 4597 15681 4631
rect 15612 4563 15637 4597
rect 15671 4563 15681 4597
rect 15612 4547 15681 4563
rect 15711 4706 15763 4747
rect 15711 4672 15721 4706
rect 15755 4672 15763 4706
rect 15711 4612 15763 4672
rect 15711 4578 15721 4612
rect 15755 4578 15763 4612
rect 15711 4547 15763 4578
rect 16402 4691 16454 4729
rect 16402 4657 16410 4691
rect 16444 4657 16454 4691
rect 16402 4601 16454 4657
rect 16402 4567 16410 4601
rect 16444 4567 16454 4601
rect 16402 4529 16454 4567
rect 16484 4613 16536 4729
rect 17651 4613 17703 4729
rect 16484 4571 16553 4613
rect 16484 4537 16494 4571
rect 16528 4537 16553 4571
rect 16484 4529 16553 4537
rect 16583 4529 16649 4613
rect 16679 4529 16721 4613
rect 16751 4583 16817 4613
rect 16751 4549 16761 4583
rect 16795 4549 16817 4583
rect 16751 4529 16817 4549
rect 16847 4588 16906 4613
rect 16847 4554 16862 4588
rect 16896 4554 16906 4588
rect 16847 4529 16906 4554
rect 16936 4571 16990 4613
rect 16936 4537 16946 4571
rect 16980 4537 16990 4571
rect 16936 4529 16990 4537
rect 17020 4588 17074 4613
rect 17020 4554 17030 4588
rect 17064 4554 17074 4588
rect 17020 4529 17074 4554
rect 17104 4575 17156 4613
rect 17104 4541 17114 4575
rect 17148 4541 17156 4575
rect 17104 4529 17156 4541
rect 17210 4588 17262 4613
rect 17210 4554 17218 4588
rect 17252 4554 17262 4588
rect 17210 4529 17262 4554
rect 17292 4571 17346 4613
rect 17292 4537 17302 4571
rect 17336 4537 17346 4571
rect 17292 4529 17346 4537
rect 17376 4588 17430 4613
rect 17376 4554 17386 4588
rect 17420 4554 17430 4588
rect 17376 4529 17430 4554
rect 17460 4588 17514 4613
rect 17460 4554 17470 4588
rect 17504 4554 17514 4588
rect 17460 4529 17514 4554
rect 17544 4529 17604 4613
rect 17634 4579 17703 4613
rect 17634 4545 17659 4579
rect 17693 4545 17703 4579
rect 17634 4529 17703 4545
rect 17733 4688 17785 4729
rect 17733 4654 17743 4688
rect 17777 4654 17785 4688
rect 17733 4594 17785 4654
rect 17733 4560 17743 4594
rect 17777 4560 17785 4594
rect 17733 4529 17785 4560
rect 1868 1953 1920 1991
rect 1868 1919 1876 1953
rect 1910 1919 1920 1953
rect 1868 1863 1920 1919
rect 1868 1829 1876 1863
rect 1910 1829 1920 1863
rect 1868 1791 1920 1829
rect 1950 1875 2002 1991
rect 3117 1875 3169 1991
rect 1950 1833 2019 1875
rect 1950 1799 1960 1833
rect 1994 1799 2019 1833
rect 1950 1791 2019 1799
rect 2049 1791 2115 1875
rect 2145 1791 2187 1875
rect 2217 1845 2283 1875
rect 2217 1811 2227 1845
rect 2261 1811 2283 1845
rect 2217 1791 2283 1811
rect 2313 1850 2372 1875
rect 2313 1816 2328 1850
rect 2362 1816 2372 1850
rect 2313 1791 2372 1816
rect 2402 1833 2456 1875
rect 2402 1799 2412 1833
rect 2446 1799 2456 1833
rect 2402 1791 2456 1799
rect 2486 1850 2540 1875
rect 2486 1816 2496 1850
rect 2530 1816 2540 1850
rect 2486 1791 2540 1816
rect 2570 1837 2622 1875
rect 2570 1803 2580 1837
rect 2614 1803 2622 1837
rect 2570 1791 2622 1803
rect 2676 1850 2728 1875
rect 2676 1816 2684 1850
rect 2718 1816 2728 1850
rect 2676 1791 2728 1816
rect 2758 1833 2812 1875
rect 2758 1799 2768 1833
rect 2802 1799 2812 1833
rect 2758 1791 2812 1799
rect 2842 1850 2896 1875
rect 2842 1816 2852 1850
rect 2886 1816 2896 1850
rect 2842 1791 2896 1816
rect 2926 1850 2980 1875
rect 2926 1816 2936 1850
rect 2970 1816 2980 1850
rect 2926 1791 2980 1816
rect 3010 1791 3070 1875
rect 3100 1841 3169 1875
rect 3100 1807 3125 1841
rect 3159 1807 3169 1841
rect 3100 1791 3169 1807
rect 3199 1950 3251 1991
rect 3199 1916 3209 1950
rect 3243 1916 3251 1950
rect 3199 1856 3251 1916
rect 3199 1822 3209 1856
rect 3243 1822 3251 1856
rect 3199 1791 3251 1822
rect 3938 1949 3990 1987
rect 3938 1915 3946 1949
rect 3980 1915 3990 1949
rect 3938 1859 3990 1915
rect 3938 1825 3946 1859
rect 3980 1825 3990 1859
rect 3938 1787 3990 1825
rect 4020 1871 4072 1987
rect 5187 1871 5239 1987
rect 4020 1829 4089 1871
rect 4020 1795 4030 1829
rect 4064 1795 4089 1829
rect 4020 1787 4089 1795
rect 4119 1787 4185 1871
rect 4215 1787 4257 1871
rect 4287 1841 4353 1871
rect 4287 1807 4297 1841
rect 4331 1807 4353 1841
rect 4287 1787 4353 1807
rect 4383 1846 4442 1871
rect 4383 1812 4398 1846
rect 4432 1812 4442 1846
rect 4383 1787 4442 1812
rect 4472 1829 4526 1871
rect 4472 1795 4482 1829
rect 4516 1795 4526 1829
rect 4472 1787 4526 1795
rect 4556 1846 4610 1871
rect 4556 1812 4566 1846
rect 4600 1812 4610 1846
rect 4556 1787 4610 1812
rect 4640 1833 4692 1871
rect 4640 1799 4650 1833
rect 4684 1799 4692 1833
rect 4640 1787 4692 1799
rect 4746 1846 4798 1871
rect 4746 1812 4754 1846
rect 4788 1812 4798 1846
rect 4746 1787 4798 1812
rect 4828 1829 4882 1871
rect 4828 1795 4838 1829
rect 4872 1795 4882 1829
rect 4828 1787 4882 1795
rect 4912 1846 4966 1871
rect 4912 1812 4922 1846
rect 4956 1812 4966 1846
rect 4912 1787 4966 1812
rect 4996 1846 5050 1871
rect 4996 1812 5006 1846
rect 5040 1812 5050 1846
rect 4996 1787 5050 1812
rect 5080 1787 5140 1871
rect 5170 1837 5239 1871
rect 5170 1803 5195 1837
rect 5229 1803 5239 1837
rect 5170 1787 5239 1803
rect 5269 1946 5321 1987
rect 5269 1912 5279 1946
rect 5313 1912 5321 1946
rect 5269 1852 5321 1912
rect 5269 1818 5279 1852
rect 5313 1818 5321 1852
rect 5269 1787 5321 1818
rect 5890 1949 5942 1987
rect 5890 1915 5898 1949
rect 5932 1915 5942 1949
rect 5890 1859 5942 1915
rect 5890 1825 5898 1859
rect 5932 1825 5942 1859
rect 5890 1787 5942 1825
rect 5972 1871 6024 1987
rect 7139 1871 7191 1987
rect 5972 1829 6041 1871
rect 5972 1795 5982 1829
rect 6016 1795 6041 1829
rect 5972 1787 6041 1795
rect 6071 1787 6137 1871
rect 6167 1787 6209 1871
rect 6239 1841 6305 1871
rect 6239 1807 6249 1841
rect 6283 1807 6305 1841
rect 6239 1787 6305 1807
rect 6335 1846 6394 1871
rect 6335 1812 6350 1846
rect 6384 1812 6394 1846
rect 6335 1787 6394 1812
rect 6424 1829 6478 1871
rect 6424 1795 6434 1829
rect 6468 1795 6478 1829
rect 6424 1787 6478 1795
rect 6508 1846 6562 1871
rect 6508 1812 6518 1846
rect 6552 1812 6562 1846
rect 6508 1787 6562 1812
rect 6592 1833 6644 1871
rect 6592 1799 6602 1833
rect 6636 1799 6644 1833
rect 6592 1787 6644 1799
rect 6698 1846 6750 1871
rect 6698 1812 6706 1846
rect 6740 1812 6750 1846
rect 6698 1787 6750 1812
rect 6780 1829 6834 1871
rect 6780 1795 6790 1829
rect 6824 1795 6834 1829
rect 6780 1787 6834 1795
rect 6864 1846 6918 1871
rect 6864 1812 6874 1846
rect 6908 1812 6918 1846
rect 6864 1787 6918 1812
rect 6948 1846 7002 1871
rect 6948 1812 6958 1846
rect 6992 1812 7002 1846
rect 6948 1787 7002 1812
rect 7032 1787 7092 1871
rect 7122 1837 7191 1871
rect 7122 1803 7147 1837
rect 7181 1803 7191 1837
rect 7122 1787 7191 1803
rect 7221 1946 7273 1987
rect 7221 1912 7231 1946
rect 7265 1912 7273 1946
rect 7221 1852 7273 1912
rect 7221 1818 7231 1852
rect 7265 1818 7273 1852
rect 7221 1787 7273 1818
rect 7892 1955 7944 1993
rect 7892 1921 7900 1955
rect 7934 1921 7944 1955
rect 7892 1865 7944 1921
rect 7892 1831 7900 1865
rect 7934 1831 7944 1865
rect 7892 1793 7944 1831
rect 7974 1877 8026 1993
rect 9141 1877 9193 1993
rect 7974 1835 8043 1877
rect 7974 1801 7984 1835
rect 8018 1801 8043 1835
rect 7974 1793 8043 1801
rect 8073 1793 8139 1877
rect 8169 1793 8211 1877
rect 8241 1847 8307 1877
rect 8241 1813 8251 1847
rect 8285 1813 8307 1847
rect 8241 1793 8307 1813
rect 8337 1852 8396 1877
rect 8337 1818 8352 1852
rect 8386 1818 8396 1852
rect 8337 1793 8396 1818
rect 8426 1835 8480 1877
rect 8426 1801 8436 1835
rect 8470 1801 8480 1835
rect 8426 1793 8480 1801
rect 8510 1852 8564 1877
rect 8510 1818 8520 1852
rect 8554 1818 8564 1852
rect 8510 1793 8564 1818
rect 8594 1839 8646 1877
rect 8594 1805 8604 1839
rect 8638 1805 8646 1839
rect 8594 1793 8646 1805
rect 8700 1852 8752 1877
rect 8700 1818 8708 1852
rect 8742 1818 8752 1852
rect 8700 1793 8752 1818
rect 8782 1835 8836 1877
rect 8782 1801 8792 1835
rect 8826 1801 8836 1835
rect 8782 1793 8836 1801
rect 8866 1852 8920 1877
rect 8866 1818 8876 1852
rect 8910 1818 8920 1852
rect 8866 1793 8920 1818
rect 8950 1852 9004 1877
rect 8950 1818 8960 1852
rect 8994 1818 9004 1852
rect 8950 1793 9004 1818
rect 9034 1793 9094 1877
rect 9124 1843 9193 1877
rect 9124 1809 9149 1843
rect 9183 1809 9193 1843
rect 9124 1793 9193 1809
rect 9223 1952 9275 1993
rect 9223 1918 9233 1952
rect 9267 1918 9275 1952
rect 9223 1858 9275 1918
rect 9223 1824 9233 1858
rect 9267 1824 9275 1858
rect 9223 1793 9275 1824
rect 9844 1955 9896 1993
rect 9844 1921 9852 1955
rect 9886 1921 9896 1955
rect 9844 1865 9896 1921
rect 9844 1831 9852 1865
rect 9886 1831 9896 1865
rect 9844 1793 9896 1831
rect 9926 1877 9978 1993
rect 11093 1877 11145 1993
rect 9926 1835 9995 1877
rect 9926 1801 9936 1835
rect 9970 1801 9995 1835
rect 9926 1793 9995 1801
rect 10025 1793 10091 1877
rect 10121 1793 10163 1877
rect 10193 1847 10259 1877
rect 10193 1813 10203 1847
rect 10237 1813 10259 1847
rect 10193 1793 10259 1813
rect 10289 1852 10348 1877
rect 10289 1818 10304 1852
rect 10338 1818 10348 1852
rect 10289 1793 10348 1818
rect 10378 1835 10432 1877
rect 10378 1801 10388 1835
rect 10422 1801 10432 1835
rect 10378 1793 10432 1801
rect 10462 1852 10516 1877
rect 10462 1818 10472 1852
rect 10506 1818 10516 1852
rect 10462 1793 10516 1818
rect 10546 1839 10598 1877
rect 10546 1805 10556 1839
rect 10590 1805 10598 1839
rect 10546 1793 10598 1805
rect 10652 1852 10704 1877
rect 10652 1818 10660 1852
rect 10694 1818 10704 1852
rect 10652 1793 10704 1818
rect 10734 1835 10788 1877
rect 10734 1801 10744 1835
rect 10778 1801 10788 1835
rect 10734 1793 10788 1801
rect 10818 1852 10872 1877
rect 10818 1818 10828 1852
rect 10862 1818 10872 1852
rect 10818 1793 10872 1818
rect 10902 1852 10956 1877
rect 10902 1818 10912 1852
rect 10946 1818 10956 1852
rect 10902 1793 10956 1818
rect 10986 1793 11046 1877
rect 11076 1843 11145 1877
rect 11076 1809 11101 1843
rect 11135 1809 11145 1843
rect 11076 1793 11145 1809
rect 11175 1952 11227 1993
rect 11175 1918 11185 1952
rect 11219 1918 11227 1952
rect 11175 1858 11227 1918
rect 11175 1824 11185 1858
rect 11219 1824 11227 1858
rect 11175 1793 11227 1824
rect 11836 1955 11888 1993
rect 11836 1921 11844 1955
rect 11878 1921 11888 1955
rect 11836 1865 11888 1921
rect 11836 1831 11844 1865
rect 11878 1831 11888 1865
rect 11836 1793 11888 1831
rect 11918 1877 11970 1993
rect 13085 1877 13137 1993
rect 11918 1835 11987 1877
rect 11918 1801 11928 1835
rect 11962 1801 11987 1835
rect 11918 1793 11987 1801
rect 12017 1793 12083 1877
rect 12113 1793 12155 1877
rect 12185 1847 12251 1877
rect 12185 1813 12195 1847
rect 12229 1813 12251 1847
rect 12185 1793 12251 1813
rect 12281 1852 12340 1877
rect 12281 1818 12296 1852
rect 12330 1818 12340 1852
rect 12281 1793 12340 1818
rect 12370 1835 12424 1877
rect 12370 1801 12380 1835
rect 12414 1801 12424 1835
rect 12370 1793 12424 1801
rect 12454 1852 12508 1877
rect 12454 1818 12464 1852
rect 12498 1818 12508 1852
rect 12454 1793 12508 1818
rect 12538 1839 12590 1877
rect 12538 1805 12548 1839
rect 12582 1805 12590 1839
rect 12538 1793 12590 1805
rect 12644 1852 12696 1877
rect 12644 1818 12652 1852
rect 12686 1818 12696 1852
rect 12644 1793 12696 1818
rect 12726 1835 12780 1877
rect 12726 1801 12736 1835
rect 12770 1801 12780 1835
rect 12726 1793 12780 1801
rect 12810 1852 12864 1877
rect 12810 1818 12820 1852
rect 12854 1818 12864 1852
rect 12810 1793 12864 1818
rect 12894 1852 12948 1877
rect 12894 1818 12904 1852
rect 12938 1818 12948 1852
rect 12894 1793 12948 1818
rect 12978 1793 13038 1877
rect 13068 1843 13137 1877
rect 13068 1809 13093 1843
rect 13127 1809 13137 1843
rect 13068 1793 13137 1809
rect 13167 1952 13219 1993
rect 13167 1918 13177 1952
rect 13211 1918 13219 1952
rect 13167 1858 13219 1918
rect 13167 1824 13177 1858
rect 13211 1824 13219 1858
rect 13167 1793 13219 1824
rect 13788 1955 13840 1993
rect 13788 1921 13796 1955
rect 13830 1921 13840 1955
rect 13788 1865 13840 1921
rect 13788 1831 13796 1865
rect 13830 1831 13840 1865
rect 13788 1793 13840 1831
rect 13870 1877 13922 1993
rect 15037 1877 15089 1993
rect 13870 1835 13939 1877
rect 13870 1801 13880 1835
rect 13914 1801 13939 1835
rect 13870 1793 13939 1801
rect 13969 1793 14035 1877
rect 14065 1793 14107 1877
rect 14137 1847 14203 1877
rect 14137 1813 14147 1847
rect 14181 1813 14203 1847
rect 14137 1793 14203 1813
rect 14233 1852 14292 1877
rect 14233 1818 14248 1852
rect 14282 1818 14292 1852
rect 14233 1793 14292 1818
rect 14322 1835 14376 1877
rect 14322 1801 14332 1835
rect 14366 1801 14376 1835
rect 14322 1793 14376 1801
rect 14406 1852 14460 1877
rect 14406 1818 14416 1852
rect 14450 1818 14460 1852
rect 14406 1793 14460 1818
rect 14490 1839 14542 1877
rect 14490 1805 14500 1839
rect 14534 1805 14542 1839
rect 14490 1793 14542 1805
rect 14596 1852 14648 1877
rect 14596 1818 14604 1852
rect 14638 1818 14648 1852
rect 14596 1793 14648 1818
rect 14678 1835 14732 1877
rect 14678 1801 14688 1835
rect 14722 1801 14732 1835
rect 14678 1793 14732 1801
rect 14762 1852 14816 1877
rect 14762 1818 14772 1852
rect 14806 1818 14816 1852
rect 14762 1793 14816 1818
rect 14846 1852 14900 1877
rect 14846 1818 14856 1852
rect 14890 1818 14900 1852
rect 14846 1793 14900 1818
rect 14930 1793 14990 1877
rect 15020 1843 15089 1877
rect 15020 1809 15045 1843
rect 15079 1809 15089 1843
rect 15020 1793 15089 1809
rect 15119 1952 15171 1993
rect 15119 1918 15129 1952
rect 15163 1918 15171 1952
rect 15119 1858 15171 1918
rect 15119 1824 15129 1858
rect 15163 1824 15171 1858
rect 15119 1793 15171 1824
rect 15852 1955 15904 1993
rect 15852 1921 15860 1955
rect 15894 1921 15904 1955
rect 15852 1865 15904 1921
rect 15852 1831 15860 1865
rect 15894 1831 15904 1865
rect 15852 1793 15904 1831
rect 15934 1877 15986 1993
rect 17101 1877 17153 1993
rect 15934 1835 16003 1877
rect 15934 1801 15944 1835
rect 15978 1801 16003 1835
rect 15934 1793 16003 1801
rect 16033 1793 16099 1877
rect 16129 1793 16171 1877
rect 16201 1847 16267 1877
rect 16201 1813 16211 1847
rect 16245 1813 16267 1847
rect 16201 1793 16267 1813
rect 16297 1852 16356 1877
rect 16297 1818 16312 1852
rect 16346 1818 16356 1852
rect 16297 1793 16356 1818
rect 16386 1835 16440 1877
rect 16386 1801 16396 1835
rect 16430 1801 16440 1835
rect 16386 1793 16440 1801
rect 16470 1852 16524 1877
rect 16470 1818 16480 1852
rect 16514 1818 16524 1852
rect 16470 1793 16524 1818
rect 16554 1839 16606 1877
rect 16554 1805 16564 1839
rect 16598 1805 16606 1839
rect 16554 1793 16606 1805
rect 16660 1852 16712 1877
rect 16660 1818 16668 1852
rect 16702 1818 16712 1852
rect 16660 1793 16712 1818
rect 16742 1835 16796 1877
rect 16742 1801 16752 1835
rect 16786 1801 16796 1835
rect 16742 1793 16796 1801
rect 16826 1852 16880 1877
rect 16826 1818 16836 1852
rect 16870 1818 16880 1852
rect 16826 1793 16880 1818
rect 16910 1852 16964 1877
rect 16910 1818 16920 1852
rect 16954 1818 16964 1852
rect 16910 1793 16964 1818
rect 16994 1793 17054 1877
rect 17084 1843 17153 1877
rect 17084 1809 17109 1843
rect 17143 1809 17153 1843
rect 17084 1793 17153 1809
rect 17183 1952 17235 1993
rect 17183 1918 17193 1952
rect 17227 1918 17235 1952
rect 17183 1858 17235 1918
rect 17183 1824 17193 1858
rect 17227 1824 17235 1858
rect 17183 1793 17235 1824
<< ndiffc >>
rect 18879 35065 18913 35099
rect 18917 34981 18951 35015
rect 18891 34886 18925 34920
rect 18846 34782 18880 34816
rect 18914 34782 18948 34816
rect 18887 34698 18921 34732
rect 18848 34614 18882 34648
rect 18916 34614 18950 34648
rect 18903 34508 18937 34542
rect 18903 34310 18937 34344
rect 18903 34207 18937 34241
rect 18909 34088 18943 34122
rect 18903 33889 18937 33923
rect 18903 33778 18937 33812
rect 18917 33693 18951 33727
rect 18891 33589 18925 33623
rect 18917 33505 18951 33539
rect 18891 33421 18925 33455
rect 18887 32759 18921 32793
rect 18925 32675 18959 32709
rect 18899 32580 18933 32614
rect 18854 32476 18888 32510
rect 18922 32476 18956 32510
rect 18895 32392 18929 32426
rect 18856 32308 18890 32342
rect 18924 32308 18958 32342
rect 18911 32202 18945 32236
rect 18911 32004 18945 32038
rect 18911 31901 18945 31935
rect 18917 31782 18951 31816
rect 18911 31583 18945 31617
rect 18911 31472 18945 31506
rect 18925 31387 18959 31421
rect 18899 31283 18933 31317
rect 18925 31199 18959 31233
rect 18899 31115 18933 31149
rect 18895 30545 18929 30579
rect 18933 30461 18967 30495
rect 18907 30366 18941 30400
rect 18862 30262 18896 30296
rect 18930 30262 18964 30296
rect 18903 30178 18937 30212
rect 18864 30094 18898 30128
rect 18932 30094 18966 30128
rect 18919 29988 18953 30022
rect 18919 29790 18953 29824
rect 18919 29687 18953 29721
rect 18925 29568 18959 29602
rect 18919 29369 18953 29403
rect 18919 29258 18953 29292
rect 18933 29173 18967 29207
rect 18907 29069 18941 29103
rect 18933 28985 18967 29019
rect 18907 28901 18941 28935
rect 18877 28345 18911 28379
rect 18915 28261 18949 28295
rect 18889 28166 18923 28200
rect 18844 28062 18878 28096
rect 18912 28062 18946 28096
rect 18885 27978 18919 28012
rect 18846 27894 18880 27928
rect 18914 27894 18948 27928
rect 18901 27788 18935 27822
rect 18901 27590 18935 27624
rect 18901 27487 18935 27521
rect 18907 27368 18941 27402
rect 18901 27169 18935 27203
rect 18901 27058 18935 27092
rect 18915 26973 18949 27007
rect 18889 26869 18923 26903
rect 18915 26785 18949 26819
rect 18889 26701 18923 26735
rect 18885 26131 18919 26165
rect 18923 26047 18957 26081
rect 18897 25952 18931 25986
rect 18852 25848 18886 25882
rect 18920 25848 18954 25882
rect 18893 25764 18927 25798
rect 18854 25680 18888 25714
rect 18922 25680 18956 25714
rect 18909 25574 18943 25608
rect 18909 25376 18943 25410
rect 18909 25273 18943 25307
rect 18915 25154 18949 25188
rect 18909 24955 18943 24989
rect 18909 24844 18943 24878
rect 18923 24759 18957 24793
rect 18897 24655 18931 24689
rect 18923 24571 18957 24605
rect 18897 24487 18931 24521
rect 7581 22929 7615 22963
rect 7665 22903 7699 22937
rect 7749 22929 7783 22963
rect 7853 22903 7887 22937
rect 7938 22917 7972 22951
rect 8049 22917 8083 22951
rect 8248 22911 8282 22945
rect 8367 22917 8401 22951
rect 8470 22917 8504 22951
rect 8668 22917 8702 22951
rect 8774 22972 8808 23006
rect 8774 22904 8808 22938
rect 8858 22933 8892 22967
rect 8942 22974 8976 23008
rect 8942 22906 8976 22940
rect 9046 22929 9080 22963
rect 9141 22903 9175 22937
rect 9225 22941 9259 22975
rect 9795 22937 9829 22971
rect 9879 22911 9913 22945
rect 9963 22937 9997 22971
rect 10067 22911 10101 22945
rect 10152 22925 10186 22959
rect 10263 22925 10297 22959
rect 10462 22919 10496 22953
rect 10581 22925 10615 22959
rect 10684 22925 10718 22959
rect 10882 22925 10916 22959
rect 10988 22980 11022 23014
rect 10988 22912 11022 22946
rect 11072 22941 11106 22975
rect 11156 22982 11190 23016
rect 11156 22914 11190 22948
rect 11260 22937 11294 22971
rect 11355 22911 11389 22945
rect 11439 22949 11473 22983
rect 11995 22919 12029 22953
rect 12079 22893 12113 22927
rect 12163 22919 12197 22953
rect 12267 22893 12301 22927
rect 12352 22907 12386 22941
rect 12463 22907 12497 22941
rect 12662 22901 12696 22935
rect 12781 22907 12815 22941
rect 12884 22907 12918 22941
rect 13082 22907 13116 22941
rect 13188 22962 13222 22996
rect 13188 22894 13222 22928
rect 13272 22923 13306 22957
rect 13356 22964 13390 22998
rect 13356 22896 13390 22930
rect 13460 22919 13494 22953
rect 13555 22893 13589 22927
rect 13639 22931 13673 22965
rect 14209 22927 14243 22961
rect 14293 22901 14327 22935
rect 14377 22927 14411 22961
rect 14481 22901 14515 22935
rect 14566 22915 14600 22949
rect 14677 22915 14711 22949
rect 14876 22909 14910 22943
rect 14995 22915 15029 22949
rect 15098 22915 15132 22949
rect 15296 22915 15330 22949
rect 15402 22970 15436 23004
rect 15402 22902 15436 22936
rect 15486 22931 15520 22965
rect 15570 22972 15604 23006
rect 15570 22904 15604 22938
rect 15674 22927 15708 22961
rect 15769 22901 15803 22935
rect 15853 22939 15887 22973
rect 16515 22935 16549 22969
rect 16599 22909 16633 22943
rect 16683 22935 16717 22969
rect 16787 22909 16821 22943
rect 16872 22923 16906 22957
rect 16983 22923 17017 22957
rect 17182 22917 17216 22951
rect 17301 22923 17335 22957
rect 17404 22923 17438 22957
rect 17602 22923 17636 22957
rect 17708 22978 17742 23012
rect 17708 22910 17742 22944
rect 17792 22939 17826 22973
rect 17876 22980 17910 23014
rect 17876 22912 17910 22946
rect 17980 22935 18014 22969
rect 18075 22909 18109 22943
rect 18159 22947 18193 22981
rect 15649 17549 15683 17583
rect 15649 17481 15683 17515
rect 15733 17549 15767 17583
rect 16427 17587 16461 17621
rect 16427 17519 16461 17553
rect 15733 17481 15767 17515
rect 16511 17587 16545 17621
rect 16511 17519 16545 17553
rect 17301 17589 17335 17623
rect 17301 17521 17335 17555
rect 17385 17589 17419 17623
rect 17385 17521 17419 17555
rect 18069 17579 18103 17613
rect 18069 17511 18103 17545
rect 18153 17579 18187 17613
rect 18153 17511 18187 17545
rect 19191 17581 19225 17615
rect 19191 17513 19225 17547
rect 19275 17581 19309 17615
rect 19275 17513 19309 17547
rect 20065 17583 20099 17617
rect 20065 17515 20099 17549
rect 20149 17583 20183 17617
rect 20149 17515 20183 17549
rect 20833 17573 20867 17607
rect 20833 17505 20867 17539
rect 20917 17573 20951 17607
rect 20917 17505 20951 17539
rect 21447 17571 21481 17605
rect 21447 17503 21481 17537
rect 21531 17571 21565 17605
rect 21531 17503 21565 17537
rect 22321 17573 22355 17607
rect 22321 17505 22355 17539
rect 22405 17573 22439 17607
rect 22405 17505 22439 17539
rect 23089 17563 23123 17597
rect 23089 17495 23123 17529
rect 23173 17563 23207 17597
rect 23173 17495 23207 17529
rect 9377 16107 9411 16141
rect 9461 16129 9495 16163
rect 9545 16107 9579 16141
rect 9713 16109 9747 16143
rect 9813 16109 9847 16143
rect 9903 16180 9937 16214
rect 9903 16112 9937 16146
rect 9503 15389 9537 15423
rect 9695 15361 9729 15395
rect 9779 15361 9813 15395
rect 11509 15259 11543 15293
rect 11950 15319 11984 15353
rect 11950 15251 11984 15285
rect 12049 15319 12083 15353
rect 12049 15251 12083 15285
rect 10687 14779 10721 14813
rect 10879 14751 10913 14785
rect 10963 14751 10997 14785
rect 9387 14543 9421 14577
rect 9471 14565 9505 14599
rect 9555 14543 9589 14577
rect 9723 14545 9757 14579
rect 9823 14545 9857 14579
rect 9913 14616 9947 14650
rect 9913 14548 9947 14582
rect 9513 13825 9547 13859
rect 9705 13797 9739 13831
rect 9789 13797 9823 13831
rect 10725 13793 10759 13827
rect 11166 13853 11200 13887
rect 11166 13785 11200 13819
rect 11265 13853 11299 13887
rect 11265 13785 11299 13819
rect 12623 13793 12657 13827
rect 12713 13787 12747 13821
rect 12803 13773 12837 13807
rect 12887 13787 12921 13821
rect 12981 13773 13015 13807
rect 13069 13811 13103 13845
rect 11724 13421 11758 13455
rect 11808 13421 11842 13455
rect 11904 13421 11938 13455
rect 11989 13481 12023 13515
rect 11989 13413 12023 13447
rect 9379 12875 9413 12909
rect 9463 12897 9497 12931
rect 9547 12875 9581 12909
rect 9715 12877 9749 12911
rect 9815 12877 9849 12911
rect 9905 12948 9939 12982
rect 10849 12943 10883 12977
rect 11121 12959 11155 12993
rect 11205 12969 11239 13003
rect 9905 12880 9939 12914
rect 9505 12157 9539 12191
rect 9697 12129 9731 12163
rect 9781 12129 9815 12163
rect 10881 11951 10915 11985
rect 11073 11923 11107 11957
rect 11157 11923 11191 11957
rect 9389 11311 9423 11345
rect 9473 11333 9507 11367
rect 9557 11311 9591 11345
rect 9725 11313 9759 11347
rect 9825 11313 9859 11347
rect 9915 11384 9949 11418
rect 9915 11316 9949 11350
rect 9515 10593 9549 10627
rect 9707 10565 9741 10599
rect 9791 10565 9825 10599
rect 6194 6503 6228 6537
rect 6194 6435 6228 6469
rect 6278 6503 6312 6537
rect 6278 6435 6312 6469
rect 10088 5839 10122 5873
rect 10187 5879 10221 5913
rect 10439 5867 10473 5901
rect 10540 5862 10574 5896
rect 10624 5879 10658 5913
rect 10708 5862 10742 5896
rect 10792 5870 10826 5904
rect 10896 5862 10930 5896
rect 10980 5879 11014 5913
rect 11064 5862 11098 5896
rect 11148 5862 11182 5896
rect 11337 5875 11371 5909
rect 1906 5419 1940 5453
rect 2005 5459 2039 5493
rect 2257 5447 2291 5481
rect 2358 5442 2392 5476
rect 2442 5459 2476 5493
rect 2526 5442 2560 5476
rect 2610 5450 2644 5484
rect 2714 5442 2748 5476
rect 2798 5459 2832 5493
rect 2882 5442 2916 5476
rect 2966 5442 3000 5476
rect 3155 5455 3189 5489
rect 3239 5419 3273 5453
rect 4040 5411 4074 5445
rect 4139 5451 4173 5485
rect 4391 5439 4425 5473
rect 4492 5434 4526 5468
rect 4576 5451 4610 5485
rect 4660 5434 4694 5468
rect 4744 5442 4778 5476
rect 4848 5434 4882 5468
rect 4932 5451 4966 5485
rect 5016 5434 5050 5468
rect 5100 5434 5134 5468
rect 5289 5447 5323 5481
rect 5373 5411 5407 5445
rect 5992 5411 6026 5445
rect 6091 5451 6125 5485
rect 6343 5439 6377 5473
rect 6444 5434 6478 5468
rect 6528 5451 6562 5485
rect 6612 5434 6646 5468
rect 6696 5442 6730 5476
rect 6800 5434 6834 5468
rect 6884 5451 6918 5485
rect 6968 5434 7002 5468
rect 7052 5434 7086 5468
rect 7241 5447 7275 5481
rect 7325 5411 7359 5445
rect 7994 5417 8028 5451
rect 8093 5457 8127 5491
rect 8345 5445 8379 5479
rect 8446 5440 8480 5474
rect 8530 5457 8564 5491
rect 8614 5440 8648 5474
rect 8698 5448 8732 5482
rect 8802 5440 8836 5474
rect 8886 5457 8920 5491
rect 8970 5440 9004 5474
rect 9054 5440 9088 5474
rect 9243 5453 9277 5487
rect 11421 5839 11455 5873
rect 12150 5827 12184 5861
rect 12249 5867 12283 5901
rect 12501 5855 12535 5889
rect 12602 5850 12636 5884
rect 12686 5867 12720 5901
rect 12770 5850 12804 5884
rect 12854 5858 12888 5892
rect 12958 5850 12992 5884
rect 13042 5867 13076 5901
rect 13126 5850 13160 5884
rect 13210 5850 13244 5884
rect 13399 5863 13433 5897
rect 9327 5417 9361 5451
rect 13483 5827 13517 5861
rect 14108 5835 14142 5869
rect 14207 5875 14241 5909
rect 14459 5863 14493 5897
rect 14560 5858 14594 5892
rect 14644 5875 14678 5909
rect 14728 5858 14762 5892
rect 14812 5866 14846 5900
rect 14916 5858 14950 5892
rect 15000 5875 15034 5909
rect 15084 5858 15118 5892
rect 15168 5858 15202 5892
rect 15357 5871 15391 5905
rect 15441 5835 15475 5869
rect 16102 5841 16136 5875
rect 16201 5881 16235 5915
rect 16453 5869 16487 5903
rect 16554 5864 16588 5898
rect 16638 5881 16672 5915
rect 16722 5864 16756 5898
rect 16806 5872 16840 5906
rect 16910 5864 16944 5898
rect 16994 5881 17028 5915
rect 17078 5864 17112 5898
rect 17162 5864 17196 5898
rect 17351 5877 17385 5911
rect 17435 5841 17469 5875
rect 10116 4965 10150 4999
rect 10215 5005 10249 5039
rect 10467 4993 10501 5027
rect 10568 4988 10602 5022
rect 10652 5005 10686 5039
rect 10736 4988 10770 5022
rect 10820 4996 10854 5030
rect 10924 4988 10958 5022
rect 11008 5005 11042 5039
rect 11092 4988 11126 5022
rect 11176 4988 11210 5022
rect 11365 5001 11399 5035
rect 11449 4965 11483 4999
rect 12386 4921 12420 4955
rect 12485 4961 12519 4995
rect 12737 4949 12771 4983
rect 12838 4944 12872 4978
rect 12922 4961 12956 4995
rect 13006 4944 13040 4978
rect 13090 4952 13124 4986
rect 13194 4944 13228 4978
rect 13278 4961 13312 4995
rect 13362 4944 13396 4978
rect 13446 4944 13480 4978
rect 13635 4957 13669 4991
rect 13719 4921 13753 4955
rect 14388 4915 14422 4949
rect 14487 4955 14521 4989
rect 14739 4943 14773 4977
rect 14840 4938 14874 4972
rect 14924 4955 14958 4989
rect 15008 4938 15042 4972
rect 15092 4946 15126 4980
rect 15196 4938 15230 4972
rect 15280 4955 15314 4989
rect 15364 4938 15398 4972
rect 15448 4938 15482 4972
rect 15637 4951 15671 4985
rect 15721 4915 15755 4949
rect 16410 4897 16444 4931
rect 16509 4937 16543 4971
rect 16761 4925 16795 4959
rect 16862 4920 16896 4954
rect 16946 4937 16980 4971
rect 17030 4920 17064 4954
rect 17114 4928 17148 4962
rect 17218 4920 17252 4954
rect 17302 4937 17336 4971
rect 17386 4920 17420 4954
rect 17470 4920 17504 4954
rect 17659 4933 17693 4967
rect 17743 4897 17777 4931
rect 1876 2159 1910 2193
rect 1975 2199 2009 2233
rect 2227 2187 2261 2221
rect 2328 2182 2362 2216
rect 2412 2199 2446 2233
rect 2496 2182 2530 2216
rect 2580 2190 2614 2224
rect 2684 2182 2718 2216
rect 2768 2199 2802 2233
rect 2852 2182 2886 2216
rect 2936 2182 2970 2216
rect 3125 2195 3159 2229
rect 3209 2159 3243 2193
rect 3946 2155 3980 2189
rect 4045 2195 4079 2229
rect 4297 2183 4331 2217
rect 4398 2178 4432 2212
rect 4482 2195 4516 2229
rect 4566 2178 4600 2212
rect 4650 2186 4684 2220
rect 4754 2178 4788 2212
rect 4838 2195 4872 2229
rect 4922 2178 4956 2212
rect 5006 2178 5040 2212
rect 5195 2191 5229 2225
rect 5279 2155 5313 2189
rect 5898 2155 5932 2189
rect 5997 2195 6031 2229
rect 6249 2183 6283 2217
rect 6350 2178 6384 2212
rect 6434 2195 6468 2229
rect 6518 2178 6552 2212
rect 6602 2186 6636 2220
rect 6706 2178 6740 2212
rect 6790 2195 6824 2229
rect 6874 2178 6908 2212
rect 6958 2178 6992 2212
rect 7147 2191 7181 2225
rect 7231 2155 7265 2189
rect 7900 2161 7934 2195
rect 7999 2201 8033 2235
rect 8251 2189 8285 2223
rect 8352 2184 8386 2218
rect 8436 2201 8470 2235
rect 8520 2184 8554 2218
rect 8604 2192 8638 2226
rect 8708 2184 8742 2218
rect 8792 2201 8826 2235
rect 8876 2184 8910 2218
rect 8960 2184 8994 2218
rect 9149 2197 9183 2231
rect 9233 2161 9267 2195
rect 9852 2161 9886 2195
rect 9951 2201 9985 2235
rect 10203 2189 10237 2223
rect 10304 2184 10338 2218
rect 10388 2201 10422 2235
rect 10472 2184 10506 2218
rect 10556 2192 10590 2226
rect 10660 2184 10694 2218
rect 10744 2201 10778 2235
rect 10828 2184 10862 2218
rect 10912 2184 10946 2218
rect 11101 2197 11135 2231
rect 11185 2161 11219 2195
rect 11844 2161 11878 2195
rect 11943 2201 11977 2235
rect 12195 2189 12229 2223
rect 12296 2184 12330 2218
rect 12380 2201 12414 2235
rect 12464 2184 12498 2218
rect 12548 2192 12582 2226
rect 12652 2184 12686 2218
rect 12736 2201 12770 2235
rect 12820 2184 12854 2218
rect 12904 2184 12938 2218
rect 13093 2197 13127 2231
rect 13177 2161 13211 2195
rect 13796 2161 13830 2195
rect 13895 2201 13929 2235
rect 14147 2189 14181 2223
rect 14248 2184 14282 2218
rect 14332 2201 14366 2235
rect 14416 2184 14450 2218
rect 14500 2192 14534 2226
rect 14604 2184 14638 2218
rect 14688 2201 14722 2235
rect 14772 2184 14806 2218
rect 14856 2184 14890 2218
rect 15045 2197 15079 2231
rect 15129 2161 15163 2195
rect 15860 2161 15894 2195
rect 15959 2201 15993 2235
rect 16211 2189 16245 2223
rect 16312 2184 16346 2218
rect 16396 2201 16430 2235
rect 16480 2184 16514 2218
rect 16564 2192 16598 2226
rect 16668 2184 16702 2218
rect 16752 2201 16786 2235
rect 16836 2184 16870 2218
rect 16920 2184 16954 2218
rect 17109 2197 17143 2231
rect 17193 2161 17227 2195
<< pdiffc >>
rect 18525 35065 18559 35099
rect 18596 35065 18630 35099
rect 18667 35065 18701 35099
rect 18525 34981 18559 35015
rect 18593 34981 18627 35015
rect 18661 34981 18695 35015
rect 18525 34884 18559 34918
rect 18593 34884 18627 34918
rect 18531 34780 18565 34814
rect 18599 34780 18633 34814
rect 18667 34780 18701 34814
rect 18555 34696 18589 34730
rect 18635 34696 18669 34730
rect 18525 34610 18559 34644
rect 18596 34610 18630 34644
rect 18667 34610 18701 34644
rect 18533 34486 18567 34520
rect 18543 34287 18577 34321
rect 18533 34192 18567 34226
rect 18525 34108 18559 34142
rect 18593 34108 18627 34142
rect 18538 33869 18572 33903
rect 18533 33777 18567 33811
rect 18525 33693 18559 33727
rect 18533 33589 18567 33623
rect 18601 33589 18635 33623
rect 18549 33505 18583 33539
rect 18533 33421 18567 33455
rect 18601 33421 18635 33455
rect 18533 32759 18567 32793
rect 18604 32759 18638 32793
rect 18675 32759 18709 32793
rect 18533 32675 18567 32709
rect 18601 32675 18635 32709
rect 18669 32675 18703 32709
rect 18533 32578 18567 32612
rect 18601 32578 18635 32612
rect 18539 32474 18573 32508
rect 18607 32474 18641 32508
rect 18675 32474 18709 32508
rect 18563 32390 18597 32424
rect 18643 32390 18677 32424
rect 18533 32304 18567 32338
rect 18604 32304 18638 32338
rect 18675 32304 18709 32338
rect 18541 32180 18575 32214
rect 18551 31981 18585 32015
rect 18541 31886 18575 31920
rect 18533 31802 18567 31836
rect 18601 31802 18635 31836
rect 18546 31563 18580 31597
rect 18541 31471 18575 31505
rect 18533 31387 18567 31421
rect 18541 31283 18575 31317
rect 18609 31283 18643 31317
rect 18557 31199 18591 31233
rect 18541 31115 18575 31149
rect 18609 31115 18643 31149
rect 18541 30545 18575 30579
rect 18612 30545 18646 30579
rect 18683 30545 18717 30579
rect 18541 30461 18575 30495
rect 18609 30461 18643 30495
rect 18677 30461 18711 30495
rect 18541 30364 18575 30398
rect 18609 30364 18643 30398
rect 18547 30260 18581 30294
rect 18615 30260 18649 30294
rect 18683 30260 18717 30294
rect 18571 30176 18605 30210
rect 18651 30176 18685 30210
rect 18541 30090 18575 30124
rect 18612 30090 18646 30124
rect 18683 30090 18717 30124
rect 18549 29966 18583 30000
rect 18559 29767 18593 29801
rect 18549 29672 18583 29706
rect 18541 29588 18575 29622
rect 18609 29588 18643 29622
rect 18554 29349 18588 29383
rect 18549 29257 18583 29291
rect 18541 29173 18575 29207
rect 18549 29069 18583 29103
rect 18617 29069 18651 29103
rect 18565 28985 18599 29019
rect 18549 28901 18583 28935
rect 18617 28901 18651 28935
rect 18523 28345 18557 28379
rect 18594 28345 18628 28379
rect 18665 28345 18699 28379
rect 18523 28261 18557 28295
rect 18591 28261 18625 28295
rect 18659 28261 18693 28295
rect 18523 28164 18557 28198
rect 18591 28164 18625 28198
rect 18529 28060 18563 28094
rect 18597 28060 18631 28094
rect 18665 28060 18699 28094
rect 18553 27976 18587 28010
rect 18633 27976 18667 28010
rect 18523 27890 18557 27924
rect 18594 27890 18628 27924
rect 18665 27890 18699 27924
rect 18531 27766 18565 27800
rect 18541 27567 18575 27601
rect 18531 27472 18565 27506
rect 18523 27388 18557 27422
rect 18591 27388 18625 27422
rect 18536 27149 18570 27183
rect 18531 27057 18565 27091
rect 18523 26973 18557 27007
rect 18531 26869 18565 26903
rect 18599 26869 18633 26903
rect 18547 26785 18581 26819
rect 18531 26701 18565 26735
rect 18599 26701 18633 26735
rect 18531 26131 18565 26165
rect 18602 26131 18636 26165
rect 18673 26131 18707 26165
rect 18531 26047 18565 26081
rect 18599 26047 18633 26081
rect 18667 26047 18701 26081
rect 18531 25950 18565 25984
rect 18599 25950 18633 25984
rect 18537 25846 18571 25880
rect 18605 25846 18639 25880
rect 18673 25846 18707 25880
rect 18561 25762 18595 25796
rect 18641 25762 18675 25796
rect 18531 25676 18565 25710
rect 18602 25676 18636 25710
rect 18673 25676 18707 25710
rect 18539 25552 18573 25586
rect 18549 25353 18583 25387
rect 18539 25258 18573 25292
rect 18531 25174 18565 25208
rect 18599 25174 18633 25208
rect 18544 24935 18578 24969
rect 18539 24843 18573 24877
rect 18531 24759 18565 24793
rect 18539 24655 18573 24689
rect 18607 24655 18641 24689
rect 18555 24571 18589 24605
rect 18539 24487 18573 24521
rect 18607 24487 18641 24521
rect 7581 23287 7615 23321
rect 7581 23219 7615 23253
rect 7665 23271 7699 23305
rect 7749 23287 7783 23321
rect 7853 23295 7887 23329
rect 7937 23287 7971 23321
rect 8029 23282 8063 23316
rect 8268 23295 8302 23329
rect 7749 23219 7783 23253
rect 8268 23227 8302 23261
rect 8352 23287 8386 23321
rect 8447 23277 8481 23311
rect 8646 23287 8680 23321
rect 8770 23295 8804 23329
rect 8770 23224 8804 23258
rect 8770 23153 8804 23187
rect 8856 23265 8890 23299
rect 8856 23185 8890 23219
rect 8940 23289 8974 23323
rect 8940 23221 8974 23255
rect 9044 23295 9078 23329
rect 9044 23227 9078 23261
rect 9141 23295 9175 23329
rect 9141 23227 9175 23261
rect 8940 23153 8974 23187
rect 9141 23159 9175 23193
rect 9225 23295 9259 23329
rect 9225 23224 9259 23258
rect 9225 23153 9259 23187
rect 9795 23295 9829 23329
rect 9795 23227 9829 23261
rect 9879 23279 9913 23313
rect 9963 23295 9997 23329
rect 10067 23303 10101 23337
rect 10151 23295 10185 23329
rect 10243 23290 10277 23324
rect 10482 23303 10516 23337
rect 9963 23227 9997 23261
rect 10482 23235 10516 23269
rect 10566 23295 10600 23329
rect 10661 23285 10695 23319
rect 10860 23295 10894 23329
rect 10984 23303 11018 23337
rect 10984 23232 11018 23266
rect 10984 23161 11018 23195
rect 11070 23273 11104 23307
rect 11070 23193 11104 23227
rect 11154 23297 11188 23331
rect 11154 23229 11188 23263
rect 11258 23303 11292 23337
rect 11258 23235 11292 23269
rect 11355 23303 11389 23337
rect 11355 23235 11389 23269
rect 11154 23161 11188 23195
rect 11355 23167 11389 23201
rect 11439 23303 11473 23337
rect 11439 23232 11473 23266
rect 11439 23161 11473 23195
rect 11995 23277 12029 23311
rect 11995 23209 12029 23243
rect 12079 23261 12113 23295
rect 12163 23277 12197 23311
rect 12267 23285 12301 23319
rect 12351 23277 12385 23311
rect 12443 23272 12477 23306
rect 12682 23285 12716 23319
rect 12163 23209 12197 23243
rect 12682 23217 12716 23251
rect 12766 23277 12800 23311
rect 12861 23267 12895 23301
rect 13060 23277 13094 23311
rect 13184 23285 13218 23319
rect 13184 23214 13218 23248
rect 13184 23143 13218 23177
rect 13270 23255 13304 23289
rect 13270 23175 13304 23209
rect 13354 23279 13388 23313
rect 13354 23211 13388 23245
rect 13458 23285 13492 23319
rect 13458 23217 13492 23251
rect 13555 23285 13589 23319
rect 13555 23217 13589 23251
rect 13354 23143 13388 23177
rect 13555 23149 13589 23183
rect 13639 23285 13673 23319
rect 13639 23214 13673 23248
rect 13639 23143 13673 23177
rect 14209 23285 14243 23319
rect 14209 23217 14243 23251
rect 14293 23269 14327 23303
rect 14377 23285 14411 23319
rect 14481 23293 14515 23327
rect 14565 23285 14599 23319
rect 14657 23280 14691 23314
rect 14896 23293 14930 23327
rect 14377 23217 14411 23251
rect 14896 23225 14930 23259
rect 14980 23285 15014 23319
rect 15075 23275 15109 23309
rect 15274 23285 15308 23319
rect 15398 23293 15432 23327
rect 15398 23222 15432 23256
rect 15398 23151 15432 23185
rect 15484 23263 15518 23297
rect 15484 23183 15518 23217
rect 15568 23287 15602 23321
rect 15568 23219 15602 23253
rect 15672 23293 15706 23327
rect 15672 23225 15706 23259
rect 15769 23293 15803 23327
rect 15769 23225 15803 23259
rect 15568 23151 15602 23185
rect 15769 23157 15803 23191
rect 15853 23293 15887 23327
rect 15853 23222 15887 23256
rect 15853 23151 15887 23185
rect 16515 23293 16549 23327
rect 16515 23225 16549 23259
rect 16599 23277 16633 23311
rect 16683 23293 16717 23327
rect 16787 23301 16821 23335
rect 16871 23293 16905 23327
rect 16963 23288 16997 23322
rect 17202 23301 17236 23335
rect 16683 23225 16717 23259
rect 17202 23233 17236 23267
rect 17286 23293 17320 23327
rect 17381 23283 17415 23317
rect 17580 23293 17614 23327
rect 17704 23301 17738 23335
rect 17704 23230 17738 23264
rect 17704 23159 17738 23193
rect 17790 23271 17824 23305
rect 17790 23191 17824 23225
rect 17874 23295 17908 23329
rect 17874 23227 17908 23261
rect 17978 23301 18012 23335
rect 17978 23233 18012 23267
rect 18075 23301 18109 23335
rect 18075 23233 18109 23267
rect 17874 23159 17908 23193
rect 18075 23165 18109 23199
rect 18159 23301 18193 23335
rect 18159 23230 18193 23264
rect 18159 23159 18193 23193
rect 15649 17297 15683 17331
rect 15649 17229 15683 17263
rect 15649 17161 15683 17195
rect 15733 17297 15767 17331
rect 15733 17229 15767 17263
rect 16427 17335 16461 17369
rect 16427 17267 16461 17301
rect 15733 17161 15767 17195
rect 16427 17199 16461 17233
rect 16511 17335 16545 17369
rect 16511 17267 16545 17301
rect 16511 17199 16545 17233
rect 17301 17337 17335 17371
rect 17301 17269 17335 17303
rect 17301 17201 17335 17235
rect 17385 17337 17419 17371
rect 17385 17269 17419 17303
rect 17385 17201 17419 17235
rect 18069 17327 18103 17361
rect 18069 17259 18103 17293
rect 18069 17191 18103 17225
rect 18153 17327 18187 17361
rect 18153 17259 18187 17293
rect 18153 17191 18187 17225
rect 19191 17329 19225 17363
rect 19191 17261 19225 17295
rect 19191 17193 19225 17227
rect 19275 17329 19309 17363
rect 19275 17261 19309 17295
rect 19275 17193 19309 17227
rect 20065 17331 20099 17365
rect 20065 17263 20099 17297
rect 20065 17195 20099 17229
rect 20149 17331 20183 17365
rect 20149 17263 20183 17297
rect 20149 17195 20183 17229
rect 20833 17321 20867 17355
rect 20833 17253 20867 17287
rect 20833 17185 20867 17219
rect 20917 17321 20951 17355
rect 20917 17253 20951 17287
rect 20917 17185 20951 17219
rect 21447 17319 21481 17353
rect 21447 17251 21481 17285
rect 21447 17183 21481 17217
rect 21531 17319 21565 17353
rect 21531 17251 21565 17285
rect 21531 17183 21565 17217
rect 22321 17321 22355 17355
rect 22321 17253 22355 17287
rect 22321 17185 22355 17219
rect 22405 17321 22439 17355
rect 22405 17253 22439 17287
rect 22405 17185 22439 17219
rect 23089 17311 23123 17345
rect 23089 17243 23123 17277
rect 23089 17175 23123 17209
rect 23173 17311 23207 17345
rect 23173 17243 23207 17277
rect 23173 17175 23207 17209
rect 9377 16497 9411 16531
rect 9377 16429 9411 16463
rect 9545 16487 9579 16521
rect 9545 16419 9579 16453
rect 9629 16487 9663 16521
rect 9629 16419 9663 16453
rect 9713 16487 9747 16521
rect 9817 16487 9851 16521
rect 9817 16419 9851 16453
rect 9901 16489 9935 16523
rect 9901 16421 9935 16455
rect 9901 16353 9935 16387
rect 9503 15711 9537 15745
rect 9587 15711 9621 15745
rect 9695 15753 9729 15787
rect 9695 15685 9729 15719
rect 9799 15753 9833 15787
rect 9799 15685 9833 15719
rect 11509 15643 11543 15677
rect 11601 15635 11635 15669
rect 11703 15643 11737 15677
rect 11798 15635 11832 15669
rect 11949 15643 11983 15677
rect 11949 15575 11983 15609
rect 12049 15643 12083 15677
rect 12049 15575 12083 15609
rect 12049 15507 12083 15541
rect 10687 15101 10721 15135
rect 10771 15101 10805 15135
rect 10879 15143 10913 15177
rect 10879 15075 10913 15109
rect 9387 14933 9421 14967
rect 9387 14865 9421 14899
rect 9555 14923 9589 14957
rect 9555 14855 9589 14889
rect 9639 14923 9673 14957
rect 9639 14855 9673 14889
rect 9723 14923 9757 14957
rect 9827 14923 9861 14957
rect 9827 14855 9861 14889
rect 9911 14925 9945 14959
rect 9911 14857 9945 14891
rect 10983 15143 11017 15177
rect 10983 15075 11017 15109
rect 9911 14789 9945 14823
rect 9513 14147 9547 14181
rect 9597 14147 9631 14181
rect 9705 14189 9739 14223
rect 9705 14121 9739 14155
rect 9809 14189 9843 14223
rect 9809 14121 9843 14155
rect 10725 14177 10759 14211
rect 10817 14169 10851 14203
rect 10919 14177 10953 14211
rect 11014 14169 11048 14203
rect 11165 14177 11199 14211
rect 11165 14109 11199 14143
rect 11265 14177 11299 14211
rect 11265 14109 11299 14143
rect 12984 14161 13018 14195
rect 12984 14093 13018 14127
rect 11265 14041 11299 14075
rect 12623 14030 12657 14064
rect 13069 14130 13103 14164
rect 13069 14062 13103 14096
rect 11905 13787 11939 13821
rect 11736 13667 11770 13701
rect 11905 13719 11939 13753
rect 12005 13803 12039 13837
rect 12005 13735 12039 13769
rect 9379 13265 9413 13299
rect 9379 13197 9413 13231
rect 9547 13255 9581 13289
rect 9547 13187 9581 13221
rect 9631 13255 9665 13289
rect 9631 13187 9665 13221
rect 9715 13255 9749 13289
rect 9819 13255 9853 13289
rect 9819 13187 9853 13221
rect 11121 13335 11155 13369
rect 9903 13257 9937 13291
rect 9903 13189 9937 13223
rect 10849 13196 10883 13230
rect 10933 13226 10967 13260
rect 11026 13207 11060 13241
rect 9903 13121 9937 13155
rect 11205 13321 11239 13355
rect 11205 13253 11239 13287
rect 9505 12479 9539 12513
rect 9589 12479 9623 12513
rect 9697 12521 9731 12555
rect 9697 12453 9731 12487
rect 9801 12521 9835 12555
rect 9801 12453 9835 12487
rect 10881 12273 10915 12307
rect 10965 12273 10999 12307
rect 11073 12315 11107 12349
rect 11073 12247 11107 12281
rect 11177 12315 11211 12349
rect 11177 12247 11211 12281
rect 9389 11701 9423 11735
rect 9389 11633 9423 11667
rect 9557 11691 9591 11725
rect 9557 11623 9591 11657
rect 9641 11691 9675 11725
rect 9641 11623 9675 11657
rect 9725 11691 9759 11725
rect 9829 11691 9863 11725
rect 9829 11623 9863 11657
rect 9913 11693 9947 11727
rect 9913 11625 9947 11659
rect 9913 11557 9947 11591
rect 9515 10915 9549 10949
rect 9599 10915 9633 10949
rect 9707 10957 9741 10991
rect 9707 10889 9741 10923
rect 9811 10957 9845 10991
rect 9811 10889 9845 10923
rect 6194 6251 6228 6285
rect 6194 6183 6228 6217
rect 6194 6115 6228 6149
rect 6278 6251 6312 6285
rect 6278 6183 6312 6217
rect 6278 6115 6312 6149
rect 10088 5599 10122 5633
rect 1906 5179 1940 5213
rect 1906 5089 1940 5123
rect 10088 5509 10122 5543
rect 1990 5059 2024 5093
rect 2257 5071 2291 5105
rect 2358 5076 2392 5110
rect 2442 5059 2476 5093
rect 2526 5076 2560 5110
rect 2610 5063 2644 5097
rect 2714 5076 2748 5110
rect 2798 5059 2832 5093
rect 2882 5076 2916 5110
rect 2966 5076 3000 5110
rect 3155 5067 3189 5101
rect 3239 5176 3273 5210
rect 3239 5082 3273 5116
rect 4040 5171 4074 5205
rect 4040 5081 4074 5115
rect 4124 5051 4158 5085
rect 4391 5063 4425 5097
rect 4492 5068 4526 5102
rect 4576 5051 4610 5085
rect 4660 5068 4694 5102
rect 4744 5055 4778 5089
rect 4848 5068 4882 5102
rect 4932 5051 4966 5085
rect 5016 5068 5050 5102
rect 5100 5068 5134 5102
rect 5289 5059 5323 5093
rect 5373 5168 5407 5202
rect 5373 5074 5407 5108
rect 5992 5171 6026 5205
rect 5992 5081 6026 5115
rect 6076 5051 6110 5085
rect 6343 5063 6377 5097
rect 6444 5068 6478 5102
rect 6528 5051 6562 5085
rect 6612 5068 6646 5102
rect 6696 5055 6730 5089
rect 6800 5068 6834 5102
rect 6884 5051 6918 5085
rect 6968 5068 7002 5102
rect 7052 5068 7086 5102
rect 7241 5059 7275 5093
rect 7325 5168 7359 5202
rect 7325 5074 7359 5108
rect 7994 5177 8028 5211
rect 7994 5087 8028 5121
rect 10172 5479 10206 5513
rect 10439 5491 10473 5525
rect 10540 5496 10574 5530
rect 10624 5479 10658 5513
rect 10708 5496 10742 5530
rect 10792 5483 10826 5517
rect 10896 5496 10930 5530
rect 10980 5479 11014 5513
rect 11064 5496 11098 5530
rect 11148 5496 11182 5530
rect 11337 5487 11371 5521
rect 11421 5596 11455 5630
rect 11421 5502 11455 5536
rect 12150 5587 12184 5621
rect 12150 5497 12184 5531
rect 12234 5467 12268 5501
rect 12501 5479 12535 5513
rect 12602 5484 12636 5518
rect 12686 5467 12720 5501
rect 12770 5484 12804 5518
rect 12854 5471 12888 5505
rect 12958 5484 12992 5518
rect 13042 5467 13076 5501
rect 13126 5484 13160 5518
rect 13210 5484 13244 5518
rect 13399 5475 13433 5509
rect 13483 5584 13517 5618
rect 13483 5490 13517 5524
rect 14108 5595 14142 5629
rect 14108 5505 14142 5539
rect 14192 5475 14226 5509
rect 14459 5487 14493 5521
rect 14560 5492 14594 5526
rect 14644 5475 14678 5509
rect 14728 5492 14762 5526
rect 14812 5479 14846 5513
rect 14916 5492 14950 5526
rect 15000 5475 15034 5509
rect 15084 5492 15118 5526
rect 15168 5492 15202 5526
rect 15357 5483 15391 5517
rect 15441 5592 15475 5626
rect 15441 5498 15475 5532
rect 16102 5601 16136 5635
rect 16102 5511 16136 5545
rect 16186 5481 16220 5515
rect 16453 5493 16487 5527
rect 16554 5498 16588 5532
rect 16638 5481 16672 5515
rect 16722 5498 16756 5532
rect 16806 5485 16840 5519
rect 16910 5498 16944 5532
rect 16994 5481 17028 5515
rect 17078 5498 17112 5532
rect 17162 5498 17196 5532
rect 17351 5489 17385 5523
rect 17435 5598 17469 5632
rect 17435 5504 17469 5538
rect 8078 5057 8112 5091
rect 8345 5069 8379 5103
rect 8446 5074 8480 5108
rect 8530 5057 8564 5091
rect 8614 5074 8648 5108
rect 8698 5061 8732 5095
rect 8802 5074 8836 5108
rect 8886 5057 8920 5091
rect 8970 5074 9004 5108
rect 9054 5074 9088 5108
rect 9243 5065 9277 5099
rect 9327 5174 9361 5208
rect 9327 5080 9361 5114
rect 10116 4725 10150 4759
rect 10116 4635 10150 4669
rect 10200 4605 10234 4639
rect 10467 4617 10501 4651
rect 10568 4622 10602 4656
rect 10652 4605 10686 4639
rect 10736 4622 10770 4656
rect 10820 4609 10854 4643
rect 10924 4622 10958 4656
rect 11008 4605 11042 4639
rect 11092 4622 11126 4656
rect 11176 4622 11210 4656
rect 11365 4613 11399 4647
rect 11449 4722 11483 4756
rect 11449 4628 11483 4662
rect 12386 4681 12420 4715
rect 12386 4591 12420 4625
rect 12470 4561 12504 4595
rect 12737 4573 12771 4607
rect 12838 4578 12872 4612
rect 12922 4561 12956 4595
rect 13006 4578 13040 4612
rect 13090 4565 13124 4599
rect 13194 4578 13228 4612
rect 13278 4561 13312 4595
rect 13362 4578 13396 4612
rect 13446 4578 13480 4612
rect 13635 4569 13669 4603
rect 13719 4678 13753 4712
rect 13719 4584 13753 4618
rect 14388 4675 14422 4709
rect 14388 4585 14422 4619
rect 14472 4555 14506 4589
rect 14739 4567 14773 4601
rect 14840 4572 14874 4606
rect 14924 4555 14958 4589
rect 15008 4572 15042 4606
rect 15092 4559 15126 4593
rect 15196 4572 15230 4606
rect 15280 4555 15314 4589
rect 15364 4572 15398 4606
rect 15448 4572 15482 4606
rect 15637 4563 15671 4597
rect 15721 4672 15755 4706
rect 15721 4578 15755 4612
rect 16410 4657 16444 4691
rect 16410 4567 16444 4601
rect 16494 4537 16528 4571
rect 16761 4549 16795 4583
rect 16862 4554 16896 4588
rect 16946 4537 16980 4571
rect 17030 4554 17064 4588
rect 17114 4541 17148 4575
rect 17218 4554 17252 4588
rect 17302 4537 17336 4571
rect 17386 4554 17420 4588
rect 17470 4554 17504 4588
rect 17659 4545 17693 4579
rect 17743 4654 17777 4688
rect 17743 4560 17777 4594
rect 1876 1919 1910 1953
rect 1876 1829 1910 1863
rect 1960 1799 1994 1833
rect 2227 1811 2261 1845
rect 2328 1816 2362 1850
rect 2412 1799 2446 1833
rect 2496 1816 2530 1850
rect 2580 1803 2614 1837
rect 2684 1816 2718 1850
rect 2768 1799 2802 1833
rect 2852 1816 2886 1850
rect 2936 1816 2970 1850
rect 3125 1807 3159 1841
rect 3209 1916 3243 1950
rect 3209 1822 3243 1856
rect 3946 1915 3980 1949
rect 3946 1825 3980 1859
rect 4030 1795 4064 1829
rect 4297 1807 4331 1841
rect 4398 1812 4432 1846
rect 4482 1795 4516 1829
rect 4566 1812 4600 1846
rect 4650 1799 4684 1833
rect 4754 1812 4788 1846
rect 4838 1795 4872 1829
rect 4922 1812 4956 1846
rect 5006 1812 5040 1846
rect 5195 1803 5229 1837
rect 5279 1912 5313 1946
rect 5279 1818 5313 1852
rect 5898 1915 5932 1949
rect 5898 1825 5932 1859
rect 5982 1795 6016 1829
rect 6249 1807 6283 1841
rect 6350 1812 6384 1846
rect 6434 1795 6468 1829
rect 6518 1812 6552 1846
rect 6602 1799 6636 1833
rect 6706 1812 6740 1846
rect 6790 1795 6824 1829
rect 6874 1812 6908 1846
rect 6958 1812 6992 1846
rect 7147 1803 7181 1837
rect 7231 1912 7265 1946
rect 7231 1818 7265 1852
rect 7900 1921 7934 1955
rect 7900 1831 7934 1865
rect 7984 1801 8018 1835
rect 8251 1813 8285 1847
rect 8352 1818 8386 1852
rect 8436 1801 8470 1835
rect 8520 1818 8554 1852
rect 8604 1805 8638 1839
rect 8708 1818 8742 1852
rect 8792 1801 8826 1835
rect 8876 1818 8910 1852
rect 8960 1818 8994 1852
rect 9149 1809 9183 1843
rect 9233 1918 9267 1952
rect 9233 1824 9267 1858
rect 9852 1921 9886 1955
rect 9852 1831 9886 1865
rect 9936 1801 9970 1835
rect 10203 1813 10237 1847
rect 10304 1818 10338 1852
rect 10388 1801 10422 1835
rect 10472 1818 10506 1852
rect 10556 1805 10590 1839
rect 10660 1818 10694 1852
rect 10744 1801 10778 1835
rect 10828 1818 10862 1852
rect 10912 1818 10946 1852
rect 11101 1809 11135 1843
rect 11185 1918 11219 1952
rect 11185 1824 11219 1858
rect 11844 1921 11878 1955
rect 11844 1831 11878 1865
rect 11928 1801 11962 1835
rect 12195 1813 12229 1847
rect 12296 1818 12330 1852
rect 12380 1801 12414 1835
rect 12464 1818 12498 1852
rect 12548 1805 12582 1839
rect 12652 1818 12686 1852
rect 12736 1801 12770 1835
rect 12820 1818 12854 1852
rect 12904 1818 12938 1852
rect 13093 1809 13127 1843
rect 13177 1918 13211 1952
rect 13177 1824 13211 1858
rect 13796 1921 13830 1955
rect 13796 1831 13830 1865
rect 13880 1801 13914 1835
rect 14147 1813 14181 1847
rect 14248 1818 14282 1852
rect 14332 1801 14366 1835
rect 14416 1818 14450 1852
rect 14500 1805 14534 1839
rect 14604 1818 14638 1852
rect 14688 1801 14722 1835
rect 14772 1818 14806 1852
rect 14856 1818 14890 1852
rect 15045 1809 15079 1843
rect 15129 1918 15163 1952
rect 15129 1824 15163 1858
rect 15860 1921 15894 1955
rect 15860 1831 15894 1865
rect 15944 1801 15978 1835
rect 16211 1813 16245 1847
rect 16312 1818 16346 1852
rect 16396 1801 16430 1835
rect 16480 1818 16514 1852
rect 16564 1805 16598 1839
rect 16668 1818 16702 1852
rect 16752 1801 16786 1835
rect 16836 1818 16870 1852
rect 16920 1818 16954 1852
rect 17109 1809 17143 1843
rect 17193 1918 17227 1952
rect 17193 1824 17227 1858
<< psubdiff >>
rect 18841 35163 18865 35197
rect 18899 35163 18946 35197
rect 18849 32857 18873 32891
rect 18907 32857 18954 32891
rect 18857 30643 18881 30677
rect 18915 30643 18962 30677
rect 18839 28443 18863 28477
rect 18897 28443 18944 28477
rect 18847 26229 18871 26263
rect 18905 26229 18952 26263
rect 9323 22989 9357 23013
rect 9323 22908 9357 22955
rect 11537 22997 11571 23021
rect 11537 22916 11571 22963
rect 13737 22979 13771 23003
rect 13737 22898 13771 22945
rect 15951 22987 15985 23011
rect 15951 22906 15985 22953
rect 18257 22995 18291 23019
rect 18257 22914 18291 22961
rect 15510 17535 15544 17582
rect 15510 17477 15544 17501
rect 16296 17573 16330 17620
rect 16296 17515 16330 17539
rect 17162 17575 17196 17622
rect 17162 17517 17196 17541
rect 17940 17565 17974 17612
rect 17940 17507 17974 17531
rect 19056 17567 19090 17614
rect 19056 17509 19090 17533
rect 19922 17569 19956 17616
rect 19922 17511 19956 17535
rect 20692 17559 20726 17606
rect 20692 17501 20726 17525
rect 21670 17557 21704 17604
rect 21670 17499 21704 17523
rect 22178 17559 22212 17606
rect 22178 17501 22212 17525
rect 23310 17549 23344 17596
rect 23310 17491 23344 17515
<< nsubdiff >>
rect 18530 35163 18554 35197
rect 18588 35163 18647 35197
rect 18681 35163 18705 35197
rect 18538 32857 18562 32891
rect 18596 32857 18655 32891
rect 18689 32857 18713 32891
rect 18546 30643 18570 30677
rect 18604 30643 18663 30677
rect 18697 30643 18721 30677
rect 18528 28443 18552 28477
rect 18586 28443 18645 28477
rect 18679 28443 18703 28477
rect 18536 26229 18560 26263
rect 18594 26229 18653 26263
rect 18687 26229 18711 26263
rect 9323 23300 9357 23324
rect 9323 23207 9357 23266
rect 9323 23149 9357 23173
rect 11537 23308 11571 23332
rect 11537 23215 11571 23274
rect 11537 23157 11571 23181
rect 13737 23290 13771 23314
rect 13737 23197 13771 23256
rect 13737 23139 13771 23163
rect 15951 23298 15985 23322
rect 15951 23205 15985 23264
rect 15951 23147 15985 23171
rect 18257 23306 18291 23330
rect 18257 23213 18291 23272
rect 18257 23155 18291 23179
rect 16296 17355 16330 17379
rect 15510 17317 15544 17341
rect 15510 17224 15544 17283
rect 15510 17166 15544 17190
rect 16296 17262 16330 17321
rect 16296 17204 16330 17228
rect 17162 17357 17196 17381
rect 17162 17264 17196 17323
rect 17162 17206 17196 17230
rect 17940 17347 17974 17371
rect 17940 17254 17974 17313
rect 17940 17196 17974 17220
rect 19056 17349 19090 17373
rect 19056 17256 19090 17315
rect 19056 17198 19090 17222
rect 19922 17351 19956 17375
rect 19922 17258 19956 17317
rect 19922 17200 19956 17224
rect 20692 17341 20726 17365
rect 20692 17248 20726 17307
rect 20692 17190 20726 17214
rect 21670 17339 21704 17363
rect 21670 17246 21704 17305
rect 21670 17188 21704 17212
rect 22178 17341 22212 17365
rect 22178 17248 22212 17307
rect 22178 17190 22212 17214
rect 23310 17331 23344 17355
rect 23310 17238 23344 17297
rect 23310 17180 23344 17204
<< psubdiffcont >>
rect 18865 35163 18899 35197
rect 18873 32857 18907 32891
rect 18881 30643 18915 30677
rect 18863 28443 18897 28477
rect 18871 26229 18905 26263
rect 9323 22955 9357 22989
rect 11537 22963 11571 22997
rect 13737 22945 13771 22979
rect 15951 22953 15985 22987
rect 18257 22961 18291 22995
rect 15510 17501 15544 17535
rect 16296 17539 16330 17573
rect 17162 17541 17196 17575
rect 17940 17531 17974 17565
rect 19056 17533 19090 17567
rect 19922 17535 19956 17569
rect 20692 17525 20726 17559
rect 21670 17523 21704 17557
rect 22178 17525 22212 17559
rect 23310 17515 23344 17549
<< nsubdiffcont >>
rect 18554 35163 18588 35197
rect 18647 35163 18681 35197
rect 18562 32857 18596 32891
rect 18655 32857 18689 32891
rect 18570 30643 18604 30677
rect 18663 30643 18697 30677
rect 18552 28443 18586 28477
rect 18645 28443 18679 28477
rect 18560 26229 18594 26263
rect 18653 26229 18687 26263
rect 9323 23266 9357 23300
rect 9323 23173 9357 23207
rect 11537 23274 11571 23308
rect 11537 23181 11571 23215
rect 13737 23256 13771 23290
rect 13737 23163 13771 23197
rect 15951 23264 15985 23298
rect 15951 23171 15985 23205
rect 18257 23272 18291 23306
rect 18257 23179 18291 23213
rect 15510 17283 15544 17317
rect 15510 17190 15544 17224
rect 16296 17321 16330 17355
rect 16296 17228 16330 17262
rect 17162 17323 17196 17357
rect 17162 17230 17196 17264
rect 17940 17313 17974 17347
rect 17940 17220 17974 17254
rect 19056 17315 19090 17349
rect 19056 17222 19090 17256
rect 19922 17317 19956 17351
rect 19922 17224 19956 17258
rect 20692 17307 20726 17341
rect 20692 17214 20726 17248
rect 21670 17305 21704 17339
rect 21670 17212 21704 17246
rect 22178 17307 22212 17341
rect 22178 17214 22212 17248
rect 23310 17297 23344 17331
rect 23310 17204 23344 17238
<< poly >>
rect 18487 35025 18513 35055
rect 18713 35035 18833 35055
rect 18713 35025 18761 35035
rect 18745 35001 18761 35025
rect 18795 35025 18833 35035
rect 18963 35025 18989 35055
rect 18795 35001 18811 35025
rect 18745 34991 18811 35001
rect 18487 34928 18513 34958
rect 18641 34949 18707 34958
rect 18840 34949 18879 34960
rect 18641 34930 18879 34949
rect 18963 34930 18989 34960
rect 18641 34928 18864 34930
rect 18677 34919 18864 34928
rect 18745 34774 18811 34919
rect 18745 34770 18761 34774
rect 18487 34740 18513 34770
rect 18713 34740 18761 34770
rect 18795 34772 18811 34774
rect 18795 34742 18833 34772
rect 18963 34742 18989 34772
rect 18795 34740 18811 34742
rect 18745 34730 18811 34740
rect 18745 34686 18833 34688
rect 18487 34656 18513 34686
rect 18713 34658 18833 34686
rect 18963 34658 18989 34688
rect 18713 34656 18811 34658
rect 18745 34590 18811 34656
rect 18745 34556 18761 34590
rect 18795 34556 18811 34590
rect 18745 34546 18811 34556
rect 18629 34516 18695 34526
rect 18629 34482 18645 34516
rect 18679 34498 18695 34516
rect 18679 34482 18879 34498
rect 18629 34475 18879 34482
rect 18487 34445 18513 34475
rect 18597 34468 18879 34475
rect 18963 34468 18989 34498
rect 18597 34445 18695 34468
rect 18635 34380 18689 34396
rect 18635 34361 18645 34380
rect 18487 34331 18513 34361
rect 18597 34346 18645 34361
rect 18679 34346 18689 34380
rect 18597 34331 18689 34346
rect 18635 34330 18689 34331
rect 18731 34373 18891 34403
rect 18963 34373 18989 34403
rect 18731 34288 18761 34373
rect 18695 34278 18761 34288
rect 18695 34277 18711 34278
rect 18487 34247 18513 34277
rect 18597 34247 18711 34277
rect 18695 34244 18711 34247
rect 18745 34244 18761 34278
rect 18803 34321 18869 34331
rect 18803 34287 18819 34321
rect 18853 34297 18869 34321
rect 18853 34287 18891 34297
rect 18803 34267 18891 34287
rect 18963 34267 18989 34297
rect 18695 34234 18761 34244
rect 18790 34182 18835 34196
rect 18487 34152 18513 34182
rect 18663 34166 18835 34182
rect 18963 34166 18989 34196
rect 18663 34152 18820 34166
rect 18701 34142 18755 34152
rect 18701 34108 18711 34142
rect 18745 34108 18755 34142
rect 18701 34092 18755 34108
rect 18797 34078 18851 34094
rect 18797 34050 18807 34078
rect 18487 34020 18513 34050
rect 18597 34044 18807 34050
rect 18841 34077 18851 34078
rect 18841 34047 18879 34077
rect 18963 34047 18989 34077
rect 18841 34044 18851 34047
rect 18597 34020 18851 34044
rect 18629 33968 18695 33978
rect 18629 33947 18645 33968
rect 18487 33917 18513 33947
rect 18597 33934 18645 33947
rect 18679 33934 18695 33968
rect 18597 33917 18695 33934
rect 18737 33948 18891 33978
rect 18963 33948 18989 33978
rect 18737 33875 18767 33948
rect 18713 33859 18767 33875
rect 18713 33852 18723 33859
rect 18487 33822 18513 33852
rect 18597 33825 18723 33852
rect 18757 33825 18767 33859
rect 18809 33879 18863 33895
rect 18809 33845 18819 33879
rect 18853 33849 18891 33879
rect 18963 33849 18989 33879
rect 18853 33845 18863 33849
rect 18809 33829 18863 33845
rect 18597 33822 18767 33825
rect 18713 33809 18767 33822
rect 18487 33737 18513 33767
rect 18597 33737 18879 33767
rect 18963 33737 18989 33767
rect 18677 33716 18743 33737
rect 18677 33682 18693 33716
rect 18727 33682 18743 33716
rect 18677 33672 18743 33682
rect 18493 33549 18519 33579
rect 18647 33554 18879 33579
rect 18647 33549 18746 33554
rect 18736 33520 18746 33549
rect 18780 33549 18879 33554
rect 18963 33549 18989 33579
rect 18780 33520 18790 33549
rect 18736 33504 18790 33520
rect 18493 33465 18519 33495
rect 18647 33465 18692 33495
rect 18662 33462 18692 33465
rect 18834 33465 18879 33495
rect 18963 33465 18989 33495
rect 18834 33462 18864 33465
rect 18662 33452 18864 33462
rect 18662 33432 18761 33452
rect 18745 33418 18761 33432
rect 18795 33432 18864 33452
rect 18795 33418 18811 33432
rect 18745 33408 18811 33418
rect 18495 32719 18521 32749
rect 18721 32729 18841 32749
rect 18721 32719 18769 32729
rect 18753 32695 18769 32719
rect 18803 32719 18841 32729
rect 18971 32719 18997 32749
rect 18803 32695 18819 32719
rect 18753 32685 18819 32695
rect 18495 32622 18521 32652
rect 18649 32643 18715 32652
rect 18848 32643 18887 32654
rect 18649 32624 18887 32643
rect 18971 32624 18997 32654
rect 18649 32622 18872 32624
rect 18685 32613 18872 32622
rect 18753 32468 18819 32613
rect 18753 32464 18769 32468
rect 18495 32434 18521 32464
rect 18721 32434 18769 32464
rect 18803 32466 18819 32468
rect 18803 32436 18841 32466
rect 18971 32436 18997 32466
rect 18803 32434 18819 32436
rect 18753 32424 18819 32434
rect 18753 32380 18841 32382
rect 18495 32350 18521 32380
rect 18721 32352 18841 32380
rect 18971 32352 18997 32382
rect 18721 32350 18819 32352
rect 18753 32284 18819 32350
rect 18753 32250 18769 32284
rect 18803 32250 18819 32284
rect 18753 32240 18819 32250
rect 18637 32210 18703 32220
rect 18637 32176 18653 32210
rect 18687 32192 18703 32210
rect 18687 32176 18887 32192
rect 18637 32169 18887 32176
rect 18495 32139 18521 32169
rect 18605 32162 18887 32169
rect 18971 32162 18997 32192
rect 18605 32139 18703 32162
rect 18643 32074 18697 32090
rect 18643 32055 18653 32074
rect 18495 32025 18521 32055
rect 18605 32040 18653 32055
rect 18687 32040 18697 32074
rect 18605 32025 18697 32040
rect 18643 32024 18697 32025
rect 18739 32067 18899 32097
rect 18971 32067 18997 32097
rect 18739 31982 18769 32067
rect 18703 31972 18769 31982
rect 18703 31971 18719 31972
rect 18495 31941 18521 31971
rect 18605 31941 18719 31971
rect 18703 31938 18719 31941
rect 18753 31938 18769 31972
rect 18811 32015 18877 32025
rect 18811 31981 18827 32015
rect 18861 31991 18877 32015
rect 18861 31981 18899 31991
rect 18811 31961 18899 31981
rect 18971 31961 18997 31991
rect 18703 31928 18769 31938
rect 18798 31876 18843 31890
rect 18495 31846 18521 31876
rect 18671 31860 18843 31876
rect 18971 31860 18997 31890
rect 18671 31846 18828 31860
rect 18709 31836 18763 31846
rect 18709 31802 18719 31836
rect 18753 31802 18763 31836
rect 18709 31786 18763 31802
rect 18805 31772 18859 31788
rect 18805 31744 18815 31772
rect 18495 31714 18521 31744
rect 18605 31738 18815 31744
rect 18849 31771 18859 31772
rect 18849 31741 18887 31771
rect 18971 31741 18997 31771
rect 18849 31738 18859 31741
rect 18605 31714 18859 31738
rect 18637 31662 18703 31672
rect 18637 31641 18653 31662
rect 18495 31611 18521 31641
rect 18605 31628 18653 31641
rect 18687 31628 18703 31662
rect 18605 31611 18703 31628
rect 18745 31642 18899 31672
rect 18971 31642 18997 31672
rect 18745 31569 18775 31642
rect 18721 31553 18775 31569
rect 18721 31546 18731 31553
rect 18495 31516 18521 31546
rect 18605 31519 18731 31546
rect 18765 31519 18775 31553
rect 18817 31573 18871 31589
rect 18817 31539 18827 31573
rect 18861 31543 18899 31573
rect 18971 31543 18997 31573
rect 18861 31539 18871 31543
rect 18817 31523 18871 31539
rect 18605 31516 18775 31519
rect 18721 31503 18775 31516
rect 18495 31431 18521 31461
rect 18605 31431 18887 31461
rect 18971 31431 18997 31461
rect 18685 31410 18751 31431
rect 18685 31376 18701 31410
rect 18735 31376 18751 31410
rect 18685 31366 18751 31376
rect 18501 31243 18527 31273
rect 18655 31248 18887 31273
rect 18655 31243 18754 31248
rect 18744 31214 18754 31243
rect 18788 31243 18887 31248
rect 18971 31243 18997 31273
rect 18788 31214 18798 31243
rect 18744 31198 18798 31214
rect 18501 31159 18527 31189
rect 18655 31159 18700 31189
rect 18670 31156 18700 31159
rect 18842 31159 18887 31189
rect 18971 31159 18997 31189
rect 18842 31156 18872 31159
rect 18670 31146 18872 31156
rect 18670 31126 18769 31146
rect 18753 31112 18769 31126
rect 18803 31126 18872 31146
rect 18803 31112 18819 31126
rect 18753 31102 18819 31112
rect 18503 30505 18529 30535
rect 18729 30515 18849 30535
rect 18729 30505 18777 30515
rect 18761 30481 18777 30505
rect 18811 30505 18849 30515
rect 18979 30505 19005 30535
rect 18811 30481 18827 30505
rect 18761 30471 18827 30481
rect 18503 30408 18529 30438
rect 18657 30429 18723 30438
rect 18856 30429 18895 30440
rect 18657 30410 18895 30429
rect 18979 30410 19005 30440
rect 18657 30408 18880 30410
rect 18693 30399 18880 30408
rect 18761 30254 18827 30399
rect 18761 30250 18777 30254
rect 18503 30220 18529 30250
rect 18729 30220 18777 30250
rect 18811 30252 18827 30254
rect 18811 30222 18849 30252
rect 18979 30222 19005 30252
rect 18811 30220 18827 30222
rect 18761 30210 18827 30220
rect 18761 30166 18849 30168
rect 18503 30136 18529 30166
rect 18729 30138 18849 30166
rect 18979 30138 19005 30168
rect 18729 30136 18827 30138
rect 18761 30070 18827 30136
rect 18761 30036 18777 30070
rect 18811 30036 18827 30070
rect 18761 30026 18827 30036
rect 18645 29996 18711 30006
rect 18645 29962 18661 29996
rect 18695 29978 18711 29996
rect 18695 29962 18895 29978
rect 18645 29955 18895 29962
rect 18503 29925 18529 29955
rect 18613 29948 18895 29955
rect 18979 29948 19005 29978
rect 18613 29925 18711 29948
rect 18651 29860 18705 29876
rect 18651 29841 18661 29860
rect 18503 29811 18529 29841
rect 18613 29826 18661 29841
rect 18695 29826 18705 29860
rect 18613 29811 18705 29826
rect 18651 29810 18705 29811
rect 18747 29853 18907 29883
rect 18979 29853 19005 29883
rect 18747 29768 18777 29853
rect 18711 29758 18777 29768
rect 18711 29757 18727 29758
rect 18503 29727 18529 29757
rect 18613 29727 18727 29757
rect 18711 29724 18727 29727
rect 18761 29724 18777 29758
rect 18819 29801 18885 29811
rect 18819 29767 18835 29801
rect 18869 29777 18885 29801
rect 18869 29767 18907 29777
rect 18819 29747 18907 29767
rect 18979 29747 19005 29777
rect 18711 29714 18777 29724
rect 18806 29662 18851 29676
rect 18503 29632 18529 29662
rect 18679 29646 18851 29662
rect 18979 29646 19005 29676
rect 18679 29632 18836 29646
rect 18717 29622 18771 29632
rect 18717 29588 18727 29622
rect 18761 29588 18771 29622
rect 18717 29572 18771 29588
rect 18813 29558 18867 29574
rect 18813 29530 18823 29558
rect 18503 29500 18529 29530
rect 18613 29524 18823 29530
rect 18857 29557 18867 29558
rect 18857 29527 18895 29557
rect 18979 29527 19005 29557
rect 18857 29524 18867 29527
rect 18613 29500 18867 29524
rect 18645 29448 18711 29458
rect 18645 29427 18661 29448
rect 18503 29397 18529 29427
rect 18613 29414 18661 29427
rect 18695 29414 18711 29448
rect 18613 29397 18711 29414
rect 18753 29428 18907 29458
rect 18979 29428 19005 29458
rect 18753 29355 18783 29428
rect 18729 29339 18783 29355
rect 18729 29332 18739 29339
rect 18503 29302 18529 29332
rect 18613 29305 18739 29332
rect 18773 29305 18783 29339
rect 18825 29359 18879 29375
rect 18825 29325 18835 29359
rect 18869 29329 18907 29359
rect 18979 29329 19005 29359
rect 18869 29325 18879 29329
rect 18825 29309 18879 29325
rect 18613 29302 18783 29305
rect 18729 29289 18783 29302
rect 18503 29217 18529 29247
rect 18613 29217 18895 29247
rect 18979 29217 19005 29247
rect 18693 29196 18759 29217
rect 18693 29162 18709 29196
rect 18743 29162 18759 29196
rect 18693 29152 18759 29162
rect 18509 29029 18535 29059
rect 18663 29034 18895 29059
rect 18663 29029 18762 29034
rect 18752 29000 18762 29029
rect 18796 29029 18895 29034
rect 18979 29029 19005 29059
rect 18796 29000 18806 29029
rect 18752 28984 18806 29000
rect 18509 28945 18535 28975
rect 18663 28945 18708 28975
rect 18678 28942 18708 28945
rect 18850 28945 18895 28975
rect 18979 28945 19005 28975
rect 18850 28942 18880 28945
rect 18678 28932 18880 28942
rect 18678 28912 18777 28932
rect 18761 28898 18777 28912
rect 18811 28912 18880 28932
rect 18811 28898 18827 28912
rect 18761 28888 18827 28898
rect 18485 28305 18511 28335
rect 18711 28315 18831 28335
rect 18711 28305 18759 28315
rect 18743 28281 18759 28305
rect 18793 28305 18831 28315
rect 18961 28305 18987 28335
rect 18793 28281 18809 28305
rect 18743 28271 18809 28281
rect 18485 28208 18511 28238
rect 18639 28229 18705 28238
rect 18838 28229 18877 28240
rect 18639 28210 18877 28229
rect 18961 28210 18987 28240
rect 18639 28208 18862 28210
rect 18675 28199 18862 28208
rect 18743 28054 18809 28199
rect 18743 28050 18759 28054
rect 18485 28020 18511 28050
rect 18711 28020 18759 28050
rect 18793 28052 18809 28054
rect 18793 28022 18831 28052
rect 18961 28022 18987 28052
rect 18793 28020 18809 28022
rect 18743 28010 18809 28020
rect 18743 27966 18831 27968
rect 18485 27936 18511 27966
rect 18711 27938 18831 27966
rect 18961 27938 18987 27968
rect 18711 27936 18809 27938
rect 18743 27870 18809 27936
rect 18743 27836 18759 27870
rect 18793 27836 18809 27870
rect 18743 27826 18809 27836
rect 18627 27796 18693 27806
rect 18627 27762 18643 27796
rect 18677 27778 18693 27796
rect 18677 27762 18877 27778
rect 18627 27755 18877 27762
rect 18485 27725 18511 27755
rect 18595 27748 18877 27755
rect 18961 27748 18987 27778
rect 18595 27725 18693 27748
rect 18633 27660 18687 27676
rect 18633 27641 18643 27660
rect 18485 27611 18511 27641
rect 18595 27626 18643 27641
rect 18677 27626 18687 27660
rect 18595 27611 18687 27626
rect 18633 27610 18687 27611
rect 18729 27653 18889 27683
rect 18961 27653 18987 27683
rect 18729 27568 18759 27653
rect 18693 27558 18759 27568
rect 18693 27557 18709 27558
rect 18485 27527 18511 27557
rect 18595 27527 18709 27557
rect 18693 27524 18709 27527
rect 18743 27524 18759 27558
rect 18801 27601 18867 27611
rect 18801 27567 18817 27601
rect 18851 27577 18867 27601
rect 18851 27567 18889 27577
rect 18801 27547 18889 27567
rect 18961 27547 18987 27577
rect 18693 27514 18759 27524
rect 18788 27462 18833 27476
rect 18485 27432 18511 27462
rect 18661 27446 18833 27462
rect 18961 27446 18987 27476
rect 18661 27432 18818 27446
rect 18699 27422 18753 27432
rect 18699 27388 18709 27422
rect 18743 27388 18753 27422
rect 18699 27372 18753 27388
rect 18795 27358 18849 27374
rect 18795 27330 18805 27358
rect 18485 27300 18511 27330
rect 18595 27324 18805 27330
rect 18839 27357 18849 27358
rect 18839 27327 18877 27357
rect 18961 27327 18987 27357
rect 18839 27324 18849 27327
rect 18595 27300 18849 27324
rect 18627 27248 18693 27258
rect 18627 27227 18643 27248
rect 18485 27197 18511 27227
rect 18595 27214 18643 27227
rect 18677 27214 18693 27248
rect 18595 27197 18693 27214
rect 18735 27228 18889 27258
rect 18961 27228 18987 27258
rect 18735 27155 18765 27228
rect 18711 27139 18765 27155
rect 18711 27132 18721 27139
rect 18485 27102 18511 27132
rect 18595 27105 18721 27132
rect 18755 27105 18765 27139
rect 18807 27159 18861 27175
rect 18807 27125 18817 27159
rect 18851 27129 18889 27159
rect 18961 27129 18987 27159
rect 18851 27125 18861 27129
rect 18807 27109 18861 27125
rect 18595 27102 18765 27105
rect 18711 27089 18765 27102
rect 18485 27017 18511 27047
rect 18595 27017 18877 27047
rect 18961 27017 18987 27047
rect 18675 26996 18741 27017
rect 18675 26962 18691 26996
rect 18725 26962 18741 26996
rect 18675 26952 18741 26962
rect 18491 26829 18517 26859
rect 18645 26834 18877 26859
rect 18645 26829 18744 26834
rect 18734 26800 18744 26829
rect 18778 26829 18877 26834
rect 18961 26829 18987 26859
rect 18778 26800 18788 26829
rect 18734 26784 18788 26800
rect 18491 26745 18517 26775
rect 18645 26745 18690 26775
rect 18660 26742 18690 26745
rect 18832 26745 18877 26775
rect 18961 26745 18987 26775
rect 18832 26742 18862 26745
rect 18660 26732 18862 26742
rect 18660 26712 18759 26732
rect 18743 26698 18759 26712
rect 18793 26712 18862 26732
rect 18793 26698 18809 26712
rect 18743 26688 18809 26698
rect 18493 26091 18519 26121
rect 18719 26101 18839 26121
rect 18719 26091 18767 26101
rect 18751 26067 18767 26091
rect 18801 26091 18839 26101
rect 18969 26091 18995 26121
rect 18801 26067 18817 26091
rect 18751 26057 18817 26067
rect 18493 25994 18519 26024
rect 18647 26015 18713 26024
rect 18846 26015 18885 26026
rect 18647 25996 18885 26015
rect 18969 25996 18995 26026
rect 18647 25994 18870 25996
rect 18683 25985 18870 25994
rect 18751 25840 18817 25985
rect 18751 25836 18767 25840
rect 18493 25806 18519 25836
rect 18719 25806 18767 25836
rect 18801 25838 18817 25840
rect 18801 25808 18839 25838
rect 18969 25808 18995 25838
rect 18801 25806 18817 25808
rect 18751 25796 18817 25806
rect 18751 25752 18839 25754
rect 18493 25722 18519 25752
rect 18719 25724 18839 25752
rect 18969 25724 18995 25754
rect 18719 25722 18817 25724
rect 18751 25656 18817 25722
rect 18751 25622 18767 25656
rect 18801 25622 18817 25656
rect 18751 25612 18817 25622
rect 18635 25582 18701 25592
rect 18635 25548 18651 25582
rect 18685 25564 18701 25582
rect 18685 25548 18885 25564
rect 18635 25541 18885 25548
rect 18493 25511 18519 25541
rect 18603 25534 18885 25541
rect 18969 25534 18995 25564
rect 18603 25511 18701 25534
rect 18641 25446 18695 25462
rect 18641 25427 18651 25446
rect 18493 25397 18519 25427
rect 18603 25412 18651 25427
rect 18685 25412 18695 25446
rect 18603 25397 18695 25412
rect 18641 25396 18695 25397
rect 18737 25439 18897 25469
rect 18969 25439 18995 25469
rect 18737 25354 18767 25439
rect 18701 25344 18767 25354
rect 18701 25343 18717 25344
rect 18493 25313 18519 25343
rect 18603 25313 18717 25343
rect 18701 25310 18717 25313
rect 18751 25310 18767 25344
rect 18809 25387 18875 25397
rect 18809 25353 18825 25387
rect 18859 25363 18875 25387
rect 18859 25353 18897 25363
rect 18809 25333 18897 25353
rect 18969 25333 18995 25363
rect 18701 25300 18767 25310
rect 18796 25248 18841 25262
rect 18493 25218 18519 25248
rect 18669 25232 18841 25248
rect 18969 25232 18995 25262
rect 18669 25218 18826 25232
rect 18707 25208 18761 25218
rect 18707 25174 18717 25208
rect 18751 25174 18761 25208
rect 18707 25158 18761 25174
rect 18803 25144 18857 25160
rect 18803 25116 18813 25144
rect 18493 25086 18519 25116
rect 18603 25110 18813 25116
rect 18847 25143 18857 25144
rect 18847 25113 18885 25143
rect 18969 25113 18995 25143
rect 18847 25110 18857 25113
rect 18603 25086 18857 25110
rect 18635 25034 18701 25044
rect 18635 25013 18651 25034
rect 18493 24983 18519 25013
rect 18603 25000 18651 25013
rect 18685 25000 18701 25034
rect 18603 24983 18701 25000
rect 18743 25014 18897 25044
rect 18969 25014 18995 25044
rect 18743 24941 18773 25014
rect 18719 24925 18773 24941
rect 18719 24918 18729 24925
rect 18493 24888 18519 24918
rect 18603 24891 18729 24918
rect 18763 24891 18773 24925
rect 18815 24945 18869 24961
rect 18815 24911 18825 24945
rect 18859 24915 18897 24945
rect 18969 24915 18995 24945
rect 18859 24911 18869 24915
rect 18815 24895 18869 24911
rect 18603 24888 18773 24891
rect 18719 24875 18773 24888
rect 18493 24803 18519 24833
rect 18603 24803 18885 24833
rect 18969 24803 18995 24833
rect 18683 24782 18749 24803
rect 18683 24748 18699 24782
rect 18733 24748 18749 24782
rect 18683 24738 18749 24748
rect 18499 24615 18525 24645
rect 18653 24620 18885 24645
rect 18653 24615 18752 24620
rect 18742 24586 18752 24615
rect 18786 24615 18885 24620
rect 18969 24615 18995 24645
rect 18786 24586 18796 24615
rect 18742 24570 18796 24586
rect 18499 24531 18525 24561
rect 18653 24531 18698 24561
rect 18668 24528 18698 24531
rect 18840 24531 18885 24561
rect 18969 24531 18995 24561
rect 18840 24528 18870 24531
rect 18668 24518 18870 24528
rect 18668 24498 18767 24518
rect 18751 24484 18767 24498
rect 18801 24498 18870 24518
rect 18801 24484 18817 24498
rect 18751 24474 18817 24484
rect 7625 23335 7655 23361
rect 7709 23335 7739 23361
rect 7897 23341 7927 23367
rect 7982 23341 8012 23367
rect 8077 23341 8107 23367
rect 8180 23341 8210 23367
rect 8312 23341 8342 23367
rect 8407 23341 8437 23367
rect 8491 23341 8521 23367
rect 8605 23341 8635 23367
rect 8816 23341 8846 23367
rect 8900 23341 8930 23367
rect 9088 23341 9118 23367
rect 9185 23341 9215 23367
rect 9839 23343 9869 23369
rect 9923 23343 9953 23369
rect 10111 23349 10141 23375
rect 10196 23349 10226 23375
rect 10291 23349 10321 23375
rect 10394 23349 10424 23375
rect 10526 23349 10556 23375
rect 10621 23349 10651 23375
rect 10705 23349 10735 23375
rect 10819 23349 10849 23375
rect 11030 23349 11060 23375
rect 11114 23349 11144 23375
rect 11302 23349 11332 23375
rect 11399 23349 11429 23375
rect 7625 23192 7655 23207
rect 7592 23162 7655 23192
rect 7592 23109 7622 23162
rect 7709 23118 7739 23207
rect 7897 23177 7927 23257
rect 7568 23093 7622 23109
rect 7568 23059 7578 23093
rect 7612 23059 7622 23093
rect 7664 23108 7739 23118
rect 7832 23161 7927 23177
rect 7832 23127 7842 23161
rect 7876 23127 7927 23161
rect 7982 23141 8012 23257
rect 8077 23225 8107 23257
rect 8077 23209 8138 23225
rect 8077 23175 8094 23209
rect 8128 23175 8138 23209
rect 8077 23159 8138 23175
rect 7832 23111 7927 23127
rect 7664 23074 7680 23108
rect 7714 23074 7739 23108
rect 7664 23064 7739 23074
rect 7568 23043 7622 23059
rect 7592 23020 7622 23043
rect 7592 22990 7655 23020
rect 7625 22975 7655 22990
rect 7709 22975 7739 23064
rect 7897 22975 7927 23111
rect 7969 23131 8035 23141
rect 7969 23097 7985 23131
rect 8019 23117 8035 23131
rect 8019 23097 8138 23117
rect 7969 23087 8138 23097
rect 7989 23035 8055 23045
rect 7989 23001 8005 23035
rect 8039 23001 8055 23035
rect 7989 22991 8055 23001
rect 8009 22963 8039 22991
rect 8108 22963 8138 23087
rect 8180 23057 8210 23257
rect 8312 23153 8342 23191
rect 8407 23159 8437 23257
rect 8491 23219 8521 23257
rect 8605 23225 8635 23257
rect 8490 23209 8556 23219
rect 8490 23175 8506 23209
rect 8540 23175 8556 23209
rect 8490 23165 8556 23175
rect 8605 23209 8686 23225
rect 8605 23175 8642 23209
rect 8676 23175 8686 23209
rect 8605 23159 8686 23175
rect 8252 23143 8342 23153
rect 8252 23109 8268 23143
rect 8302 23109 8342 23143
rect 8252 23099 8342 23109
rect 8312 23064 8342 23099
rect 8394 23143 8448 23159
rect 8394 23109 8404 23143
rect 8438 23123 8448 23143
rect 8438 23109 8563 23123
rect 8394 23093 8563 23109
rect 8180 23047 8254 23057
rect 8180 23013 8204 23047
rect 8238 23013 8254 23047
rect 8312 23034 8356 23064
rect 8326 23019 8356 23034
rect 8427 23035 8491 23051
rect 8180 23003 8254 23013
rect 8207 22975 8237 23003
rect 8427 23001 8447 23035
rect 8481 23001 8491 23035
rect 8427 22985 8491 23001
rect 8427 22963 8457 22985
rect 8533 22963 8563 23093
rect 8628 22975 8658 23159
rect 9088 23177 9118 23213
rect 9079 23147 9118 23177
rect 8816 23109 8846 23141
rect 8900 23109 8930 23141
rect 9079 23109 9109 23147
rect 9839 23200 9869 23215
rect 9806 23170 9869 23200
rect 9185 23109 9215 23141
rect 9806 23117 9836 23170
rect 9923 23126 9953 23215
rect 10111 23185 10141 23265
rect 8706 23093 8848 23109
rect 8706 23059 8716 23093
rect 8750 23059 8848 23093
rect 8706 23043 8848 23059
rect 8890 23093 9109 23109
rect 8890 23059 8900 23093
rect 8934 23059 9109 23093
rect 8890 23043 9109 23059
rect 9151 23093 9215 23109
rect 9151 23059 9161 23093
rect 9195 23059 9215 23093
rect 9151 23043 9215 23059
rect 9782 23101 9836 23117
rect 9782 23067 9792 23101
rect 9826 23067 9836 23101
rect 9878 23116 9953 23126
rect 10046 23169 10141 23185
rect 10046 23135 10056 23169
rect 10090 23135 10141 23169
rect 10196 23149 10226 23265
rect 10291 23233 10321 23265
rect 10291 23217 10352 23233
rect 10291 23183 10308 23217
rect 10342 23183 10352 23217
rect 10291 23167 10352 23183
rect 10046 23119 10141 23135
rect 9878 23082 9894 23116
rect 9928 23082 9953 23116
rect 9878 23072 9953 23082
rect 9782 23051 9836 23067
rect 8818 23021 8848 23043
rect 8902 23021 8932 23043
rect 9079 23014 9109 23043
rect 9185 23021 9215 23043
rect 9806 23028 9836 23051
rect 9079 22990 9120 23014
rect 9090 22975 9120 22990
rect 9806 22998 9869 23028
rect 9839 22983 9869 22998
rect 9923 22983 9953 23072
rect 10111 22983 10141 23119
rect 10183 23139 10249 23149
rect 10183 23105 10199 23139
rect 10233 23125 10249 23139
rect 10233 23105 10352 23125
rect 10183 23095 10352 23105
rect 10203 23043 10269 23053
rect 10203 23009 10219 23043
rect 10253 23009 10269 23043
rect 10203 22999 10269 23009
rect 10223 22971 10253 22999
rect 10322 22971 10352 23095
rect 10394 23065 10424 23265
rect 10526 23161 10556 23199
rect 10621 23167 10651 23265
rect 10705 23227 10735 23265
rect 10819 23233 10849 23265
rect 10704 23217 10770 23227
rect 10704 23183 10720 23217
rect 10754 23183 10770 23217
rect 10704 23173 10770 23183
rect 10819 23217 10900 23233
rect 10819 23183 10856 23217
rect 10890 23183 10900 23217
rect 10819 23167 10900 23183
rect 10466 23151 10556 23161
rect 10466 23117 10482 23151
rect 10516 23117 10556 23151
rect 10466 23107 10556 23117
rect 10526 23072 10556 23107
rect 10608 23151 10662 23167
rect 10608 23117 10618 23151
rect 10652 23131 10662 23151
rect 10652 23117 10777 23131
rect 10608 23101 10777 23117
rect 10394 23055 10468 23065
rect 10394 23021 10418 23055
rect 10452 23021 10468 23055
rect 10526 23042 10570 23072
rect 10540 23027 10570 23042
rect 10641 23043 10705 23059
rect 10394 23011 10468 23021
rect 10421 22983 10451 23011
rect 10641 23009 10661 23043
rect 10695 23009 10705 23043
rect 10641 22993 10705 23009
rect 10641 22971 10671 22993
rect 10747 22971 10777 23101
rect 10842 22983 10872 23167
rect 11302 23185 11332 23221
rect 11293 23155 11332 23185
rect 11030 23117 11060 23149
rect 11114 23117 11144 23149
rect 11293 23117 11323 23155
rect 12039 23325 12069 23351
rect 12123 23325 12153 23351
rect 12311 23331 12341 23357
rect 12396 23331 12426 23357
rect 12491 23331 12521 23357
rect 12594 23331 12624 23357
rect 12726 23331 12756 23357
rect 12821 23331 12851 23357
rect 12905 23331 12935 23357
rect 13019 23331 13049 23357
rect 13230 23331 13260 23357
rect 13314 23331 13344 23357
rect 13502 23331 13532 23357
rect 13599 23331 13629 23357
rect 14253 23333 14283 23359
rect 14337 23333 14367 23359
rect 14525 23339 14555 23365
rect 14610 23339 14640 23365
rect 14705 23339 14735 23365
rect 14808 23339 14838 23365
rect 14940 23339 14970 23365
rect 15035 23339 15065 23365
rect 15119 23339 15149 23365
rect 15233 23339 15263 23365
rect 15444 23339 15474 23365
rect 15528 23339 15558 23365
rect 15716 23339 15746 23365
rect 15813 23339 15843 23365
rect 16559 23341 16589 23367
rect 16643 23341 16673 23367
rect 16831 23347 16861 23373
rect 16916 23347 16946 23373
rect 17011 23347 17041 23373
rect 17114 23347 17144 23373
rect 17246 23347 17276 23373
rect 17341 23347 17371 23373
rect 17425 23347 17455 23373
rect 17539 23347 17569 23373
rect 17750 23347 17780 23373
rect 17834 23347 17864 23373
rect 18022 23347 18052 23373
rect 18119 23347 18149 23373
rect 12039 23182 12069 23197
rect 12006 23152 12069 23182
rect 11399 23117 11429 23149
rect 10920 23101 11062 23117
rect 10920 23067 10930 23101
rect 10964 23067 11062 23101
rect 10920 23051 11062 23067
rect 11104 23101 11323 23117
rect 11104 23067 11114 23101
rect 11148 23067 11323 23101
rect 11104 23051 11323 23067
rect 11365 23101 11429 23117
rect 11365 23067 11375 23101
rect 11409 23067 11429 23101
rect 12006 23099 12036 23152
rect 12123 23108 12153 23197
rect 12311 23167 12341 23247
rect 11365 23051 11429 23067
rect 11032 23029 11062 23051
rect 11116 23029 11146 23051
rect 11293 23022 11323 23051
rect 11399 23029 11429 23051
rect 11982 23083 12036 23099
rect 11982 23049 11992 23083
rect 12026 23049 12036 23083
rect 12078 23098 12153 23108
rect 12246 23151 12341 23167
rect 12246 23117 12256 23151
rect 12290 23117 12341 23151
rect 12396 23131 12426 23247
rect 12491 23215 12521 23247
rect 12491 23199 12552 23215
rect 12491 23165 12508 23199
rect 12542 23165 12552 23199
rect 12491 23149 12552 23165
rect 12246 23101 12341 23117
rect 12078 23064 12094 23098
rect 12128 23064 12153 23098
rect 12078 23054 12153 23064
rect 11982 23033 12036 23049
rect 11293 22998 11334 23022
rect 11304 22983 11334 22998
rect 12006 23010 12036 23033
rect 12006 22980 12069 23010
rect 12039 22965 12069 22980
rect 12123 22965 12153 23054
rect 12311 22965 12341 23101
rect 12383 23121 12449 23131
rect 12383 23087 12399 23121
rect 12433 23107 12449 23121
rect 12433 23087 12552 23107
rect 12383 23077 12552 23087
rect 12403 23025 12469 23035
rect 12403 22991 12419 23025
rect 12453 22991 12469 23025
rect 12403 22981 12469 22991
rect 7625 22865 7655 22891
rect 7709 22865 7739 22891
rect 7897 22865 7927 22891
rect 8009 22865 8039 22891
rect 8108 22865 8138 22891
rect 8207 22865 8237 22891
rect 8326 22865 8356 22891
rect 8427 22865 8457 22891
rect 8533 22865 8563 22891
rect 8628 22865 8658 22891
rect 8818 22865 8848 22891
rect 8902 22865 8932 22891
rect 9090 22865 9120 22891
rect 9185 22865 9215 22891
rect 9839 22873 9869 22899
rect 9923 22873 9953 22899
rect 10111 22873 10141 22899
rect 10223 22873 10253 22899
rect 10322 22873 10352 22899
rect 10421 22873 10451 22899
rect 10540 22873 10570 22899
rect 10641 22873 10671 22899
rect 10747 22873 10777 22899
rect 10842 22873 10872 22899
rect 11032 22873 11062 22899
rect 11116 22873 11146 22899
rect 11304 22873 11334 22899
rect 11399 22873 11429 22899
rect 12423 22953 12453 22981
rect 12522 22953 12552 23077
rect 12594 23047 12624 23247
rect 12726 23143 12756 23181
rect 12821 23149 12851 23247
rect 12905 23209 12935 23247
rect 13019 23215 13049 23247
rect 12904 23199 12970 23209
rect 12904 23165 12920 23199
rect 12954 23165 12970 23199
rect 12904 23155 12970 23165
rect 13019 23199 13100 23215
rect 13019 23165 13056 23199
rect 13090 23165 13100 23199
rect 13019 23149 13100 23165
rect 12666 23133 12756 23143
rect 12666 23099 12682 23133
rect 12716 23099 12756 23133
rect 12666 23089 12756 23099
rect 12726 23054 12756 23089
rect 12808 23133 12862 23149
rect 12808 23099 12818 23133
rect 12852 23113 12862 23133
rect 12852 23099 12977 23113
rect 12808 23083 12977 23099
rect 12594 23037 12668 23047
rect 12594 23003 12618 23037
rect 12652 23003 12668 23037
rect 12726 23024 12770 23054
rect 12740 23009 12770 23024
rect 12841 23025 12905 23041
rect 12594 22993 12668 23003
rect 12621 22965 12651 22993
rect 12841 22991 12861 23025
rect 12895 22991 12905 23025
rect 12841 22975 12905 22991
rect 12841 22953 12871 22975
rect 12947 22953 12977 23083
rect 13042 22965 13072 23149
rect 13502 23167 13532 23203
rect 13493 23137 13532 23167
rect 13230 23099 13260 23131
rect 13314 23099 13344 23131
rect 13493 23099 13523 23137
rect 14253 23190 14283 23205
rect 14220 23160 14283 23190
rect 13599 23099 13629 23131
rect 14220 23107 14250 23160
rect 14337 23116 14367 23205
rect 14525 23175 14555 23255
rect 13120 23083 13262 23099
rect 13120 23049 13130 23083
rect 13164 23049 13262 23083
rect 13120 23033 13262 23049
rect 13304 23083 13523 23099
rect 13304 23049 13314 23083
rect 13348 23049 13523 23083
rect 13304 23033 13523 23049
rect 13565 23083 13629 23099
rect 13565 23049 13575 23083
rect 13609 23049 13629 23083
rect 13565 23033 13629 23049
rect 14196 23091 14250 23107
rect 14196 23057 14206 23091
rect 14240 23057 14250 23091
rect 14292 23106 14367 23116
rect 14460 23159 14555 23175
rect 14460 23125 14470 23159
rect 14504 23125 14555 23159
rect 14610 23139 14640 23255
rect 14705 23223 14735 23255
rect 14705 23207 14766 23223
rect 14705 23173 14722 23207
rect 14756 23173 14766 23207
rect 14705 23157 14766 23173
rect 14460 23109 14555 23125
rect 14292 23072 14308 23106
rect 14342 23072 14367 23106
rect 14292 23062 14367 23072
rect 14196 23041 14250 23057
rect 13232 23011 13262 23033
rect 13316 23011 13346 23033
rect 13493 23004 13523 23033
rect 13599 23011 13629 23033
rect 14220 23018 14250 23041
rect 13493 22980 13534 23004
rect 13504 22965 13534 22980
rect 14220 22988 14283 23018
rect 14253 22973 14283 22988
rect 14337 22973 14367 23062
rect 14525 22973 14555 23109
rect 14597 23129 14663 23139
rect 14597 23095 14613 23129
rect 14647 23115 14663 23129
rect 14647 23095 14766 23115
rect 14597 23085 14766 23095
rect 14617 23033 14683 23043
rect 14617 22999 14633 23033
rect 14667 22999 14683 23033
rect 14617 22989 14683 22999
rect 14637 22961 14667 22989
rect 14736 22961 14766 23085
rect 14808 23055 14838 23255
rect 14940 23151 14970 23189
rect 15035 23157 15065 23255
rect 15119 23217 15149 23255
rect 15233 23223 15263 23255
rect 15118 23207 15184 23217
rect 15118 23173 15134 23207
rect 15168 23173 15184 23207
rect 15118 23163 15184 23173
rect 15233 23207 15314 23223
rect 15233 23173 15270 23207
rect 15304 23173 15314 23207
rect 15233 23157 15314 23173
rect 14880 23141 14970 23151
rect 14880 23107 14896 23141
rect 14930 23107 14970 23141
rect 14880 23097 14970 23107
rect 14940 23062 14970 23097
rect 15022 23141 15076 23157
rect 15022 23107 15032 23141
rect 15066 23121 15076 23141
rect 15066 23107 15191 23121
rect 15022 23091 15191 23107
rect 14808 23045 14882 23055
rect 14808 23011 14832 23045
rect 14866 23011 14882 23045
rect 14940 23032 14984 23062
rect 14954 23017 14984 23032
rect 15055 23033 15119 23049
rect 14808 23001 14882 23011
rect 14835 22973 14865 23001
rect 15055 22999 15075 23033
rect 15109 22999 15119 23033
rect 15055 22983 15119 22999
rect 15055 22961 15085 22983
rect 15161 22961 15191 23091
rect 15256 22973 15286 23157
rect 15716 23175 15746 23211
rect 15707 23145 15746 23175
rect 15444 23107 15474 23139
rect 15528 23107 15558 23139
rect 15707 23107 15737 23145
rect 16559 23198 16589 23213
rect 16526 23168 16589 23198
rect 15813 23107 15843 23139
rect 16526 23115 16556 23168
rect 16643 23124 16673 23213
rect 16831 23183 16861 23263
rect 15334 23091 15476 23107
rect 15334 23057 15344 23091
rect 15378 23057 15476 23091
rect 15334 23041 15476 23057
rect 15518 23091 15737 23107
rect 15518 23057 15528 23091
rect 15562 23057 15737 23091
rect 15518 23041 15737 23057
rect 15779 23091 15843 23107
rect 15779 23057 15789 23091
rect 15823 23057 15843 23091
rect 15779 23041 15843 23057
rect 16502 23099 16556 23115
rect 16502 23065 16512 23099
rect 16546 23065 16556 23099
rect 16598 23114 16673 23124
rect 16766 23167 16861 23183
rect 16766 23133 16776 23167
rect 16810 23133 16861 23167
rect 16916 23147 16946 23263
rect 17011 23231 17041 23263
rect 17011 23215 17072 23231
rect 17011 23181 17028 23215
rect 17062 23181 17072 23215
rect 17011 23165 17072 23181
rect 16766 23117 16861 23133
rect 16598 23080 16614 23114
rect 16648 23080 16673 23114
rect 16598 23070 16673 23080
rect 16502 23049 16556 23065
rect 15446 23019 15476 23041
rect 15530 23019 15560 23041
rect 15707 23012 15737 23041
rect 15813 23019 15843 23041
rect 16526 23026 16556 23049
rect 15707 22988 15748 23012
rect 15718 22973 15748 22988
rect 16526 22996 16589 23026
rect 16559 22981 16589 22996
rect 16643 22981 16673 23070
rect 16831 22981 16861 23117
rect 16903 23137 16969 23147
rect 16903 23103 16919 23137
rect 16953 23123 16969 23137
rect 16953 23103 17072 23123
rect 16903 23093 17072 23103
rect 16923 23041 16989 23051
rect 16923 23007 16939 23041
rect 16973 23007 16989 23041
rect 16923 22997 16989 23007
rect 16943 22969 16973 22997
rect 17042 22969 17072 23093
rect 17114 23063 17144 23263
rect 17246 23159 17276 23197
rect 17341 23165 17371 23263
rect 17425 23225 17455 23263
rect 17539 23231 17569 23263
rect 17424 23215 17490 23225
rect 17424 23181 17440 23215
rect 17474 23181 17490 23215
rect 17424 23171 17490 23181
rect 17539 23215 17620 23231
rect 17539 23181 17576 23215
rect 17610 23181 17620 23215
rect 17539 23165 17620 23181
rect 17186 23149 17276 23159
rect 17186 23115 17202 23149
rect 17236 23115 17276 23149
rect 17186 23105 17276 23115
rect 17246 23070 17276 23105
rect 17328 23149 17382 23165
rect 17328 23115 17338 23149
rect 17372 23129 17382 23149
rect 17372 23115 17497 23129
rect 17328 23099 17497 23115
rect 17114 23053 17188 23063
rect 17114 23019 17138 23053
rect 17172 23019 17188 23053
rect 17246 23040 17290 23070
rect 17260 23025 17290 23040
rect 17361 23041 17425 23057
rect 17114 23009 17188 23019
rect 17141 22981 17171 23009
rect 17361 23007 17381 23041
rect 17415 23007 17425 23041
rect 17361 22991 17425 23007
rect 17361 22969 17391 22991
rect 17467 22969 17497 23099
rect 17562 22981 17592 23165
rect 18022 23183 18052 23219
rect 18013 23153 18052 23183
rect 17750 23115 17780 23147
rect 17834 23115 17864 23147
rect 18013 23115 18043 23153
rect 18119 23115 18149 23147
rect 17640 23099 17782 23115
rect 17640 23065 17650 23099
rect 17684 23065 17782 23099
rect 17640 23049 17782 23065
rect 17824 23099 18043 23115
rect 17824 23065 17834 23099
rect 17868 23065 18043 23099
rect 17824 23049 18043 23065
rect 18085 23099 18149 23115
rect 18085 23065 18095 23099
rect 18129 23065 18149 23099
rect 18085 23049 18149 23065
rect 17752 23027 17782 23049
rect 17836 23027 17866 23049
rect 18013 23020 18043 23049
rect 18119 23027 18149 23049
rect 18013 22996 18054 23020
rect 18024 22981 18054 22996
rect 12039 22855 12069 22881
rect 12123 22855 12153 22881
rect 12311 22855 12341 22881
rect 12423 22855 12453 22881
rect 12522 22855 12552 22881
rect 12621 22855 12651 22881
rect 12740 22855 12770 22881
rect 12841 22855 12871 22881
rect 12947 22855 12977 22881
rect 13042 22855 13072 22881
rect 13232 22855 13262 22881
rect 13316 22855 13346 22881
rect 13504 22855 13534 22881
rect 13599 22855 13629 22881
rect 14253 22863 14283 22889
rect 14337 22863 14367 22889
rect 14525 22863 14555 22889
rect 14637 22863 14667 22889
rect 14736 22863 14766 22889
rect 14835 22863 14865 22889
rect 14954 22863 14984 22889
rect 15055 22863 15085 22889
rect 15161 22863 15191 22889
rect 15256 22863 15286 22889
rect 15446 22863 15476 22889
rect 15530 22863 15560 22889
rect 15718 22863 15748 22889
rect 15813 22863 15843 22889
rect 16559 22871 16589 22897
rect 16643 22871 16673 22897
rect 16831 22871 16861 22897
rect 16943 22871 16973 22897
rect 17042 22871 17072 22897
rect 17141 22871 17171 22897
rect 17260 22871 17290 22897
rect 17361 22871 17391 22897
rect 17467 22871 17497 22897
rect 17562 22871 17592 22897
rect 17752 22871 17782 22897
rect 17836 22871 17866 22897
rect 18024 22871 18054 22897
rect 18119 22871 18149 22897
rect 16471 17637 16501 17663
rect 17345 17639 17375 17665
rect 15693 17599 15723 17625
rect 18113 17629 18143 17655
rect 19235 17631 19265 17657
rect 20109 17633 20139 17659
rect 16471 17485 16501 17507
rect 17345 17487 17375 17509
rect 20877 17623 20907 17649
rect 16471 17469 16557 17485
rect 15693 17447 15723 17469
rect 15693 17431 15779 17447
rect 15693 17397 15729 17431
rect 15763 17397 15779 17431
rect 15693 17381 15779 17397
rect 16471 17435 16507 17469
rect 16541 17435 16557 17469
rect 16471 17419 16557 17435
rect 17345 17471 17431 17487
rect 17345 17437 17381 17471
rect 17415 17437 17431 17471
rect 17345 17421 17431 17437
rect 18113 17477 18143 17499
rect 19235 17479 19265 17501
rect 20109 17481 20139 17503
rect 21491 17621 21521 17647
rect 22365 17623 22395 17649
rect 18113 17461 18199 17477
rect 18113 17427 18149 17461
rect 18183 17427 18199 17461
rect 16471 17387 16501 17419
rect 17345 17389 17375 17421
rect 18113 17411 18199 17427
rect 19235 17463 19321 17479
rect 19235 17429 19271 17463
rect 19305 17429 19321 17463
rect 19235 17413 19321 17429
rect 20109 17465 20195 17481
rect 20109 17431 20145 17465
rect 20179 17431 20195 17465
rect 20109 17415 20195 17431
rect 20877 17471 20907 17493
rect 23133 17613 23163 17639
rect 20877 17455 20963 17471
rect 20877 17421 20913 17455
rect 20947 17421 20963 17455
rect 15693 17349 15723 17381
rect 18113 17379 18143 17411
rect 19235 17381 19265 17413
rect 20109 17383 20139 17415
rect 20877 17405 20963 17421
rect 21491 17469 21521 17491
rect 22365 17471 22395 17493
rect 21491 17453 21577 17469
rect 21491 17419 21527 17453
rect 21561 17419 21577 17453
rect 16471 17161 16501 17187
rect 17345 17163 17375 17189
rect 20877 17373 20907 17405
rect 21491 17403 21577 17419
rect 22365 17455 22451 17471
rect 22365 17421 22401 17455
rect 22435 17421 22451 17455
rect 22365 17405 22451 17421
rect 23133 17461 23163 17483
rect 23133 17445 23219 17461
rect 23133 17411 23169 17445
rect 23203 17411 23219 17445
rect 18113 17153 18143 17179
rect 19235 17155 19265 17181
rect 20109 17157 20139 17183
rect 21491 17371 21521 17403
rect 22365 17373 22395 17405
rect 23133 17395 23219 17411
rect 15693 17123 15723 17149
rect 20877 17147 20907 17173
rect 23133 17363 23163 17395
rect 21491 17145 21521 17171
rect 22365 17147 22395 17173
rect 23133 17137 23163 17163
rect 9421 16543 9451 16569
rect 9505 16543 9535 16569
rect 9589 16543 9619 16569
rect 9673 16543 9703 16569
rect 9861 16543 9891 16569
rect 9421 16311 9451 16343
rect 9505 16311 9535 16343
rect 9589 16311 9619 16343
rect 9673 16311 9703 16343
rect 9861 16311 9891 16343
rect 9409 16295 9463 16311
rect 9409 16261 9419 16295
rect 9453 16261 9463 16295
rect 9409 16245 9463 16261
rect 9505 16295 9619 16311
rect 9505 16261 9536 16295
rect 9570 16261 9619 16295
rect 9505 16245 9619 16261
rect 9661 16295 9715 16311
rect 9661 16261 9671 16295
rect 9705 16261 9715 16295
rect 9661 16245 9715 16261
rect 9757 16295 9891 16311
rect 9757 16261 9767 16295
rect 9801 16278 9891 16295
rect 9801 16261 9887 16278
rect 9757 16245 9887 16261
rect 9421 16223 9451 16245
rect 9505 16223 9535 16245
rect 9589 16223 9619 16245
rect 9673 16223 9703 16245
rect 9857 16223 9887 16245
rect 9421 16067 9451 16093
rect 9505 16067 9535 16093
rect 9589 16067 9619 16093
rect 9673 16067 9703 16093
rect 9857 16067 9887 16093
rect 9739 15799 9769 15825
rect 9547 15757 9577 15783
rect 9631 15757 9661 15783
rect 9547 15567 9577 15673
rect 9490 15551 9577 15567
rect 9490 15517 9506 15551
rect 9540 15517 9577 15551
rect 9490 15501 9577 15517
rect 9547 15461 9577 15501
rect 9631 15567 9661 15673
rect 11553 15689 11583 15715
rect 11653 15689 11683 15715
rect 11757 15689 11787 15715
rect 11843 15689 11873 15715
rect 12009 15689 12039 15715
rect 9739 15567 9769 15599
rect 9631 15551 9697 15567
rect 9631 15517 9647 15551
rect 9681 15517 9697 15551
rect 9631 15501 9697 15517
rect 9739 15551 9805 15567
rect 9739 15517 9755 15551
rect 9789 15517 9805 15551
rect 9739 15501 9805 15517
rect 9631 15461 9661 15501
rect 9739 15479 9769 15501
rect 9547 15351 9577 15377
rect 9631 15351 9661 15377
rect 11553 15457 11583 15605
rect 11653 15457 11683 15605
rect 11757 15457 11787 15605
rect 11843 15457 11873 15605
rect 12009 15457 12039 15489
rect 11495 15441 11583 15457
rect 11495 15407 11505 15441
rect 11539 15407 11583 15441
rect 11495 15391 11583 15407
rect 9739 15323 9769 15349
rect 11553 15323 11583 15391
rect 11641 15441 11695 15457
rect 11641 15407 11651 15441
rect 11685 15407 11695 15441
rect 11641 15391 11695 15407
rect 11747 15441 11801 15457
rect 11747 15407 11757 15441
rect 11791 15407 11801 15441
rect 11747 15391 11801 15407
rect 11843 15441 11907 15457
rect 11843 15407 11853 15441
rect 11887 15407 11907 15441
rect 11843 15391 11907 15407
rect 11954 15441 12039 15457
rect 11954 15407 11964 15441
rect 11998 15407 12039 15441
rect 11954 15391 12039 15407
rect 11641 15323 11671 15391
rect 11747 15323 11777 15391
rect 11843 15323 11873 15391
rect 12009 15369 12039 15391
rect 10923 15189 10953 15215
rect 11553 15213 11583 15239
rect 11641 15213 11671 15239
rect 11747 15213 11777 15239
rect 11843 15213 11873 15239
rect 12009 15213 12039 15239
rect 10731 15147 10761 15173
rect 10815 15147 10845 15173
rect 9431 14979 9461 15005
rect 9515 14979 9545 15005
rect 9599 14979 9629 15005
rect 9683 14979 9713 15005
rect 9871 14979 9901 15005
rect 10731 14957 10761 15063
rect 10674 14941 10761 14957
rect 10674 14907 10690 14941
rect 10724 14907 10761 14941
rect 10674 14891 10761 14907
rect 10731 14851 10761 14891
rect 10815 14957 10845 15063
rect 10923 14957 10953 14989
rect 10815 14941 10881 14957
rect 10815 14907 10831 14941
rect 10865 14907 10881 14941
rect 10815 14891 10881 14907
rect 10923 14941 10989 14957
rect 10923 14907 10939 14941
rect 10973 14907 10989 14941
rect 10923 14891 10989 14907
rect 10815 14851 10845 14891
rect 10923 14869 10953 14891
rect 9431 14747 9461 14779
rect 9515 14747 9545 14779
rect 9599 14747 9629 14779
rect 9683 14747 9713 14779
rect 9871 14747 9901 14779
rect 9419 14731 9473 14747
rect 9419 14697 9429 14731
rect 9463 14697 9473 14731
rect 9419 14681 9473 14697
rect 9515 14731 9629 14747
rect 9515 14697 9546 14731
rect 9580 14697 9629 14731
rect 9515 14681 9629 14697
rect 9671 14731 9725 14747
rect 9671 14697 9681 14731
rect 9715 14697 9725 14731
rect 9671 14681 9725 14697
rect 9767 14731 9901 14747
rect 10731 14741 10761 14767
rect 10815 14741 10845 14767
rect 9767 14697 9777 14731
rect 9811 14714 9901 14731
rect 9811 14697 9897 14714
rect 10923 14713 10953 14739
rect 9767 14681 9897 14697
rect 9431 14659 9461 14681
rect 9515 14659 9545 14681
rect 9599 14659 9629 14681
rect 9683 14659 9713 14681
rect 9867 14659 9897 14681
rect 9431 14503 9461 14529
rect 9515 14503 9545 14529
rect 9599 14503 9629 14529
rect 9683 14503 9713 14529
rect 9867 14503 9897 14529
rect 9749 14235 9779 14261
rect 9557 14193 9587 14219
rect 9641 14193 9671 14219
rect 9557 14003 9587 14109
rect 9500 13987 9587 14003
rect 9500 13953 9516 13987
rect 9550 13953 9587 13987
rect 9500 13937 9587 13953
rect 9557 13897 9587 13937
rect 9641 14003 9671 14109
rect 10769 14223 10799 14249
rect 10869 14223 10899 14249
rect 10973 14223 11003 14249
rect 11059 14223 11089 14249
rect 11225 14223 11255 14249
rect 9749 14003 9779 14035
rect 9641 13987 9707 14003
rect 9641 13953 9657 13987
rect 9691 13953 9707 13987
rect 9641 13937 9707 13953
rect 9749 13987 9815 14003
rect 10769 13991 10799 14139
rect 10869 13991 10899 14139
rect 10973 13991 11003 14139
rect 11059 13991 11089 14139
rect 13029 14207 13059 14233
rect 12829 14183 12895 14193
rect 12829 14149 12845 14183
rect 12879 14149 12895 14183
rect 12829 14139 12895 14149
rect 12667 14091 12697 14117
rect 12763 14091 12793 14117
rect 12835 14091 12865 14139
rect 12931 14091 12961 14117
rect 11225 13991 11255 14023
rect 9749 13953 9765 13987
rect 9799 13953 9815 13987
rect 9749 13937 9815 13953
rect 10711 13975 10799 13991
rect 10711 13941 10721 13975
rect 10755 13941 10799 13975
rect 9641 13897 9671 13937
rect 9749 13915 9779 13937
rect 10711 13925 10799 13941
rect 9557 13787 9587 13813
rect 9641 13787 9671 13813
rect 10769 13857 10799 13925
rect 10857 13975 10911 13991
rect 10857 13941 10867 13975
rect 10901 13941 10911 13975
rect 10857 13925 10911 13941
rect 10963 13975 11017 13991
rect 10963 13941 10973 13975
rect 11007 13941 11017 13975
rect 10963 13925 11017 13941
rect 11059 13975 11123 13991
rect 11059 13941 11069 13975
rect 11103 13941 11123 13975
rect 11059 13925 11123 13941
rect 11170 13975 11255 13991
rect 12667 13975 12697 14007
rect 12763 13975 12793 14007
rect 11170 13941 11180 13975
rect 11214 13941 11255 13975
rect 11170 13925 11255 13941
rect 10857 13857 10887 13925
rect 10963 13857 10993 13925
rect 11059 13857 11089 13925
rect 11225 13903 11255 13925
rect 12613 13959 12697 13975
rect 12613 13925 12623 13959
rect 12657 13925 12697 13959
rect 12613 13909 12697 13925
rect 12739 13959 12793 13975
rect 12739 13925 12749 13959
rect 12783 13925 12793 13959
rect 12739 13909 12793 13925
rect 9749 13759 9779 13785
rect 11949 13849 11979 13875
rect 10769 13747 10799 13773
rect 10857 13747 10887 13773
rect 10963 13747 10993 13773
rect 11059 13747 11089 13773
rect 11225 13747 11255 13773
rect 11780 13733 11810 13759
rect 11852 13733 11882 13759
rect 12667 13847 12697 13909
rect 12763 13847 12793 13909
rect 12835 13892 12865 14007
rect 12931 13975 12961 14007
rect 13029 13975 13059 14007
rect 12915 13959 12969 13975
rect 12915 13925 12925 13959
rect 12959 13925 12969 13959
rect 12915 13909 12969 13925
rect 13011 13959 13066 13975
rect 13011 13925 13021 13959
rect 13055 13925 13066 13959
rect 13011 13909 13066 13925
rect 12835 13891 12876 13892
rect 12835 13862 12877 13891
rect 12847 13847 12877 13862
rect 12931 13847 12961 13909
rect 13029 13887 13059 13909
rect 12667 13737 12697 13763
rect 12763 13737 12793 13763
rect 12847 13737 12877 13763
rect 12931 13737 12961 13763
rect 13029 13731 13059 13757
rect 11780 13617 11810 13649
rect 11710 13601 11810 13617
rect 11710 13567 11726 13601
rect 11760 13567 11810 13601
rect 11710 13551 11810 13567
rect 11852 13617 11882 13649
rect 11949 13617 11979 13649
rect 11852 13601 11906 13617
rect 11852 13567 11862 13601
rect 11896 13567 11906 13601
rect 11852 13551 11906 13567
rect 11949 13601 12015 13617
rect 11949 13567 11965 13601
rect 11999 13567 12015 13601
rect 11949 13551 12015 13567
rect 11768 13483 11798 13551
rect 11852 13483 11882 13551
rect 11949 13529 11979 13551
rect 11165 13381 11195 13407
rect 10977 13360 11031 13376
rect 9423 13311 9453 13337
rect 9507 13311 9537 13337
rect 9591 13311 9621 13337
rect 9675 13311 9705 13337
rect 9863 13311 9893 13337
rect 10977 13326 10987 13360
rect 11021 13326 11031 13360
rect 10977 13310 11031 13326
rect 10893 13268 10923 13309
rect 10977 13268 11007 13310
rect 11070 13268 11100 13294
rect 10893 13135 10923 13184
rect 10977 13166 11007 13184
rect 9423 13079 9453 13111
rect 9507 13079 9537 13111
rect 9591 13079 9621 13111
rect 9675 13079 9705 13111
rect 9863 13079 9893 13111
rect 9411 13063 9465 13079
rect 9411 13029 9421 13063
rect 9455 13029 9465 13063
rect 9411 13013 9465 13029
rect 9507 13063 9621 13079
rect 9507 13029 9538 13063
rect 9572 13029 9621 13063
rect 9507 13013 9621 13029
rect 9663 13063 9717 13079
rect 9663 13029 9673 13063
rect 9707 13029 9717 13063
rect 9663 13013 9717 13029
rect 9759 13063 9893 13079
rect 9759 13029 9769 13063
rect 9803 13046 9893 13063
rect 10839 13087 10923 13135
rect 10839 13053 10849 13087
rect 10883 13053 10923 13087
rect 9803 13029 9889 13046
rect 10839 13030 10923 13053
rect 9759 13013 9889 13029
rect 10893 13015 10923 13030
rect 10965 13141 11007 13166
rect 11070 13143 11100 13184
rect 11768 13373 11798 13399
rect 11852 13373 11882 13399
rect 11949 13373 11979 13399
rect 11165 13149 11195 13181
rect 10965 13015 10995 13141
rect 11049 13127 11103 13143
rect 11049 13110 11059 13127
rect 11037 13093 11059 13110
rect 11093 13093 11103 13127
rect 11037 13077 11103 13093
rect 11145 13133 11199 13149
rect 11145 13099 11155 13133
rect 11189 13099 11199 13133
rect 11145 13083 11199 13099
rect 11037 13054 11079 13077
rect 11165 13061 11195 13083
rect 11037 13030 11074 13054
rect 11037 13015 11067 13030
rect 9423 12991 9453 13013
rect 9507 12991 9537 13013
rect 9591 12991 9621 13013
rect 9675 12991 9705 13013
rect 9859 12991 9889 13013
rect 10893 12905 10923 12931
rect 10965 12905 10995 12931
rect 11037 12905 11067 12931
rect 11165 12905 11195 12931
rect 9423 12835 9453 12861
rect 9507 12835 9537 12861
rect 9591 12835 9621 12861
rect 9675 12835 9705 12861
rect 9859 12835 9889 12861
rect 9741 12567 9771 12593
rect 9549 12525 9579 12551
rect 9633 12525 9663 12551
rect 9549 12335 9579 12441
rect 9492 12319 9579 12335
rect 9492 12285 9508 12319
rect 9542 12285 9579 12319
rect 9492 12269 9579 12285
rect 9549 12229 9579 12269
rect 9633 12335 9663 12441
rect 9741 12335 9771 12367
rect 11117 12361 11147 12387
rect 9633 12319 9699 12335
rect 9633 12285 9649 12319
rect 9683 12285 9699 12319
rect 9633 12269 9699 12285
rect 9741 12319 9807 12335
rect 10925 12319 10955 12345
rect 11009 12319 11039 12345
rect 9741 12285 9757 12319
rect 9791 12285 9807 12319
rect 9741 12269 9807 12285
rect 9633 12229 9663 12269
rect 9741 12247 9771 12269
rect 9549 12119 9579 12145
rect 9633 12119 9663 12145
rect 10925 12129 10955 12235
rect 9741 12091 9771 12117
rect 10868 12113 10955 12129
rect 10868 12079 10884 12113
rect 10918 12079 10955 12113
rect 10868 12063 10955 12079
rect 10925 12023 10955 12063
rect 11009 12129 11039 12235
rect 11117 12129 11147 12161
rect 11009 12113 11075 12129
rect 11009 12079 11025 12113
rect 11059 12079 11075 12113
rect 11009 12063 11075 12079
rect 11117 12113 11183 12129
rect 11117 12079 11133 12113
rect 11167 12079 11183 12113
rect 11117 12063 11183 12079
rect 11009 12023 11039 12063
rect 11117 12041 11147 12063
rect 10925 11913 10955 11939
rect 11009 11913 11039 11939
rect 11117 11885 11147 11911
rect 9433 11747 9463 11773
rect 9517 11747 9547 11773
rect 9601 11747 9631 11773
rect 9685 11747 9715 11773
rect 9873 11747 9903 11773
rect 9433 11515 9463 11547
rect 9517 11515 9547 11547
rect 9601 11515 9631 11547
rect 9685 11515 9715 11547
rect 9873 11515 9903 11547
rect 9421 11499 9475 11515
rect 9421 11465 9431 11499
rect 9465 11465 9475 11499
rect 9421 11449 9475 11465
rect 9517 11499 9631 11515
rect 9517 11465 9548 11499
rect 9582 11465 9631 11499
rect 9517 11449 9631 11465
rect 9673 11499 9727 11515
rect 9673 11465 9683 11499
rect 9717 11465 9727 11499
rect 9673 11449 9727 11465
rect 9769 11499 9903 11515
rect 9769 11465 9779 11499
rect 9813 11482 9903 11499
rect 9813 11465 9899 11482
rect 9769 11449 9899 11465
rect 9433 11427 9463 11449
rect 9517 11427 9547 11449
rect 9601 11427 9631 11449
rect 9685 11427 9715 11449
rect 9869 11427 9899 11449
rect 9433 11271 9463 11297
rect 9517 11271 9547 11297
rect 9601 11271 9631 11297
rect 9685 11271 9715 11297
rect 9869 11271 9899 11297
rect 9751 11003 9781 11029
rect 9559 10961 9589 10987
rect 9643 10961 9673 10987
rect 9559 10771 9589 10877
rect 9502 10755 9589 10771
rect 9502 10721 9518 10755
rect 9552 10721 9589 10755
rect 9502 10705 9589 10721
rect 9559 10665 9589 10705
rect 9643 10771 9673 10877
rect 9751 10771 9781 10803
rect 9643 10755 9709 10771
rect 9643 10721 9659 10755
rect 9693 10721 9709 10755
rect 9643 10705 9709 10721
rect 9751 10755 9817 10771
rect 9751 10721 9767 10755
rect 9801 10721 9817 10755
rect 9751 10705 9817 10721
rect 9643 10665 9673 10705
rect 9751 10683 9781 10705
rect 9559 10555 9589 10581
rect 9643 10555 9673 10581
rect 9751 10527 9781 10553
rect 6238 6553 6268 6579
rect 6238 6401 6268 6423
rect 6238 6385 6324 6401
rect 6238 6351 6274 6385
rect 6308 6351 6324 6385
rect 6238 6335 6324 6351
rect 6238 6303 6268 6335
rect 6238 6077 6268 6103
rect 10132 5921 10162 5947
rect 10231 5921 10261 5947
rect 10327 5921 10357 5947
rect 10399 5921 10429 5947
rect 10495 5921 10525 5947
rect 10584 5921 10614 5947
rect 10668 5921 10698 5947
rect 10752 5921 10782 5947
rect 10940 5921 10970 5947
rect 11024 5921 11054 5947
rect 11108 5921 11138 5947
rect 11192 5921 11222 5947
rect 11282 5921 11312 5947
rect 11381 5921 11411 5947
rect 10132 5769 10162 5791
rect 10231 5777 10261 5837
rect 10132 5753 10186 5769
rect 10132 5719 10142 5753
rect 10176 5719 10186 5753
rect 10132 5703 10186 5719
rect 10231 5761 10285 5777
rect 10231 5727 10241 5761
rect 10275 5727 10285 5761
rect 10231 5711 10285 5727
rect 10132 5671 10162 5703
rect 1950 5501 1980 5527
rect 2049 5501 2079 5527
rect 2145 5501 2175 5527
rect 2217 5501 2247 5527
rect 2313 5501 2343 5527
rect 2402 5501 2432 5527
rect 2486 5501 2516 5527
rect 2570 5501 2600 5527
rect 2758 5501 2788 5527
rect 2842 5501 2872 5527
rect 2926 5501 2956 5527
rect 3010 5501 3040 5527
rect 3100 5501 3130 5527
rect 3199 5501 3229 5527
rect 1950 5349 1980 5371
rect 2049 5357 2079 5417
rect 1950 5333 2004 5349
rect 1950 5299 1960 5333
rect 1994 5299 2004 5333
rect 1950 5283 2004 5299
rect 2049 5341 2103 5357
rect 2049 5307 2059 5341
rect 2093 5307 2103 5341
rect 2049 5291 2103 5307
rect 1950 5251 1980 5283
rect 2049 5135 2079 5291
rect 2145 5245 2175 5417
rect 2121 5229 2175 5245
rect 2121 5195 2131 5229
rect 2165 5195 2175 5229
rect 2121 5179 2175 5195
rect 2145 5135 2175 5179
rect 2217 5245 2247 5417
rect 2313 5373 2343 5417
rect 2402 5373 2432 5417
rect 2486 5402 2516 5417
rect 2289 5357 2343 5373
rect 2289 5323 2299 5357
rect 2333 5323 2343 5357
rect 2289 5307 2343 5323
rect 2389 5357 2443 5373
rect 2389 5323 2399 5357
rect 2433 5323 2443 5357
rect 2389 5307 2443 5323
rect 2485 5372 2516 5402
rect 2570 5402 2600 5417
rect 2758 5402 2788 5417
rect 2570 5372 2788 5402
rect 2217 5229 2271 5245
rect 2217 5195 2227 5229
rect 2261 5195 2271 5229
rect 2217 5179 2271 5195
rect 2217 5135 2247 5179
rect 2313 5135 2343 5307
rect 2402 5135 2432 5307
rect 2485 5261 2515 5372
rect 2570 5357 2611 5372
rect 2581 5261 2611 5357
rect 2842 5342 2872 5417
rect 2926 5343 2956 5417
rect 2818 5326 2872 5342
rect 2818 5292 2828 5326
rect 2862 5292 2872 5326
rect 2818 5276 2872 5292
rect 2914 5327 2968 5343
rect 2914 5293 2924 5327
rect 2958 5293 2968 5327
rect 2914 5277 2968 5293
rect 2474 5245 2528 5261
rect 2474 5211 2484 5245
rect 2518 5211 2528 5245
rect 2474 5195 2528 5211
rect 2581 5245 2645 5261
rect 2581 5211 2601 5245
rect 2635 5211 2645 5245
rect 2486 5135 2516 5195
rect 2581 5180 2645 5211
rect 2570 5150 2788 5180
rect 2570 5135 2600 5150
rect 2758 5135 2788 5150
rect 2842 5135 2872 5276
rect 2926 5135 2956 5277
rect 3010 5238 3040 5417
rect 3100 5349 3130 5417
rect 4084 5493 4114 5519
rect 4183 5493 4213 5519
rect 4279 5493 4309 5519
rect 4351 5493 4381 5519
rect 4447 5493 4477 5519
rect 4536 5493 4566 5519
rect 4620 5493 4650 5519
rect 4704 5493 4734 5519
rect 4892 5493 4922 5519
rect 4976 5493 5006 5519
rect 5060 5493 5090 5519
rect 5144 5493 5174 5519
rect 5234 5493 5264 5519
rect 5333 5493 5363 5519
rect 6036 5493 6066 5519
rect 6135 5493 6165 5519
rect 6231 5493 6261 5519
rect 6303 5493 6333 5519
rect 6399 5493 6429 5519
rect 6488 5493 6518 5519
rect 6572 5493 6602 5519
rect 6656 5493 6686 5519
rect 6844 5493 6874 5519
rect 6928 5493 6958 5519
rect 7012 5493 7042 5519
rect 7096 5493 7126 5519
rect 7186 5493 7216 5519
rect 7285 5493 7315 5519
rect 8038 5499 8068 5525
rect 8137 5499 8167 5525
rect 8233 5499 8263 5525
rect 8305 5499 8335 5525
rect 8401 5499 8431 5525
rect 8490 5499 8520 5525
rect 8574 5499 8604 5525
rect 8658 5499 8688 5525
rect 8846 5499 8876 5525
rect 8930 5499 8960 5525
rect 9014 5499 9044 5525
rect 9098 5499 9128 5525
rect 9188 5499 9218 5525
rect 9287 5499 9317 5525
rect 3199 5349 3229 5371
rect 3082 5333 3136 5349
rect 3082 5299 3092 5333
rect 3126 5299 3136 5333
rect 3082 5283 3136 5299
rect 3178 5333 3232 5349
rect 3178 5299 3188 5333
rect 3222 5299 3232 5333
rect 3178 5283 3232 5299
rect 4084 5341 4114 5363
rect 4183 5349 4213 5409
rect 4084 5325 4138 5341
rect 4084 5291 4094 5325
rect 4128 5291 4138 5325
rect 3004 5222 3058 5238
rect 3004 5188 3014 5222
rect 3048 5188 3058 5222
rect 3004 5172 3058 5188
rect 3010 5135 3040 5172
rect 3100 5135 3130 5283
rect 3199 5251 3229 5283
rect 4084 5275 4138 5291
rect 4183 5333 4237 5349
rect 4183 5299 4193 5333
rect 4227 5299 4237 5333
rect 4183 5283 4237 5299
rect 4084 5243 4114 5275
rect 1950 5025 1980 5051
rect 2049 5025 2079 5051
rect 2145 5025 2175 5051
rect 2217 5025 2247 5051
rect 2313 5025 2343 5051
rect 2402 5025 2432 5051
rect 2486 5025 2516 5051
rect 2570 5025 2600 5051
rect 2758 5025 2788 5051
rect 2842 5025 2872 5051
rect 2926 5025 2956 5051
rect 3010 5025 3040 5051
rect 3100 5025 3130 5051
rect 3199 5025 3229 5051
rect 4183 5127 4213 5283
rect 4279 5237 4309 5409
rect 4255 5221 4309 5237
rect 4255 5187 4265 5221
rect 4299 5187 4309 5221
rect 4255 5171 4309 5187
rect 4279 5127 4309 5171
rect 4351 5237 4381 5409
rect 4447 5365 4477 5409
rect 4536 5365 4566 5409
rect 4620 5394 4650 5409
rect 4423 5349 4477 5365
rect 4423 5315 4433 5349
rect 4467 5315 4477 5349
rect 4423 5299 4477 5315
rect 4523 5349 4577 5365
rect 4523 5315 4533 5349
rect 4567 5315 4577 5349
rect 4523 5299 4577 5315
rect 4619 5364 4650 5394
rect 4704 5394 4734 5409
rect 4892 5394 4922 5409
rect 4704 5364 4922 5394
rect 4351 5221 4405 5237
rect 4351 5187 4361 5221
rect 4395 5187 4405 5221
rect 4351 5171 4405 5187
rect 4351 5127 4381 5171
rect 4447 5127 4477 5299
rect 4536 5127 4566 5299
rect 4619 5253 4649 5364
rect 4704 5349 4745 5364
rect 4715 5253 4745 5349
rect 4976 5334 5006 5409
rect 5060 5335 5090 5409
rect 4952 5318 5006 5334
rect 4952 5284 4962 5318
rect 4996 5284 5006 5318
rect 4952 5268 5006 5284
rect 5048 5319 5102 5335
rect 5048 5285 5058 5319
rect 5092 5285 5102 5319
rect 5048 5269 5102 5285
rect 4608 5237 4662 5253
rect 4608 5203 4618 5237
rect 4652 5203 4662 5237
rect 4608 5187 4662 5203
rect 4715 5237 4779 5253
rect 4715 5203 4735 5237
rect 4769 5203 4779 5237
rect 4620 5127 4650 5187
rect 4715 5172 4779 5203
rect 4704 5142 4922 5172
rect 4704 5127 4734 5142
rect 4892 5127 4922 5142
rect 4976 5127 5006 5268
rect 5060 5127 5090 5269
rect 5144 5230 5174 5409
rect 5234 5341 5264 5409
rect 5333 5341 5363 5363
rect 6036 5341 6066 5363
rect 6135 5349 6165 5409
rect 5216 5325 5270 5341
rect 5216 5291 5226 5325
rect 5260 5291 5270 5325
rect 5216 5275 5270 5291
rect 5312 5325 5366 5341
rect 5312 5291 5322 5325
rect 5356 5291 5366 5325
rect 5312 5275 5366 5291
rect 6036 5325 6090 5341
rect 6036 5291 6046 5325
rect 6080 5291 6090 5325
rect 6036 5275 6090 5291
rect 6135 5333 6189 5349
rect 6135 5299 6145 5333
rect 6179 5299 6189 5333
rect 6135 5283 6189 5299
rect 5138 5214 5192 5230
rect 5138 5180 5148 5214
rect 5182 5180 5192 5214
rect 5138 5164 5192 5180
rect 5144 5127 5174 5164
rect 5234 5127 5264 5275
rect 5333 5243 5363 5275
rect 6036 5243 6066 5275
rect 6135 5127 6165 5283
rect 6231 5237 6261 5409
rect 6207 5221 6261 5237
rect 6207 5187 6217 5221
rect 6251 5187 6261 5221
rect 6207 5171 6261 5187
rect 6231 5127 6261 5171
rect 6303 5237 6333 5409
rect 6399 5365 6429 5409
rect 6488 5365 6518 5409
rect 6572 5394 6602 5409
rect 6375 5349 6429 5365
rect 6375 5315 6385 5349
rect 6419 5315 6429 5349
rect 6375 5299 6429 5315
rect 6475 5349 6529 5365
rect 6475 5315 6485 5349
rect 6519 5315 6529 5349
rect 6475 5299 6529 5315
rect 6571 5364 6602 5394
rect 6656 5394 6686 5409
rect 6844 5394 6874 5409
rect 6656 5364 6874 5394
rect 6303 5221 6357 5237
rect 6303 5187 6313 5221
rect 6347 5187 6357 5221
rect 6303 5171 6357 5187
rect 6303 5127 6333 5171
rect 6399 5127 6429 5299
rect 6488 5127 6518 5299
rect 6571 5253 6601 5364
rect 6656 5349 6697 5364
rect 6667 5253 6697 5349
rect 6928 5334 6958 5409
rect 7012 5335 7042 5409
rect 6904 5318 6958 5334
rect 6904 5284 6914 5318
rect 6948 5284 6958 5318
rect 6904 5268 6958 5284
rect 7000 5319 7054 5335
rect 7000 5285 7010 5319
rect 7044 5285 7054 5319
rect 7000 5269 7054 5285
rect 6560 5237 6614 5253
rect 6560 5203 6570 5237
rect 6604 5203 6614 5237
rect 6560 5187 6614 5203
rect 6667 5237 6731 5253
rect 6667 5203 6687 5237
rect 6721 5203 6731 5237
rect 6572 5127 6602 5187
rect 6667 5172 6731 5203
rect 6656 5142 6874 5172
rect 6656 5127 6686 5142
rect 6844 5127 6874 5142
rect 6928 5127 6958 5268
rect 7012 5127 7042 5269
rect 7096 5230 7126 5409
rect 7186 5341 7216 5409
rect 7285 5341 7315 5363
rect 8038 5347 8068 5369
rect 8137 5355 8167 5415
rect 7168 5325 7222 5341
rect 7168 5291 7178 5325
rect 7212 5291 7222 5325
rect 7168 5275 7222 5291
rect 7264 5325 7318 5341
rect 7264 5291 7274 5325
rect 7308 5291 7318 5325
rect 7264 5275 7318 5291
rect 8038 5331 8092 5347
rect 8038 5297 8048 5331
rect 8082 5297 8092 5331
rect 8038 5281 8092 5297
rect 8137 5339 8191 5355
rect 8137 5305 8147 5339
rect 8181 5305 8191 5339
rect 8137 5289 8191 5305
rect 7090 5214 7144 5230
rect 7090 5180 7100 5214
rect 7134 5180 7144 5214
rect 7090 5164 7144 5180
rect 7096 5127 7126 5164
rect 7186 5127 7216 5275
rect 7285 5243 7315 5275
rect 8038 5249 8068 5281
rect 8137 5133 8167 5289
rect 8233 5243 8263 5415
rect 8209 5227 8263 5243
rect 8209 5193 8219 5227
rect 8253 5193 8263 5227
rect 8209 5177 8263 5193
rect 8233 5133 8263 5177
rect 8305 5243 8335 5415
rect 8401 5371 8431 5415
rect 8490 5371 8520 5415
rect 8574 5400 8604 5415
rect 8377 5355 8431 5371
rect 8377 5321 8387 5355
rect 8421 5321 8431 5355
rect 8377 5305 8431 5321
rect 8477 5355 8531 5371
rect 8477 5321 8487 5355
rect 8521 5321 8531 5355
rect 8477 5305 8531 5321
rect 8573 5370 8604 5400
rect 8658 5400 8688 5415
rect 8846 5400 8876 5415
rect 8658 5370 8876 5400
rect 8305 5227 8359 5243
rect 8305 5193 8315 5227
rect 8349 5193 8359 5227
rect 8305 5177 8359 5193
rect 8305 5133 8335 5177
rect 8401 5133 8431 5305
rect 8490 5133 8520 5305
rect 8573 5259 8603 5370
rect 8658 5355 8699 5370
rect 8669 5259 8699 5355
rect 8930 5340 8960 5415
rect 9014 5341 9044 5415
rect 8906 5324 8960 5340
rect 8906 5290 8916 5324
rect 8950 5290 8960 5324
rect 8906 5274 8960 5290
rect 9002 5325 9056 5341
rect 9002 5291 9012 5325
rect 9046 5291 9056 5325
rect 9002 5275 9056 5291
rect 8562 5243 8616 5259
rect 8562 5209 8572 5243
rect 8606 5209 8616 5243
rect 8562 5193 8616 5209
rect 8669 5243 8733 5259
rect 8669 5209 8689 5243
rect 8723 5209 8733 5243
rect 8574 5133 8604 5193
rect 8669 5178 8733 5209
rect 8658 5148 8876 5178
rect 8658 5133 8688 5148
rect 8846 5133 8876 5148
rect 8930 5133 8960 5274
rect 9014 5133 9044 5275
rect 9098 5236 9128 5415
rect 9188 5347 9218 5415
rect 10231 5555 10261 5711
rect 10327 5665 10357 5837
rect 10303 5649 10357 5665
rect 10303 5615 10313 5649
rect 10347 5615 10357 5649
rect 10303 5599 10357 5615
rect 10327 5555 10357 5599
rect 10399 5665 10429 5837
rect 10495 5793 10525 5837
rect 10584 5793 10614 5837
rect 10668 5822 10698 5837
rect 10471 5777 10525 5793
rect 10471 5743 10481 5777
rect 10515 5743 10525 5777
rect 10471 5727 10525 5743
rect 10571 5777 10625 5793
rect 10571 5743 10581 5777
rect 10615 5743 10625 5777
rect 10571 5727 10625 5743
rect 10667 5792 10698 5822
rect 10752 5822 10782 5837
rect 10940 5822 10970 5837
rect 10752 5792 10970 5822
rect 10399 5649 10453 5665
rect 10399 5615 10409 5649
rect 10443 5615 10453 5649
rect 10399 5599 10453 5615
rect 10399 5555 10429 5599
rect 10495 5555 10525 5727
rect 10584 5555 10614 5727
rect 10667 5681 10697 5792
rect 10752 5777 10793 5792
rect 10763 5681 10793 5777
rect 11024 5762 11054 5837
rect 11108 5763 11138 5837
rect 11000 5746 11054 5762
rect 11000 5712 11010 5746
rect 11044 5712 11054 5746
rect 11000 5696 11054 5712
rect 11096 5747 11150 5763
rect 11096 5713 11106 5747
rect 11140 5713 11150 5747
rect 11096 5697 11150 5713
rect 10656 5665 10710 5681
rect 10656 5631 10666 5665
rect 10700 5631 10710 5665
rect 10656 5615 10710 5631
rect 10763 5665 10827 5681
rect 10763 5631 10783 5665
rect 10817 5631 10827 5665
rect 10668 5555 10698 5615
rect 10763 5600 10827 5631
rect 10752 5570 10970 5600
rect 10752 5555 10782 5570
rect 10940 5555 10970 5570
rect 11024 5555 11054 5696
rect 11108 5555 11138 5697
rect 11192 5658 11222 5837
rect 11282 5769 11312 5837
rect 12194 5909 12224 5935
rect 12293 5909 12323 5935
rect 12389 5909 12419 5935
rect 12461 5909 12491 5935
rect 12557 5909 12587 5935
rect 12646 5909 12676 5935
rect 12730 5909 12760 5935
rect 12814 5909 12844 5935
rect 13002 5909 13032 5935
rect 13086 5909 13116 5935
rect 13170 5909 13200 5935
rect 13254 5909 13284 5935
rect 13344 5909 13374 5935
rect 13443 5909 13473 5935
rect 14152 5917 14182 5943
rect 14251 5917 14281 5943
rect 14347 5917 14377 5943
rect 14419 5917 14449 5943
rect 14515 5917 14545 5943
rect 14604 5917 14634 5943
rect 14688 5917 14718 5943
rect 14772 5917 14802 5943
rect 14960 5917 14990 5943
rect 15044 5917 15074 5943
rect 15128 5917 15158 5943
rect 15212 5917 15242 5943
rect 15302 5917 15332 5943
rect 15401 5917 15431 5943
rect 16146 5923 16176 5949
rect 16245 5923 16275 5949
rect 16341 5923 16371 5949
rect 16413 5923 16443 5949
rect 16509 5923 16539 5949
rect 16598 5923 16628 5949
rect 16682 5923 16712 5949
rect 16766 5923 16796 5949
rect 16954 5923 16984 5949
rect 17038 5923 17068 5949
rect 17122 5923 17152 5949
rect 17206 5923 17236 5949
rect 17296 5923 17326 5949
rect 17395 5923 17425 5949
rect 11381 5769 11411 5791
rect 11264 5753 11318 5769
rect 11264 5719 11274 5753
rect 11308 5719 11318 5753
rect 11264 5703 11318 5719
rect 11360 5753 11414 5769
rect 11360 5719 11370 5753
rect 11404 5719 11414 5753
rect 11360 5703 11414 5719
rect 12194 5757 12224 5779
rect 12293 5765 12323 5825
rect 12194 5741 12248 5757
rect 12194 5707 12204 5741
rect 12238 5707 12248 5741
rect 11186 5642 11240 5658
rect 11186 5608 11196 5642
rect 11230 5608 11240 5642
rect 11186 5592 11240 5608
rect 11192 5555 11222 5592
rect 11282 5555 11312 5703
rect 11381 5671 11411 5703
rect 12194 5691 12248 5707
rect 12293 5749 12347 5765
rect 12293 5715 12303 5749
rect 12337 5715 12347 5749
rect 12293 5699 12347 5715
rect 12194 5659 12224 5691
rect 10132 5445 10162 5471
rect 10231 5445 10261 5471
rect 10327 5445 10357 5471
rect 10399 5445 10429 5471
rect 10495 5445 10525 5471
rect 10584 5445 10614 5471
rect 10668 5445 10698 5471
rect 10752 5445 10782 5471
rect 10940 5445 10970 5471
rect 11024 5445 11054 5471
rect 11108 5445 11138 5471
rect 11192 5445 11222 5471
rect 11282 5445 11312 5471
rect 11381 5445 11411 5471
rect 12293 5543 12323 5699
rect 12389 5653 12419 5825
rect 12365 5637 12419 5653
rect 12365 5603 12375 5637
rect 12409 5603 12419 5637
rect 12365 5587 12419 5603
rect 12389 5543 12419 5587
rect 12461 5653 12491 5825
rect 12557 5781 12587 5825
rect 12646 5781 12676 5825
rect 12730 5810 12760 5825
rect 12533 5765 12587 5781
rect 12533 5731 12543 5765
rect 12577 5731 12587 5765
rect 12533 5715 12587 5731
rect 12633 5765 12687 5781
rect 12633 5731 12643 5765
rect 12677 5731 12687 5765
rect 12633 5715 12687 5731
rect 12729 5780 12760 5810
rect 12814 5810 12844 5825
rect 13002 5810 13032 5825
rect 12814 5780 13032 5810
rect 12461 5637 12515 5653
rect 12461 5603 12471 5637
rect 12505 5603 12515 5637
rect 12461 5587 12515 5603
rect 12461 5543 12491 5587
rect 12557 5543 12587 5715
rect 12646 5543 12676 5715
rect 12729 5669 12759 5780
rect 12814 5765 12855 5780
rect 12825 5669 12855 5765
rect 13086 5750 13116 5825
rect 13170 5751 13200 5825
rect 13062 5734 13116 5750
rect 13062 5700 13072 5734
rect 13106 5700 13116 5734
rect 13062 5684 13116 5700
rect 13158 5735 13212 5751
rect 13158 5701 13168 5735
rect 13202 5701 13212 5735
rect 13158 5685 13212 5701
rect 12718 5653 12772 5669
rect 12718 5619 12728 5653
rect 12762 5619 12772 5653
rect 12718 5603 12772 5619
rect 12825 5653 12889 5669
rect 12825 5619 12845 5653
rect 12879 5619 12889 5653
rect 12730 5543 12760 5603
rect 12825 5588 12889 5619
rect 12814 5558 13032 5588
rect 12814 5543 12844 5558
rect 13002 5543 13032 5558
rect 13086 5543 13116 5684
rect 13170 5543 13200 5685
rect 13254 5646 13284 5825
rect 13344 5757 13374 5825
rect 13443 5757 13473 5779
rect 14152 5765 14182 5787
rect 14251 5773 14281 5833
rect 13326 5741 13380 5757
rect 13326 5707 13336 5741
rect 13370 5707 13380 5741
rect 13326 5691 13380 5707
rect 13422 5741 13476 5757
rect 13422 5707 13432 5741
rect 13466 5707 13476 5741
rect 13422 5691 13476 5707
rect 14152 5749 14206 5765
rect 14152 5715 14162 5749
rect 14196 5715 14206 5749
rect 14152 5699 14206 5715
rect 14251 5757 14305 5773
rect 14251 5723 14261 5757
rect 14295 5723 14305 5757
rect 14251 5707 14305 5723
rect 13248 5630 13302 5646
rect 13248 5596 13258 5630
rect 13292 5596 13302 5630
rect 13248 5580 13302 5596
rect 13254 5543 13284 5580
rect 13344 5543 13374 5691
rect 13443 5659 13473 5691
rect 14152 5667 14182 5699
rect 14251 5551 14281 5707
rect 14347 5661 14377 5833
rect 14323 5645 14377 5661
rect 14323 5611 14333 5645
rect 14367 5611 14377 5645
rect 14323 5595 14377 5611
rect 14347 5551 14377 5595
rect 14419 5661 14449 5833
rect 14515 5789 14545 5833
rect 14604 5789 14634 5833
rect 14688 5818 14718 5833
rect 14491 5773 14545 5789
rect 14491 5739 14501 5773
rect 14535 5739 14545 5773
rect 14491 5723 14545 5739
rect 14591 5773 14645 5789
rect 14591 5739 14601 5773
rect 14635 5739 14645 5773
rect 14591 5723 14645 5739
rect 14687 5788 14718 5818
rect 14772 5818 14802 5833
rect 14960 5818 14990 5833
rect 14772 5788 14990 5818
rect 14419 5645 14473 5661
rect 14419 5611 14429 5645
rect 14463 5611 14473 5645
rect 14419 5595 14473 5611
rect 14419 5551 14449 5595
rect 14515 5551 14545 5723
rect 14604 5551 14634 5723
rect 14687 5677 14717 5788
rect 14772 5773 14813 5788
rect 14783 5677 14813 5773
rect 15044 5758 15074 5833
rect 15128 5759 15158 5833
rect 15020 5742 15074 5758
rect 15020 5708 15030 5742
rect 15064 5708 15074 5742
rect 15020 5692 15074 5708
rect 15116 5743 15170 5759
rect 15116 5709 15126 5743
rect 15160 5709 15170 5743
rect 15116 5693 15170 5709
rect 14676 5661 14730 5677
rect 14676 5627 14686 5661
rect 14720 5627 14730 5661
rect 14676 5611 14730 5627
rect 14783 5661 14847 5677
rect 14783 5627 14803 5661
rect 14837 5627 14847 5661
rect 14688 5551 14718 5611
rect 14783 5596 14847 5627
rect 14772 5566 14990 5596
rect 14772 5551 14802 5566
rect 14960 5551 14990 5566
rect 15044 5551 15074 5692
rect 15128 5551 15158 5693
rect 15212 5654 15242 5833
rect 15302 5765 15332 5833
rect 15401 5765 15431 5787
rect 16146 5771 16176 5793
rect 16245 5779 16275 5839
rect 15284 5749 15338 5765
rect 15284 5715 15294 5749
rect 15328 5715 15338 5749
rect 15284 5699 15338 5715
rect 15380 5749 15434 5765
rect 15380 5715 15390 5749
rect 15424 5715 15434 5749
rect 15380 5699 15434 5715
rect 16146 5755 16200 5771
rect 16146 5721 16156 5755
rect 16190 5721 16200 5755
rect 16146 5705 16200 5721
rect 16245 5763 16299 5779
rect 16245 5729 16255 5763
rect 16289 5729 16299 5763
rect 16245 5713 16299 5729
rect 15206 5638 15260 5654
rect 15206 5604 15216 5638
rect 15250 5604 15260 5638
rect 15206 5588 15260 5604
rect 15212 5551 15242 5588
rect 15302 5551 15332 5699
rect 15401 5667 15431 5699
rect 16146 5673 16176 5705
rect 16245 5557 16275 5713
rect 16341 5667 16371 5839
rect 16317 5651 16371 5667
rect 16317 5617 16327 5651
rect 16361 5617 16371 5651
rect 16317 5601 16371 5617
rect 16341 5557 16371 5601
rect 16413 5667 16443 5839
rect 16509 5795 16539 5839
rect 16598 5795 16628 5839
rect 16682 5824 16712 5839
rect 16485 5779 16539 5795
rect 16485 5745 16495 5779
rect 16529 5745 16539 5779
rect 16485 5729 16539 5745
rect 16585 5779 16639 5795
rect 16585 5745 16595 5779
rect 16629 5745 16639 5779
rect 16585 5729 16639 5745
rect 16681 5794 16712 5824
rect 16766 5824 16796 5839
rect 16954 5824 16984 5839
rect 16766 5794 16984 5824
rect 16413 5651 16467 5667
rect 16413 5617 16423 5651
rect 16457 5617 16467 5651
rect 16413 5601 16467 5617
rect 16413 5557 16443 5601
rect 16509 5557 16539 5729
rect 16598 5557 16628 5729
rect 16681 5683 16711 5794
rect 16766 5779 16807 5794
rect 16777 5683 16807 5779
rect 17038 5764 17068 5839
rect 17122 5765 17152 5839
rect 17014 5748 17068 5764
rect 17014 5714 17024 5748
rect 17058 5714 17068 5748
rect 17014 5698 17068 5714
rect 17110 5749 17164 5765
rect 17110 5715 17120 5749
rect 17154 5715 17164 5749
rect 17110 5699 17164 5715
rect 16670 5667 16724 5683
rect 16670 5633 16680 5667
rect 16714 5633 16724 5667
rect 16670 5617 16724 5633
rect 16777 5667 16841 5683
rect 16777 5633 16797 5667
rect 16831 5633 16841 5667
rect 16682 5557 16712 5617
rect 16777 5602 16841 5633
rect 16766 5572 16984 5602
rect 16766 5557 16796 5572
rect 16954 5557 16984 5572
rect 17038 5557 17068 5698
rect 17122 5557 17152 5699
rect 17206 5660 17236 5839
rect 17296 5771 17326 5839
rect 17395 5771 17425 5793
rect 17278 5755 17332 5771
rect 17278 5721 17288 5755
rect 17322 5721 17332 5755
rect 17278 5705 17332 5721
rect 17374 5755 17428 5771
rect 17374 5721 17384 5755
rect 17418 5721 17428 5755
rect 17374 5705 17428 5721
rect 17200 5644 17254 5660
rect 17200 5610 17210 5644
rect 17244 5610 17254 5644
rect 17200 5594 17254 5610
rect 17206 5557 17236 5594
rect 17296 5557 17326 5705
rect 17395 5673 17425 5705
rect 12194 5433 12224 5459
rect 12293 5433 12323 5459
rect 12389 5433 12419 5459
rect 12461 5433 12491 5459
rect 12557 5433 12587 5459
rect 12646 5433 12676 5459
rect 12730 5433 12760 5459
rect 12814 5433 12844 5459
rect 13002 5433 13032 5459
rect 13086 5433 13116 5459
rect 13170 5433 13200 5459
rect 13254 5433 13284 5459
rect 13344 5433 13374 5459
rect 13443 5433 13473 5459
rect 14152 5441 14182 5467
rect 14251 5441 14281 5467
rect 14347 5441 14377 5467
rect 14419 5441 14449 5467
rect 14515 5441 14545 5467
rect 14604 5441 14634 5467
rect 14688 5441 14718 5467
rect 14772 5441 14802 5467
rect 14960 5441 14990 5467
rect 15044 5441 15074 5467
rect 15128 5441 15158 5467
rect 15212 5441 15242 5467
rect 15302 5441 15332 5467
rect 15401 5441 15431 5467
rect 16146 5447 16176 5473
rect 16245 5447 16275 5473
rect 16341 5447 16371 5473
rect 16413 5447 16443 5473
rect 16509 5447 16539 5473
rect 16598 5447 16628 5473
rect 16682 5447 16712 5473
rect 16766 5447 16796 5473
rect 16954 5447 16984 5473
rect 17038 5447 17068 5473
rect 17122 5447 17152 5473
rect 17206 5447 17236 5473
rect 17296 5447 17326 5473
rect 17395 5447 17425 5473
rect 9287 5347 9317 5369
rect 9170 5331 9224 5347
rect 9170 5297 9180 5331
rect 9214 5297 9224 5331
rect 9170 5281 9224 5297
rect 9266 5331 9320 5347
rect 9266 5297 9276 5331
rect 9310 5297 9320 5331
rect 9266 5281 9320 5297
rect 9092 5220 9146 5236
rect 9092 5186 9102 5220
rect 9136 5186 9146 5220
rect 9092 5170 9146 5186
rect 9098 5133 9128 5170
rect 9188 5133 9218 5281
rect 9287 5249 9317 5281
rect 4084 5017 4114 5043
rect 4183 5017 4213 5043
rect 4279 5017 4309 5043
rect 4351 5017 4381 5043
rect 4447 5017 4477 5043
rect 4536 5017 4566 5043
rect 4620 5017 4650 5043
rect 4704 5017 4734 5043
rect 4892 5017 4922 5043
rect 4976 5017 5006 5043
rect 5060 5017 5090 5043
rect 5144 5017 5174 5043
rect 5234 5017 5264 5043
rect 5333 5017 5363 5043
rect 6036 5017 6066 5043
rect 6135 5017 6165 5043
rect 6231 5017 6261 5043
rect 6303 5017 6333 5043
rect 6399 5017 6429 5043
rect 6488 5017 6518 5043
rect 6572 5017 6602 5043
rect 6656 5017 6686 5043
rect 6844 5017 6874 5043
rect 6928 5017 6958 5043
rect 7012 5017 7042 5043
rect 7096 5017 7126 5043
rect 7186 5017 7216 5043
rect 7285 5017 7315 5043
rect 8038 5023 8068 5049
rect 8137 5023 8167 5049
rect 8233 5023 8263 5049
rect 8305 5023 8335 5049
rect 8401 5023 8431 5049
rect 8490 5023 8520 5049
rect 8574 5023 8604 5049
rect 8658 5023 8688 5049
rect 8846 5023 8876 5049
rect 8930 5023 8960 5049
rect 9014 5023 9044 5049
rect 9098 5023 9128 5049
rect 9188 5023 9218 5049
rect 9287 5023 9317 5049
rect 10160 5047 10190 5073
rect 10259 5047 10289 5073
rect 10355 5047 10385 5073
rect 10427 5047 10457 5073
rect 10523 5047 10553 5073
rect 10612 5047 10642 5073
rect 10696 5047 10726 5073
rect 10780 5047 10810 5073
rect 10968 5047 10998 5073
rect 11052 5047 11082 5073
rect 11136 5047 11166 5073
rect 11220 5047 11250 5073
rect 11310 5047 11340 5073
rect 11409 5047 11439 5073
rect 10160 4895 10190 4917
rect 10259 4903 10289 4963
rect 10160 4879 10214 4895
rect 10160 4845 10170 4879
rect 10204 4845 10214 4879
rect 10160 4829 10214 4845
rect 10259 4887 10313 4903
rect 10259 4853 10269 4887
rect 10303 4853 10313 4887
rect 10259 4837 10313 4853
rect 10160 4797 10190 4829
rect 10259 4681 10289 4837
rect 10355 4791 10385 4963
rect 10331 4775 10385 4791
rect 10331 4741 10341 4775
rect 10375 4741 10385 4775
rect 10331 4725 10385 4741
rect 10355 4681 10385 4725
rect 10427 4791 10457 4963
rect 10523 4919 10553 4963
rect 10612 4919 10642 4963
rect 10696 4948 10726 4963
rect 10499 4903 10553 4919
rect 10499 4869 10509 4903
rect 10543 4869 10553 4903
rect 10499 4853 10553 4869
rect 10599 4903 10653 4919
rect 10599 4869 10609 4903
rect 10643 4869 10653 4903
rect 10599 4853 10653 4869
rect 10695 4918 10726 4948
rect 10780 4948 10810 4963
rect 10968 4948 10998 4963
rect 10780 4918 10998 4948
rect 10427 4775 10481 4791
rect 10427 4741 10437 4775
rect 10471 4741 10481 4775
rect 10427 4725 10481 4741
rect 10427 4681 10457 4725
rect 10523 4681 10553 4853
rect 10612 4681 10642 4853
rect 10695 4807 10725 4918
rect 10780 4903 10821 4918
rect 10791 4807 10821 4903
rect 11052 4888 11082 4963
rect 11136 4889 11166 4963
rect 11028 4872 11082 4888
rect 11028 4838 11038 4872
rect 11072 4838 11082 4872
rect 11028 4822 11082 4838
rect 11124 4873 11178 4889
rect 11124 4839 11134 4873
rect 11168 4839 11178 4873
rect 11124 4823 11178 4839
rect 10684 4791 10738 4807
rect 10684 4757 10694 4791
rect 10728 4757 10738 4791
rect 10684 4741 10738 4757
rect 10791 4791 10855 4807
rect 10791 4757 10811 4791
rect 10845 4757 10855 4791
rect 10696 4681 10726 4741
rect 10791 4726 10855 4757
rect 10780 4696 10998 4726
rect 10780 4681 10810 4696
rect 10968 4681 10998 4696
rect 11052 4681 11082 4822
rect 11136 4681 11166 4823
rect 11220 4784 11250 4963
rect 11310 4895 11340 4963
rect 12430 5003 12460 5029
rect 12529 5003 12559 5029
rect 12625 5003 12655 5029
rect 12697 5003 12727 5029
rect 12793 5003 12823 5029
rect 12882 5003 12912 5029
rect 12966 5003 12996 5029
rect 13050 5003 13080 5029
rect 13238 5003 13268 5029
rect 13322 5003 13352 5029
rect 13406 5003 13436 5029
rect 13490 5003 13520 5029
rect 13580 5003 13610 5029
rect 13679 5003 13709 5029
rect 11409 4895 11439 4917
rect 11292 4879 11346 4895
rect 11292 4845 11302 4879
rect 11336 4845 11346 4879
rect 11292 4829 11346 4845
rect 11388 4879 11442 4895
rect 11388 4845 11398 4879
rect 11432 4845 11442 4879
rect 11388 4829 11442 4845
rect 12430 4851 12460 4873
rect 12529 4859 12559 4919
rect 12430 4835 12484 4851
rect 11214 4768 11268 4784
rect 11214 4734 11224 4768
rect 11258 4734 11268 4768
rect 11214 4718 11268 4734
rect 11220 4681 11250 4718
rect 11310 4681 11340 4829
rect 11409 4797 11439 4829
rect 12430 4801 12440 4835
rect 12474 4801 12484 4835
rect 12430 4785 12484 4801
rect 12529 4843 12583 4859
rect 12529 4809 12539 4843
rect 12573 4809 12583 4843
rect 12529 4793 12583 4809
rect 12430 4753 12460 4785
rect 10160 4571 10190 4597
rect 10259 4571 10289 4597
rect 10355 4571 10385 4597
rect 10427 4571 10457 4597
rect 10523 4571 10553 4597
rect 10612 4571 10642 4597
rect 10696 4571 10726 4597
rect 10780 4571 10810 4597
rect 10968 4571 10998 4597
rect 11052 4571 11082 4597
rect 11136 4571 11166 4597
rect 11220 4571 11250 4597
rect 11310 4571 11340 4597
rect 11409 4571 11439 4597
rect 12529 4637 12559 4793
rect 12625 4747 12655 4919
rect 12601 4731 12655 4747
rect 12601 4697 12611 4731
rect 12645 4697 12655 4731
rect 12601 4681 12655 4697
rect 12625 4637 12655 4681
rect 12697 4747 12727 4919
rect 12793 4875 12823 4919
rect 12882 4875 12912 4919
rect 12966 4904 12996 4919
rect 12769 4859 12823 4875
rect 12769 4825 12779 4859
rect 12813 4825 12823 4859
rect 12769 4809 12823 4825
rect 12869 4859 12923 4875
rect 12869 4825 12879 4859
rect 12913 4825 12923 4859
rect 12869 4809 12923 4825
rect 12965 4874 12996 4904
rect 13050 4904 13080 4919
rect 13238 4904 13268 4919
rect 13050 4874 13268 4904
rect 12697 4731 12751 4747
rect 12697 4697 12707 4731
rect 12741 4697 12751 4731
rect 12697 4681 12751 4697
rect 12697 4637 12727 4681
rect 12793 4637 12823 4809
rect 12882 4637 12912 4809
rect 12965 4763 12995 4874
rect 13050 4859 13091 4874
rect 13061 4763 13091 4859
rect 13322 4844 13352 4919
rect 13406 4845 13436 4919
rect 13298 4828 13352 4844
rect 13298 4794 13308 4828
rect 13342 4794 13352 4828
rect 13298 4778 13352 4794
rect 13394 4829 13448 4845
rect 13394 4795 13404 4829
rect 13438 4795 13448 4829
rect 13394 4779 13448 4795
rect 12954 4747 13008 4763
rect 12954 4713 12964 4747
rect 12998 4713 13008 4747
rect 12954 4697 13008 4713
rect 13061 4747 13125 4763
rect 13061 4713 13081 4747
rect 13115 4713 13125 4747
rect 12966 4637 12996 4697
rect 13061 4682 13125 4713
rect 13050 4652 13268 4682
rect 13050 4637 13080 4652
rect 13238 4637 13268 4652
rect 13322 4637 13352 4778
rect 13406 4637 13436 4779
rect 13490 4740 13520 4919
rect 13580 4851 13610 4919
rect 14432 4997 14462 5023
rect 14531 4997 14561 5023
rect 14627 4997 14657 5023
rect 14699 4997 14729 5023
rect 14795 4997 14825 5023
rect 14884 4997 14914 5023
rect 14968 4997 14998 5023
rect 15052 4997 15082 5023
rect 15240 4997 15270 5023
rect 15324 4997 15354 5023
rect 15408 4997 15438 5023
rect 15492 4997 15522 5023
rect 15582 4997 15612 5023
rect 15681 4997 15711 5023
rect 13679 4851 13709 4873
rect 13562 4835 13616 4851
rect 13562 4801 13572 4835
rect 13606 4801 13616 4835
rect 13562 4785 13616 4801
rect 13658 4835 13712 4851
rect 13658 4801 13668 4835
rect 13702 4801 13712 4835
rect 13658 4785 13712 4801
rect 14432 4845 14462 4867
rect 14531 4853 14561 4913
rect 14432 4829 14486 4845
rect 14432 4795 14442 4829
rect 14476 4795 14486 4829
rect 13484 4724 13538 4740
rect 13484 4690 13494 4724
rect 13528 4690 13538 4724
rect 13484 4674 13538 4690
rect 13490 4637 13520 4674
rect 13580 4637 13610 4785
rect 13679 4753 13709 4785
rect 14432 4779 14486 4795
rect 14531 4837 14585 4853
rect 14531 4803 14541 4837
rect 14575 4803 14585 4837
rect 14531 4787 14585 4803
rect 14432 4747 14462 4779
rect 12430 4527 12460 4553
rect 12529 4527 12559 4553
rect 12625 4527 12655 4553
rect 12697 4527 12727 4553
rect 12793 4527 12823 4553
rect 12882 4527 12912 4553
rect 12966 4527 12996 4553
rect 13050 4527 13080 4553
rect 13238 4527 13268 4553
rect 13322 4527 13352 4553
rect 13406 4527 13436 4553
rect 13490 4527 13520 4553
rect 13580 4527 13610 4553
rect 13679 4527 13709 4553
rect 14531 4631 14561 4787
rect 14627 4741 14657 4913
rect 14603 4725 14657 4741
rect 14603 4691 14613 4725
rect 14647 4691 14657 4725
rect 14603 4675 14657 4691
rect 14627 4631 14657 4675
rect 14699 4741 14729 4913
rect 14795 4869 14825 4913
rect 14884 4869 14914 4913
rect 14968 4898 14998 4913
rect 14771 4853 14825 4869
rect 14771 4819 14781 4853
rect 14815 4819 14825 4853
rect 14771 4803 14825 4819
rect 14871 4853 14925 4869
rect 14871 4819 14881 4853
rect 14915 4819 14925 4853
rect 14871 4803 14925 4819
rect 14967 4868 14998 4898
rect 15052 4898 15082 4913
rect 15240 4898 15270 4913
rect 15052 4868 15270 4898
rect 14699 4725 14753 4741
rect 14699 4691 14709 4725
rect 14743 4691 14753 4725
rect 14699 4675 14753 4691
rect 14699 4631 14729 4675
rect 14795 4631 14825 4803
rect 14884 4631 14914 4803
rect 14967 4757 14997 4868
rect 15052 4853 15093 4868
rect 15063 4757 15093 4853
rect 15324 4838 15354 4913
rect 15408 4839 15438 4913
rect 15300 4822 15354 4838
rect 15300 4788 15310 4822
rect 15344 4788 15354 4822
rect 15300 4772 15354 4788
rect 15396 4823 15450 4839
rect 15396 4789 15406 4823
rect 15440 4789 15450 4823
rect 15396 4773 15450 4789
rect 14956 4741 15010 4757
rect 14956 4707 14966 4741
rect 15000 4707 15010 4741
rect 14956 4691 15010 4707
rect 15063 4741 15127 4757
rect 15063 4707 15083 4741
rect 15117 4707 15127 4741
rect 14968 4631 14998 4691
rect 15063 4676 15127 4707
rect 15052 4646 15270 4676
rect 15052 4631 15082 4646
rect 15240 4631 15270 4646
rect 15324 4631 15354 4772
rect 15408 4631 15438 4773
rect 15492 4734 15522 4913
rect 15582 4845 15612 4913
rect 16454 4979 16484 5005
rect 16553 4979 16583 5005
rect 16649 4979 16679 5005
rect 16721 4979 16751 5005
rect 16817 4979 16847 5005
rect 16906 4979 16936 5005
rect 16990 4979 17020 5005
rect 17074 4979 17104 5005
rect 17262 4979 17292 5005
rect 17346 4979 17376 5005
rect 17430 4979 17460 5005
rect 17514 4979 17544 5005
rect 17604 4979 17634 5005
rect 17703 4979 17733 5005
rect 15681 4845 15711 4867
rect 15564 4829 15618 4845
rect 15564 4795 15574 4829
rect 15608 4795 15618 4829
rect 15564 4779 15618 4795
rect 15660 4829 15714 4845
rect 15660 4795 15670 4829
rect 15704 4795 15714 4829
rect 15660 4779 15714 4795
rect 16454 4827 16484 4849
rect 16553 4835 16583 4895
rect 16454 4811 16508 4827
rect 15486 4718 15540 4734
rect 15486 4684 15496 4718
rect 15530 4684 15540 4718
rect 15486 4668 15540 4684
rect 15492 4631 15522 4668
rect 15582 4631 15612 4779
rect 15681 4747 15711 4779
rect 16454 4777 16464 4811
rect 16498 4777 16508 4811
rect 16454 4761 16508 4777
rect 16553 4819 16607 4835
rect 16553 4785 16563 4819
rect 16597 4785 16607 4819
rect 16553 4769 16607 4785
rect 16454 4729 16484 4761
rect 14432 4521 14462 4547
rect 14531 4521 14561 4547
rect 14627 4521 14657 4547
rect 14699 4521 14729 4547
rect 14795 4521 14825 4547
rect 14884 4521 14914 4547
rect 14968 4521 14998 4547
rect 15052 4521 15082 4547
rect 15240 4521 15270 4547
rect 15324 4521 15354 4547
rect 15408 4521 15438 4547
rect 15492 4521 15522 4547
rect 15582 4521 15612 4547
rect 15681 4521 15711 4547
rect 16553 4613 16583 4769
rect 16649 4723 16679 4895
rect 16625 4707 16679 4723
rect 16625 4673 16635 4707
rect 16669 4673 16679 4707
rect 16625 4657 16679 4673
rect 16649 4613 16679 4657
rect 16721 4723 16751 4895
rect 16817 4851 16847 4895
rect 16906 4851 16936 4895
rect 16990 4880 17020 4895
rect 16793 4835 16847 4851
rect 16793 4801 16803 4835
rect 16837 4801 16847 4835
rect 16793 4785 16847 4801
rect 16893 4835 16947 4851
rect 16893 4801 16903 4835
rect 16937 4801 16947 4835
rect 16893 4785 16947 4801
rect 16989 4850 17020 4880
rect 17074 4880 17104 4895
rect 17262 4880 17292 4895
rect 17074 4850 17292 4880
rect 16721 4707 16775 4723
rect 16721 4673 16731 4707
rect 16765 4673 16775 4707
rect 16721 4657 16775 4673
rect 16721 4613 16751 4657
rect 16817 4613 16847 4785
rect 16906 4613 16936 4785
rect 16989 4739 17019 4850
rect 17074 4835 17115 4850
rect 17085 4739 17115 4835
rect 17346 4820 17376 4895
rect 17430 4821 17460 4895
rect 17322 4804 17376 4820
rect 17322 4770 17332 4804
rect 17366 4770 17376 4804
rect 17322 4754 17376 4770
rect 17418 4805 17472 4821
rect 17418 4771 17428 4805
rect 17462 4771 17472 4805
rect 17418 4755 17472 4771
rect 16978 4723 17032 4739
rect 16978 4689 16988 4723
rect 17022 4689 17032 4723
rect 16978 4673 17032 4689
rect 17085 4723 17149 4739
rect 17085 4689 17105 4723
rect 17139 4689 17149 4723
rect 16990 4613 17020 4673
rect 17085 4658 17149 4689
rect 17074 4628 17292 4658
rect 17074 4613 17104 4628
rect 17262 4613 17292 4628
rect 17346 4613 17376 4754
rect 17430 4613 17460 4755
rect 17514 4716 17544 4895
rect 17604 4827 17634 4895
rect 17703 4827 17733 4849
rect 17586 4811 17640 4827
rect 17586 4777 17596 4811
rect 17630 4777 17640 4811
rect 17586 4761 17640 4777
rect 17682 4811 17736 4827
rect 17682 4777 17692 4811
rect 17726 4777 17736 4811
rect 17682 4761 17736 4777
rect 17508 4700 17562 4716
rect 17508 4666 17518 4700
rect 17552 4666 17562 4700
rect 17508 4650 17562 4666
rect 17514 4613 17544 4650
rect 17604 4613 17634 4761
rect 17703 4729 17733 4761
rect 16454 4503 16484 4529
rect 16553 4503 16583 4529
rect 16649 4503 16679 4529
rect 16721 4503 16751 4529
rect 16817 4503 16847 4529
rect 16906 4503 16936 4529
rect 16990 4503 17020 4529
rect 17074 4503 17104 4529
rect 17262 4503 17292 4529
rect 17346 4503 17376 4529
rect 17430 4503 17460 4529
rect 17514 4503 17544 4529
rect 17604 4503 17634 4529
rect 17703 4503 17733 4529
rect 1920 2241 1950 2267
rect 2019 2241 2049 2267
rect 2115 2241 2145 2267
rect 2187 2241 2217 2267
rect 2283 2241 2313 2267
rect 2372 2241 2402 2267
rect 2456 2241 2486 2267
rect 2540 2241 2570 2267
rect 2728 2241 2758 2267
rect 2812 2241 2842 2267
rect 2896 2241 2926 2267
rect 2980 2241 3010 2267
rect 3070 2241 3100 2267
rect 3169 2241 3199 2267
rect 1920 2089 1950 2111
rect 2019 2097 2049 2157
rect 1920 2073 1974 2089
rect 1920 2039 1930 2073
rect 1964 2039 1974 2073
rect 1920 2023 1974 2039
rect 2019 2081 2073 2097
rect 2019 2047 2029 2081
rect 2063 2047 2073 2081
rect 2019 2031 2073 2047
rect 1920 1991 1950 2023
rect 2019 1875 2049 2031
rect 2115 1985 2145 2157
rect 2091 1969 2145 1985
rect 2091 1935 2101 1969
rect 2135 1935 2145 1969
rect 2091 1919 2145 1935
rect 2115 1875 2145 1919
rect 2187 1985 2217 2157
rect 2283 2113 2313 2157
rect 2372 2113 2402 2157
rect 2456 2142 2486 2157
rect 2259 2097 2313 2113
rect 2259 2063 2269 2097
rect 2303 2063 2313 2097
rect 2259 2047 2313 2063
rect 2359 2097 2413 2113
rect 2359 2063 2369 2097
rect 2403 2063 2413 2097
rect 2359 2047 2413 2063
rect 2455 2112 2486 2142
rect 2540 2142 2570 2157
rect 2728 2142 2758 2157
rect 2540 2112 2758 2142
rect 2187 1969 2241 1985
rect 2187 1935 2197 1969
rect 2231 1935 2241 1969
rect 2187 1919 2241 1935
rect 2187 1875 2217 1919
rect 2283 1875 2313 2047
rect 2372 1875 2402 2047
rect 2455 2001 2485 2112
rect 2540 2097 2581 2112
rect 2551 2001 2581 2097
rect 2812 2082 2842 2157
rect 2896 2083 2926 2157
rect 2788 2066 2842 2082
rect 2788 2032 2798 2066
rect 2832 2032 2842 2066
rect 2788 2016 2842 2032
rect 2884 2067 2938 2083
rect 2884 2033 2894 2067
rect 2928 2033 2938 2067
rect 2884 2017 2938 2033
rect 2444 1985 2498 2001
rect 2444 1951 2454 1985
rect 2488 1951 2498 1985
rect 2444 1935 2498 1951
rect 2551 1985 2615 2001
rect 2551 1951 2571 1985
rect 2605 1951 2615 1985
rect 2456 1875 2486 1935
rect 2551 1920 2615 1951
rect 2540 1890 2758 1920
rect 2540 1875 2570 1890
rect 2728 1875 2758 1890
rect 2812 1875 2842 2016
rect 2896 1875 2926 2017
rect 2980 1978 3010 2157
rect 3070 2089 3100 2157
rect 3990 2237 4020 2263
rect 4089 2237 4119 2263
rect 4185 2237 4215 2263
rect 4257 2237 4287 2263
rect 4353 2237 4383 2263
rect 4442 2237 4472 2263
rect 4526 2237 4556 2263
rect 4610 2237 4640 2263
rect 4798 2237 4828 2263
rect 4882 2237 4912 2263
rect 4966 2237 4996 2263
rect 5050 2237 5080 2263
rect 5140 2237 5170 2263
rect 5239 2237 5269 2263
rect 5942 2237 5972 2263
rect 6041 2237 6071 2263
rect 6137 2237 6167 2263
rect 6209 2237 6239 2263
rect 6305 2237 6335 2263
rect 6394 2237 6424 2263
rect 6478 2237 6508 2263
rect 6562 2237 6592 2263
rect 6750 2237 6780 2263
rect 6834 2237 6864 2263
rect 6918 2237 6948 2263
rect 7002 2237 7032 2263
rect 7092 2237 7122 2263
rect 7191 2237 7221 2263
rect 7944 2243 7974 2269
rect 8043 2243 8073 2269
rect 8139 2243 8169 2269
rect 8211 2243 8241 2269
rect 8307 2243 8337 2269
rect 8396 2243 8426 2269
rect 8480 2243 8510 2269
rect 8564 2243 8594 2269
rect 8752 2243 8782 2269
rect 8836 2243 8866 2269
rect 8920 2243 8950 2269
rect 9004 2243 9034 2269
rect 9094 2243 9124 2269
rect 9193 2243 9223 2269
rect 9896 2243 9926 2269
rect 9995 2243 10025 2269
rect 10091 2243 10121 2269
rect 10163 2243 10193 2269
rect 10259 2243 10289 2269
rect 10348 2243 10378 2269
rect 10432 2243 10462 2269
rect 10516 2243 10546 2269
rect 10704 2243 10734 2269
rect 10788 2243 10818 2269
rect 10872 2243 10902 2269
rect 10956 2243 10986 2269
rect 11046 2243 11076 2269
rect 11145 2243 11175 2269
rect 11888 2243 11918 2269
rect 11987 2243 12017 2269
rect 12083 2243 12113 2269
rect 12155 2243 12185 2269
rect 12251 2243 12281 2269
rect 12340 2243 12370 2269
rect 12424 2243 12454 2269
rect 12508 2243 12538 2269
rect 12696 2243 12726 2269
rect 12780 2243 12810 2269
rect 12864 2243 12894 2269
rect 12948 2243 12978 2269
rect 13038 2243 13068 2269
rect 13137 2243 13167 2269
rect 13840 2243 13870 2269
rect 13939 2243 13969 2269
rect 14035 2243 14065 2269
rect 14107 2243 14137 2269
rect 14203 2243 14233 2269
rect 14292 2243 14322 2269
rect 14376 2243 14406 2269
rect 14460 2243 14490 2269
rect 14648 2243 14678 2269
rect 14732 2243 14762 2269
rect 14816 2243 14846 2269
rect 14900 2243 14930 2269
rect 14990 2243 15020 2269
rect 15089 2243 15119 2269
rect 15904 2243 15934 2269
rect 16003 2243 16033 2269
rect 16099 2243 16129 2269
rect 16171 2243 16201 2269
rect 16267 2243 16297 2269
rect 16356 2243 16386 2269
rect 16440 2243 16470 2269
rect 16524 2243 16554 2269
rect 16712 2243 16742 2269
rect 16796 2243 16826 2269
rect 16880 2243 16910 2269
rect 16964 2243 16994 2269
rect 17054 2243 17084 2269
rect 17153 2243 17183 2269
rect 3169 2089 3199 2111
rect 3052 2073 3106 2089
rect 3052 2039 3062 2073
rect 3096 2039 3106 2073
rect 3052 2023 3106 2039
rect 3148 2073 3202 2089
rect 3148 2039 3158 2073
rect 3192 2039 3202 2073
rect 3148 2023 3202 2039
rect 3990 2085 4020 2107
rect 4089 2093 4119 2153
rect 3990 2069 4044 2085
rect 3990 2035 4000 2069
rect 4034 2035 4044 2069
rect 2974 1962 3028 1978
rect 2974 1928 2984 1962
rect 3018 1928 3028 1962
rect 2974 1912 3028 1928
rect 2980 1875 3010 1912
rect 3070 1875 3100 2023
rect 3169 1991 3199 2023
rect 3990 2019 4044 2035
rect 4089 2077 4143 2093
rect 4089 2043 4099 2077
rect 4133 2043 4143 2077
rect 4089 2027 4143 2043
rect 3990 1987 4020 2019
rect 1920 1765 1950 1791
rect 2019 1765 2049 1791
rect 2115 1765 2145 1791
rect 2187 1765 2217 1791
rect 2283 1765 2313 1791
rect 2372 1765 2402 1791
rect 2456 1765 2486 1791
rect 2540 1765 2570 1791
rect 2728 1765 2758 1791
rect 2812 1765 2842 1791
rect 2896 1765 2926 1791
rect 2980 1765 3010 1791
rect 3070 1765 3100 1791
rect 3169 1765 3199 1791
rect 4089 1871 4119 2027
rect 4185 1981 4215 2153
rect 4161 1965 4215 1981
rect 4161 1931 4171 1965
rect 4205 1931 4215 1965
rect 4161 1915 4215 1931
rect 4185 1871 4215 1915
rect 4257 1981 4287 2153
rect 4353 2109 4383 2153
rect 4442 2109 4472 2153
rect 4526 2138 4556 2153
rect 4329 2093 4383 2109
rect 4329 2059 4339 2093
rect 4373 2059 4383 2093
rect 4329 2043 4383 2059
rect 4429 2093 4483 2109
rect 4429 2059 4439 2093
rect 4473 2059 4483 2093
rect 4429 2043 4483 2059
rect 4525 2108 4556 2138
rect 4610 2138 4640 2153
rect 4798 2138 4828 2153
rect 4610 2108 4828 2138
rect 4257 1965 4311 1981
rect 4257 1931 4267 1965
rect 4301 1931 4311 1965
rect 4257 1915 4311 1931
rect 4257 1871 4287 1915
rect 4353 1871 4383 2043
rect 4442 1871 4472 2043
rect 4525 1997 4555 2108
rect 4610 2093 4651 2108
rect 4621 1997 4651 2093
rect 4882 2078 4912 2153
rect 4966 2079 4996 2153
rect 4858 2062 4912 2078
rect 4858 2028 4868 2062
rect 4902 2028 4912 2062
rect 4858 2012 4912 2028
rect 4954 2063 5008 2079
rect 4954 2029 4964 2063
rect 4998 2029 5008 2063
rect 4954 2013 5008 2029
rect 4514 1981 4568 1997
rect 4514 1947 4524 1981
rect 4558 1947 4568 1981
rect 4514 1931 4568 1947
rect 4621 1981 4685 1997
rect 4621 1947 4641 1981
rect 4675 1947 4685 1981
rect 4526 1871 4556 1931
rect 4621 1916 4685 1947
rect 4610 1886 4828 1916
rect 4610 1871 4640 1886
rect 4798 1871 4828 1886
rect 4882 1871 4912 2012
rect 4966 1871 4996 2013
rect 5050 1974 5080 2153
rect 5140 2085 5170 2153
rect 5239 2085 5269 2107
rect 5942 2085 5972 2107
rect 6041 2093 6071 2153
rect 5122 2069 5176 2085
rect 5122 2035 5132 2069
rect 5166 2035 5176 2069
rect 5122 2019 5176 2035
rect 5218 2069 5272 2085
rect 5218 2035 5228 2069
rect 5262 2035 5272 2069
rect 5218 2019 5272 2035
rect 5942 2069 5996 2085
rect 5942 2035 5952 2069
rect 5986 2035 5996 2069
rect 5942 2019 5996 2035
rect 6041 2077 6095 2093
rect 6041 2043 6051 2077
rect 6085 2043 6095 2077
rect 6041 2027 6095 2043
rect 5044 1958 5098 1974
rect 5044 1924 5054 1958
rect 5088 1924 5098 1958
rect 5044 1908 5098 1924
rect 5050 1871 5080 1908
rect 5140 1871 5170 2019
rect 5239 1987 5269 2019
rect 5942 1987 5972 2019
rect 6041 1871 6071 2027
rect 6137 1981 6167 2153
rect 6113 1965 6167 1981
rect 6113 1931 6123 1965
rect 6157 1931 6167 1965
rect 6113 1915 6167 1931
rect 6137 1871 6167 1915
rect 6209 1981 6239 2153
rect 6305 2109 6335 2153
rect 6394 2109 6424 2153
rect 6478 2138 6508 2153
rect 6281 2093 6335 2109
rect 6281 2059 6291 2093
rect 6325 2059 6335 2093
rect 6281 2043 6335 2059
rect 6381 2093 6435 2109
rect 6381 2059 6391 2093
rect 6425 2059 6435 2093
rect 6381 2043 6435 2059
rect 6477 2108 6508 2138
rect 6562 2138 6592 2153
rect 6750 2138 6780 2153
rect 6562 2108 6780 2138
rect 6209 1965 6263 1981
rect 6209 1931 6219 1965
rect 6253 1931 6263 1965
rect 6209 1915 6263 1931
rect 6209 1871 6239 1915
rect 6305 1871 6335 2043
rect 6394 1871 6424 2043
rect 6477 1997 6507 2108
rect 6562 2093 6603 2108
rect 6573 1997 6603 2093
rect 6834 2078 6864 2153
rect 6918 2079 6948 2153
rect 6810 2062 6864 2078
rect 6810 2028 6820 2062
rect 6854 2028 6864 2062
rect 6810 2012 6864 2028
rect 6906 2063 6960 2079
rect 6906 2029 6916 2063
rect 6950 2029 6960 2063
rect 6906 2013 6960 2029
rect 6466 1981 6520 1997
rect 6466 1947 6476 1981
rect 6510 1947 6520 1981
rect 6466 1931 6520 1947
rect 6573 1981 6637 1997
rect 6573 1947 6593 1981
rect 6627 1947 6637 1981
rect 6478 1871 6508 1931
rect 6573 1916 6637 1947
rect 6562 1886 6780 1916
rect 6562 1871 6592 1886
rect 6750 1871 6780 1886
rect 6834 1871 6864 2012
rect 6918 1871 6948 2013
rect 7002 1974 7032 2153
rect 7092 2085 7122 2153
rect 7191 2085 7221 2107
rect 7944 2091 7974 2113
rect 8043 2099 8073 2159
rect 7074 2069 7128 2085
rect 7074 2035 7084 2069
rect 7118 2035 7128 2069
rect 7074 2019 7128 2035
rect 7170 2069 7224 2085
rect 7170 2035 7180 2069
rect 7214 2035 7224 2069
rect 7170 2019 7224 2035
rect 7944 2075 7998 2091
rect 7944 2041 7954 2075
rect 7988 2041 7998 2075
rect 7944 2025 7998 2041
rect 8043 2083 8097 2099
rect 8043 2049 8053 2083
rect 8087 2049 8097 2083
rect 8043 2033 8097 2049
rect 6996 1958 7050 1974
rect 6996 1924 7006 1958
rect 7040 1924 7050 1958
rect 6996 1908 7050 1924
rect 7002 1871 7032 1908
rect 7092 1871 7122 2019
rect 7191 1987 7221 2019
rect 7944 1993 7974 2025
rect 8043 1877 8073 2033
rect 8139 1987 8169 2159
rect 8115 1971 8169 1987
rect 8115 1937 8125 1971
rect 8159 1937 8169 1971
rect 8115 1921 8169 1937
rect 8139 1877 8169 1921
rect 8211 1987 8241 2159
rect 8307 2115 8337 2159
rect 8396 2115 8426 2159
rect 8480 2144 8510 2159
rect 8283 2099 8337 2115
rect 8283 2065 8293 2099
rect 8327 2065 8337 2099
rect 8283 2049 8337 2065
rect 8383 2099 8437 2115
rect 8383 2065 8393 2099
rect 8427 2065 8437 2099
rect 8383 2049 8437 2065
rect 8479 2114 8510 2144
rect 8564 2144 8594 2159
rect 8752 2144 8782 2159
rect 8564 2114 8782 2144
rect 8211 1971 8265 1987
rect 8211 1937 8221 1971
rect 8255 1937 8265 1971
rect 8211 1921 8265 1937
rect 8211 1877 8241 1921
rect 8307 1877 8337 2049
rect 8396 1877 8426 2049
rect 8479 2003 8509 2114
rect 8564 2099 8605 2114
rect 8575 2003 8605 2099
rect 8836 2084 8866 2159
rect 8920 2085 8950 2159
rect 8812 2068 8866 2084
rect 8812 2034 8822 2068
rect 8856 2034 8866 2068
rect 8812 2018 8866 2034
rect 8908 2069 8962 2085
rect 8908 2035 8918 2069
rect 8952 2035 8962 2069
rect 8908 2019 8962 2035
rect 8468 1987 8522 2003
rect 8468 1953 8478 1987
rect 8512 1953 8522 1987
rect 8468 1937 8522 1953
rect 8575 1987 8639 2003
rect 8575 1953 8595 1987
rect 8629 1953 8639 1987
rect 8480 1877 8510 1937
rect 8575 1922 8639 1953
rect 8564 1892 8782 1922
rect 8564 1877 8594 1892
rect 8752 1877 8782 1892
rect 8836 1877 8866 2018
rect 8920 1877 8950 2019
rect 9004 1980 9034 2159
rect 9094 2091 9124 2159
rect 9193 2091 9223 2113
rect 9896 2091 9926 2113
rect 9995 2099 10025 2159
rect 9076 2075 9130 2091
rect 9076 2041 9086 2075
rect 9120 2041 9130 2075
rect 9076 2025 9130 2041
rect 9172 2075 9226 2091
rect 9172 2041 9182 2075
rect 9216 2041 9226 2075
rect 9172 2025 9226 2041
rect 9896 2075 9950 2091
rect 9896 2041 9906 2075
rect 9940 2041 9950 2075
rect 9896 2025 9950 2041
rect 9995 2083 10049 2099
rect 9995 2049 10005 2083
rect 10039 2049 10049 2083
rect 9995 2033 10049 2049
rect 8998 1964 9052 1980
rect 8998 1930 9008 1964
rect 9042 1930 9052 1964
rect 8998 1914 9052 1930
rect 9004 1877 9034 1914
rect 9094 1877 9124 2025
rect 9193 1993 9223 2025
rect 9896 1993 9926 2025
rect 9995 1877 10025 2033
rect 10091 1987 10121 2159
rect 10067 1971 10121 1987
rect 10067 1937 10077 1971
rect 10111 1937 10121 1971
rect 10067 1921 10121 1937
rect 10091 1877 10121 1921
rect 10163 1987 10193 2159
rect 10259 2115 10289 2159
rect 10348 2115 10378 2159
rect 10432 2144 10462 2159
rect 10235 2099 10289 2115
rect 10235 2065 10245 2099
rect 10279 2065 10289 2099
rect 10235 2049 10289 2065
rect 10335 2099 10389 2115
rect 10335 2065 10345 2099
rect 10379 2065 10389 2099
rect 10335 2049 10389 2065
rect 10431 2114 10462 2144
rect 10516 2144 10546 2159
rect 10704 2144 10734 2159
rect 10516 2114 10734 2144
rect 10163 1971 10217 1987
rect 10163 1937 10173 1971
rect 10207 1937 10217 1971
rect 10163 1921 10217 1937
rect 10163 1877 10193 1921
rect 10259 1877 10289 2049
rect 10348 1877 10378 2049
rect 10431 2003 10461 2114
rect 10516 2099 10557 2114
rect 10527 2003 10557 2099
rect 10788 2084 10818 2159
rect 10872 2085 10902 2159
rect 10764 2068 10818 2084
rect 10764 2034 10774 2068
rect 10808 2034 10818 2068
rect 10764 2018 10818 2034
rect 10860 2069 10914 2085
rect 10860 2035 10870 2069
rect 10904 2035 10914 2069
rect 10860 2019 10914 2035
rect 10420 1987 10474 2003
rect 10420 1953 10430 1987
rect 10464 1953 10474 1987
rect 10420 1937 10474 1953
rect 10527 1987 10591 2003
rect 10527 1953 10547 1987
rect 10581 1953 10591 1987
rect 10432 1877 10462 1937
rect 10527 1922 10591 1953
rect 10516 1892 10734 1922
rect 10516 1877 10546 1892
rect 10704 1877 10734 1892
rect 10788 1877 10818 2018
rect 10872 1877 10902 2019
rect 10956 1980 10986 2159
rect 11046 2091 11076 2159
rect 11145 2091 11175 2113
rect 11888 2091 11918 2113
rect 11987 2099 12017 2159
rect 11028 2075 11082 2091
rect 11028 2041 11038 2075
rect 11072 2041 11082 2075
rect 11028 2025 11082 2041
rect 11124 2075 11178 2091
rect 11124 2041 11134 2075
rect 11168 2041 11178 2075
rect 11124 2025 11178 2041
rect 11888 2075 11942 2091
rect 11888 2041 11898 2075
rect 11932 2041 11942 2075
rect 11888 2025 11942 2041
rect 11987 2083 12041 2099
rect 11987 2049 11997 2083
rect 12031 2049 12041 2083
rect 11987 2033 12041 2049
rect 10950 1964 11004 1980
rect 10950 1930 10960 1964
rect 10994 1930 11004 1964
rect 10950 1914 11004 1930
rect 10956 1877 10986 1914
rect 11046 1877 11076 2025
rect 11145 1993 11175 2025
rect 11888 1993 11918 2025
rect 11987 1877 12017 2033
rect 12083 1987 12113 2159
rect 12059 1971 12113 1987
rect 12059 1937 12069 1971
rect 12103 1937 12113 1971
rect 12059 1921 12113 1937
rect 12083 1877 12113 1921
rect 12155 1987 12185 2159
rect 12251 2115 12281 2159
rect 12340 2115 12370 2159
rect 12424 2144 12454 2159
rect 12227 2099 12281 2115
rect 12227 2065 12237 2099
rect 12271 2065 12281 2099
rect 12227 2049 12281 2065
rect 12327 2099 12381 2115
rect 12327 2065 12337 2099
rect 12371 2065 12381 2099
rect 12327 2049 12381 2065
rect 12423 2114 12454 2144
rect 12508 2144 12538 2159
rect 12696 2144 12726 2159
rect 12508 2114 12726 2144
rect 12155 1971 12209 1987
rect 12155 1937 12165 1971
rect 12199 1937 12209 1971
rect 12155 1921 12209 1937
rect 12155 1877 12185 1921
rect 12251 1877 12281 2049
rect 12340 1877 12370 2049
rect 12423 2003 12453 2114
rect 12508 2099 12549 2114
rect 12519 2003 12549 2099
rect 12780 2084 12810 2159
rect 12864 2085 12894 2159
rect 12756 2068 12810 2084
rect 12756 2034 12766 2068
rect 12800 2034 12810 2068
rect 12756 2018 12810 2034
rect 12852 2069 12906 2085
rect 12852 2035 12862 2069
rect 12896 2035 12906 2069
rect 12852 2019 12906 2035
rect 12412 1987 12466 2003
rect 12412 1953 12422 1987
rect 12456 1953 12466 1987
rect 12412 1937 12466 1953
rect 12519 1987 12583 2003
rect 12519 1953 12539 1987
rect 12573 1953 12583 1987
rect 12424 1877 12454 1937
rect 12519 1922 12583 1953
rect 12508 1892 12726 1922
rect 12508 1877 12538 1892
rect 12696 1877 12726 1892
rect 12780 1877 12810 2018
rect 12864 1877 12894 2019
rect 12948 1980 12978 2159
rect 13038 2091 13068 2159
rect 13137 2091 13167 2113
rect 13840 2091 13870 2113
rect 13939 2099 13969 2159
rect 13020 2075 13074 2091
rect 13020 2041 13030 2075
rect 13064 2041 13074 2075
rect 13020 2025 13074 2041
rect 13116 2075 13170 2091
rect 13116 2041 13126 2075
rect 13160 2041 13170 2075
rect 13116 2025 13170 2041
rect 13840 2075 13894 2091
rect 13840 2041 13850 2075
rect 13884 2041 13894 2075
rect 13840 2025 13894 2041
rect 13939 2083 13993 2099
rect 13939 2049 13949 2083
rect 13983 2049 13993 2083
rect 13939 2033 13993 2049
rect 12942 1964 12996 1980
rect 12942 1930 12952 1964
rect 12986 1930 12996 1964
rect 12942 1914 12996 1930
rect 12948 1877 12978 1914
rect 13038 1877 13068 2025
rect 13137 1993 13167 2025
rect 13840 1993 13870 2025
rect 13939 1877 13969 2033
rect 14035 1987 14065 2159
rect 14011 1971 14065 1987
rect 14011 1937 14021 1971
rect 14055 1937 14065 1971
rect 14011 1921 14065 1937
rect 14035 1877 14065 1921
rect 14107 1987 14137 2159
rect 14203 2115 14233 2159
rect 14292 2115 14322 2159
rect 14376 2144 14406 2159
rect 14179 2099 14233 2115
rect 14179 2065 14189 2099
rect 14223 2065 14233 2099
rect 14179 2049 14233 2065
rect 14279 2099 14333 2115
rect 14279 2065 14289 2099
rect 14323 2065 14333 2099
rect 14279 2049 14333 2065
rect 14375 2114 14406 2144
rect 14460 2144 14490 2159
rect 14648 2144 14678 2159
rect 14460 2114 14678 2144
rect 14107 1971 14161 1987
rect 14107 1937 14117 1971
rect 14151 1937 14161 1971
rect 14107 1921 14161 1937
rect 14107 1877 14137 1921
rect 14203 1877 14233 2049
rect 14292 1877 14322 2049
rect 14375 2003 14405 2114
rect 14460 2099 14501 2114
rect 14471 2003 14501 2099
rect 14732 2084 14762 2159
rect 14816 2085 14846 2159
rect 14708 2068 14762 2084
rect 14708 2034 14718 2068
rect 14752 2034 14762 2068
rect 14708 2018 14762 2034
rect 14804 2069 14858 2085
rect 14804 2035 14814 2069
rect 14848 2035 14858 2069
rect 14804 2019 14858 2035
rect 14364 1987 14418 2003
rect 14364 1953 14374 1987
rect 14408 1953 14418 1987
rect 14364 1937 14418 1953
rect 14471 1987 14535 2003
rect 14471 1953 14491 1987
rect 14525 1953 14535 1987
rect 14376 1877 14406 1937
rect 14471 1922 14535 1953
rect 14460 1892 14678 1922
rect 14460 1877 14490 1892
rect 14648 1877 14678 1892
rect 14732 1877 14762 2018
rect 14816 1877 14846 2019
rect 14900 1980 14930 2159
rect 14990 2091 15020 2159
rect 15089 2091 15119 2113
rect 15904 2091 15934 2113
rect 16003 2099 16033 2159
rect 14972 2075 15026 2091
rect 14972 2041 14982 2075
rect 15016 2041 15026 2075
rect 14972 2025 15026 2041
rect 15068 2075 15122 2091
rect 15068 2041 15078 2075
rect 15112 2041 15122 2075
rect 15068 2025 15122 2041
rect 15904 2075 15958 2091
rect 15904 2041 15914 2075
rect 15948 2041 15958 2075
rect 15904 2025 15958 2041
rect 16003 2083 16057 2099
rect 16003 2049 16013 2083
rect 16047 2049 16057 2083
rect 16003 2033 16057 2049
rect 14894 1964 14948 1980
rect 14894 1930 14904 1964
rect 14938 1930 14948 1964
rect 14894 1914 14948 1930
rect 14900 1877 14930 1914
rect 14990 1877 15020 2025
rect 15089 1993 15119 2025
rect 15904 1993 15934 2025
rect 16003 1877 16033 2033
rect 16099 1987 16129 2159
rect 16075 1971 16129 1987
rect 16075 1937 16085 1971
rect 16119 1937 16129 1971
rect 16075 1921 16129 1937
rect 16099 1877 16129 1921
rect 16171 1987 16201 2159
rect 16267 2115 16297 2159
rect 16356 2115 16386 2159
rect 16440 2144 16470 2159
rect 16243 2099 16297 2115
rect 16243 2065 16253 2099
rect 16287 2065 16297 2099
rect 16243 2049 16297 2065
rect 16343 2099 16397 2115
rect 16343 2065 16353 2099
rect 16387 2065 16397 2099
rect 16343 2049 16397 2065
rect 16439 2114 16470 2144
rect 16524 2144 16554 2159
rect 16712 2144 16742 2159
rect 16524 2114 16742 2144
rect 16171 1971 16225 1987
rect 16171 1937 16181 1971
rect 16215 1937 16225 1971
rect 16171 1921 16225 1937
rect 16171 1877 16201 1921
rect 16267 1877 16297 2049
rect 16356 1877 16386 2049
rect 16439 2003 16469 2114
rect 16524 2099 16565 2114
rect 16535 2003 16565 2099
rect 16796 2084 16826 2159
rect 16880 2085 16910 2159
rect 16772 2068 16826 2084
rect 16772 2034 16782 2068
rect 16816 2034 16826 2068
rect 16772 2018 16826 2034
rect 16868 2069 16922 2085
rect 16868 2035 16878 2069
rect 16912 2035 16922 2069
rect 16868 2019 16922 2035
rect 16428 1987 16482 2003
rect 16428 1953 16438 1987
rect 16472 1953 16482 1987
rect 16428 1937 16482 1953
rect 16535 1987 16599 2003
rect 16535 1953 16555 1987
rect 16589 1953 16599 1987
rect 16440 1877 16470 1937
rect 16535 1922 16599 1953
rect 16524 1892 16742 1922
rect 16524 1877 16554 1892
rect 16712 1877 16742 1892
rect 16796 1877 16826 2018
rect 16880 1877 16910 2019
rect 16964 1980 16994 2159
rect 17054 2091 17084 2159
rect 17153 2091 17183 2113
rect 17036 2075 17090 2091
rect 17036 2041 17046 2075
rect 17080 2041 17090 2075
rect 17036 2025 17090 2041
rect 17132 2075 17186 2091
rect 17132 2041 17142 2075
rect 17176 2041 17186 2075
rect 17132 2025 17186 2041
rect 16958 1964 17012 1980
rect 16958 1930 16968 1964
rect 17002 1930 17012 1964
rect 16958 1914 17012 1930
rect 16964 1877 16994 1914
rect 17054 1877 17084 2025
rect 17153 1993 17183 2025
rect 3990 1761 4020 1787
rect 4089 1761 4119 1787
rect 4185 1761 4215 1787
rect 4257 1761 4287 1787
rect 4353 1761 4383 1787
rect 4442 1761 4472 1787
rect 4526 1761 4556 1787
rect 4610 1761 4640 1787
rect 4798 1761 4828 1787
rect 4882 1761 4912 1787
rect 4966 1761 4996 1787
rect 5050 1761 5080 1787
rect 5140 1761 5170 1787
rect 5239 1761 5269 1787
rect 5942 1761 5972 1787
rect 6041 1761 6071 1787
rect 6137 1761 6167 1787
rect 6209 1761 6239 1787
rect 6305 1761 6335 1787
rect 6394 1761 6424 1787
rect 6478 1761 6508 1787
rect 6562 1761 6592 1787
rect 6750 1761 6780 1787
rect 6834 1761 6864 1787
rect 6918 1761 6948 1787
rect 7002 1761 7032 1787
rect 7092 1761 7122 1787
rect 7191 1761 7221 1787
rect 7944 1767 7974 1793
rect 8043 1767 8073 1793
rect 8139 1767 8169 1793
rect 8211 1767 8241 1793
rect 8307 1767 8337 1793
rect 8396 1767 8426 1793
rect 8480 1767 8510 1793
rect 8564 1767 8594 1793
rect 8752 1767 8782 1793
rect 8836 1767 8866 1793
rect 8920 1767 8950 1793
rect 9004 1767 9034 1793
rect 9094 1767 9124 1793
rect 9193 1767 9223 1793
rect 9896 1767 9926 1793
rect 9995 1767 10025 1793
rect 10091 1767 10121 1793
rect 10163 1767 10193 1793
rect 10259 1767 10289 1793
rect 10348 1767 10378 1793
rect 10432 1767 10462 1793
rect 10516 1767 10546 1793
rect 10704 1767 10734 1793
rect 10788 1767 10818 1793
rect 10872 1767 10902 1793
rect 10956 1767 10986 1793
rect 11046 1767 11076 1793
rect 11145 1767 11175 1793
rect 11888 1767 11918 1793
rect 11987 1767 12017 1793
rect 12083 1767 12113 1793
rect 12155 1767 12185 1793
rect 12251 1767 12281 1793
rect 12340 1767 12370 1793
rect 12424 1767 12454 1793
rect 12508 1767 12538 1793
rect 12696 1767 12726 1793
rect 12780 1767 12810 1793
rect 12864 1767 12894 1793
rect 12948 1767 12978 1793
rect 13038 1767 13068 1793
rect 13137 1767 13167 1793
rect 13840 1767 13870 1793
rect 13939 1767 13969 1793
rect 14035 1767 14065 1793
rect 14107 1767 14137 1793
rect 14203 1767 14233 1793
rect 14292 1767 14322 1793
rect 14376 1767 14406 1793
rect 14460 1767 14490 1793
rect 14648 1767 14678 1793
rect 14732 1767 14762 1793
rect 14816 1767 14846 1793
rect 14900 1767 14930 1793
rect 14990 1767 15020 1793
rect 15089 1767 15119 1793
rect 15904 1767 15934 1793
rect 16003 1767 16033 1793
rect 16099 1767 16129 1793
rect 16171 1767 16201 1793
rect 16267 1767 16297 1793
rect 16356 1767 16386 1793
rect 16440 1767 16470 1793
rect 16524 1767 16554 1793
rect 16712 1767 16742 1793
rect 16796 1767 16826 1793
rect 16880 1767 16910 1793
rect 16964 1767 16994 1793
rect 17054 1767 17084 1793
rect 17153 1767 17183 1793
<< polycont >>
rect 18761 35001 18795 35035
rect 18761 34740 18795 34774
rect 18761 34556 18795 34590
rect 18645 34482 18679 34516
rect 18645 34346 18679 34380
rect 18711 34244 18745 34278
rect 18819 34287 18853 34321
rect 18711 34108 18745 34142
rect 18807 34044 18841 34078
rect 18645 33934 18679 33968
rect 18723 33825 18757 33859
rect 18819 33845 18853 33879
rect 18693 33682 18727 33716
rect 18746 33520 18780 33554
rect 18761 33418 18795 33452
rect 18769 32695 18803 32729
rect 18769 32434 18803 32468
rect 18769 32250 18803 32284
rect 18653 32176 18687 32210
rect 18653 32040 18687 32074
rect 18719 31938 18753 31972
rect 18827 31981 18861 32015
rect 18719 31802 18753 31836
rect 18815 31738 18849 31772
rect 18653 31628 18687 31662
rect 18731 31519 18765 31553
rect 18827 31539 18861 31573
rect 18701 31376 18735 31410
rect 18754 31214 18788 31248
rect 18769 31112 18803 31146
rect 18777 30481 18811 30515
rect 18777 30220 18811 30254
rect 18777 30036 18811 30070
rect 18661 29962 18695 29996
rect 18661 29826 18695 29860
rect 18727 29724 18761 29758
rect 18835 29767 18869 29801
rect 18727 29588 18761 29622
rect 18823 29524 18857 29558
rect 18661 29414 18695 29448
rect 18739 29305 18773 29339
rect 18835 29325 18869 29359
rect 18709 29162 18743 29196
rect 18762 29000 18796 29034
rect 18777 28898 18811 28932
rect 18759 28281 18793 28315
rect 18759 28020 18793 28054
rect 18759 27836 18793 27870
rect 18643 27762 18677 27796
rect 18643 27626 18677 27660
rect 18709 27524 18743 27558
rect 18817 27567 18851 27601
rect 18709 27388 18743 27422
rect 18805 27324 18839 27358
rect 18643 27214 18677 27248
rect 18721 27105 18755 27139
rect 18817 27125 18851 27159
rect 18691 26962 18725 26996
rect 18744 26800 18778 26834
rect 18759 26698 18793 26732
rect 18767 26067 18801 26101
rect 18767 25806 18801 25840
rect 18767 25622 18801 25656
rect 18651 25548 18685 25582
rect 18651 25412 18685 25446
rect 18717 25310 18751 25344
rect 18825 25353 18859 25387
rect 18717 25174 18751 25208
rect 18813 25110 18847 25144
rect 18651 25000 18685 25034
rect 18729 24891 18763 24925
rect 18825 24911 18859 24945
rect 18699 24748 18733 24782
rect 18752 24586 18786 24620
rect 18767 24484 18801 24518
rect 7578 23059 7612 23093
rect 7842 23127 7876 23161
rect 8094 23175 8128 23209
rect 7680 23074 7714 23108
rect 7985 23097 8019 23131
rect 8005 23001 8039 23035
rect 8506 23175 8540 23209
rect 8642 23175 8676 23209
rect 8268 23109 8302 23143
rect 8404 23109 8438 23143
rect 8204 23013 8238 23047
rect 8447 23001 8481 23035
rect 8716 23059 8750 23093
rect 8900 23059 8934 23093
rect 9161 23059 9195 23093
rect 9792 23067 9826 23101
rect 10056 23135 10090 23169
rect 10308 23183 10342 23217
rect 9894 23082 9928 23116
rect 10199 23105 10233 23139
rect 10219 23009 10253 23043
rect 10720 23183 10754 23217
rect 10856 23183 10890 23217
rect 10482 23117 10516 23151
rect 10618 23117 10652 23151
rect 10418 23021 10452 23055
rect 10661 23009 10695 23043
rect 10930 23067 10964 23101
rect 11114 23067 11148 23101
rect 11375 23067 11409 23101
rect 11992 23049 12026 23083
rect 12256 23117 12290 23151
rect 12508 23165 12542 23199
rect 12094 23064 12128 23098
rect 12399 23087 12433 23121
rect 12419 22991 12453 23025
rect 12920 23165 12954 23199
rect 13056 23165 13090 23199
rect 12682 23099 12716 23133
rect 12818 23099 12852 23133
rect 12618 23003 12652 23037
rect 12861 22991 12895 23025
rect 13130 23049 13164 23083
rect 13314 23049 13348 23083
rect 13575 23049 13609 23083
rect 14206 23057 14240 23091
rect 14470 23125 14504 23159
rect 14722 23173 14756 23207
rect 14308 23072 14342 23106
rect 14613 23095 14647 23129
rect 14633 22999 14667 23033
rect 15134 23173 15168 23207
rect 15270 23173 15304 23207
rect 14896 23107 14930 23141
rect 15032 23107 15066 23141
rect 14832 23011 14866 23045
rect 15075 22999 15109 23033
rect 15344 23057 15378 23091
rect 15528 23057 15562 23091
rect 15789 23057 15823 23091
rect 16512 23065 16546 23099
rect 16776 23133 16810 23167
rect 17028 23181 17062 23215
rect 16614 23080 16648 23114
rect 16919 23103 16953 23137
rect 16939 23007 16973 23041
rect 17440 23181 17474 23215
rect 17576 23181 17610 23215
rect 17202 23115 17236 23149
rect 17338 23115 17372 23149
rect 17138 23019 17172 23053
rect 17381 23007 17415 23041
rect 17650 23065 17684 23099
rect 17834 23065 17868 23099
rect 18095 23065 18129 23099
rect 15729 17397 15763 17431
rect 16507 17435 16541 17469
rect 17381 17437 17415 17471
rect 18149 17427 18183 17461
rect 19271 17429 19305 17463
rect 20145 17431 20179 17465
rect 20913 17421 20947 17455
rect 21527 17419 21561 17453
rect 22401 17421 22435 17455
rect 23169 17411 23203 17445
rect 9419 16261 9453 16295
rect 9536 16261 9570 16295
rect 9671 16261 9705 16295
rect 9767 16261 9801 16295
rect 9506 15517 9540 15551
rect 9647 15517 9681 15551
rect 9755 15517 9789 15551
rect 11505 15407 11539 15441
rect 11651 15407 11685 15441
rect 11757 15407 11791 15441
rect 11853 15407 11887 15441
rect 11964 15407 11998 15441
rect 10690 14907 10724 14941
rect 10831 14907 10865 14941
rect 10939 14907 10973 14941
rect 9429 14697 9463 14731
rect 9546 14697 9580 14731
rect 9681 14697 9715 14731
rect 9777 14697 9811 14731
rect 9516 13953 9550 13987
rect 9657 13953 9691 13987
rect 12845 14149 12879 14183
rect 9765 13953 9799 13987
rect 10721 13941 10755 13975
rect 10867 13941 10901 13975
rect 10973 13941 11007 13975
rect 11069 13941 11103 13975
rect 11180 13941 11214 13975
rect 12623 13925 12657 13959
rect 12749 13925 12783 13959
rect 12925 13925 12959 13959
rect 13021 13925 13055 13959
rect 11726 13567 11760 13601
rect 11862 13567 11896 13601
rect 11965 13567 11999 13601
rect 10987 13326 11021 13360
rect 9421 13029 9455 13063
rect 9538 13029 9572 13063
rect 9673 13029 9707 13063
rect 9769 13029 9803 13063
rect 10849 13053 10883 13087
rect 11059 13093 11093 13127
rect 11155 13099 11189 13133
rect 9508 12285 9542 12319
rect 9649 12285 9683 12319
rect 9757 12285 9791 12319
rect 10884 12079 10918 12113
rect 11025 12079 11059 12113
rect 11133 12079 11167 12113
rect 9431 11465 9465 11499
rect 9548 11465 9582 11499
rect 9683 11465 9717 11499
rect 9779 11465 9813 11499
rect 9518 10721 9552 10755
rect 9659 10721 9693 10755
rect 9767 10721 9801 10755
rect 6274 6351 6308 6385
rect 10142 5719 10176 5753
rect 10241 5727 10275 5761
rect 1960 5299 1994 5333
rect 2059 5307 2093 5341
rect 2131 5195 2165 5229
rect 2299 5323 2333 5357
rect 2399 5323 2433 5357
rect 2227 5195 2261 5229
rect 2828 5292 2862 5326
rect 2924 5293 2958 5327
rect 2484 5211 2518 5245
rect 2601 5211 2635 5245
rect 3092 5299 3126 5333
rect 3188 5299 3222 5333
rect 4094 5291 4128 5325
rect 3014 5188 3048 5222
rect 4193 5299 4227 5333
rect 4265 5187 4299 5221
rect 4433 5315 4467 5349
rect 4533 5315 4567 5349
rect 4361 5187 4395 5221
rect 4962 5284 4996 5318
rect 5058 5285 5092 5319
rect 4618 5203 4652 5237
rect 4735 5203 4769 5237
rect 5226 5291 5260 5325
rect 5322 5291 5356 5325
rect 6046 5291 6080 5325
rect 6145 5299 6179 5333
rect 5148 5180 5182 5214
rect 6217 5187 6251 5221
rect 6385 5315 6419 5349
rect 6485 5315 6519 5349
rect 6313 5187 6347 5221
rect 6914 5284 6948 5318
rect 7010 5285 7044 5319
rect 6570 5203 6604 5237
rect 6687 5203 6721 5237
rect 7178 5291 7212 5325
rect 7274 5291 7308 5325
rect 8048 5297 8082 5331
rect 8147 5305 8181 5339
rect 7100 5180 7134 5214
rect 8219 5193 8253 5227
rect 8387 5321 8421 5355
rect 8487 5321 8521 5355
rect 8315 5193 8349 5227
rect 8916 5290 8950 5324
rect 9012 5291 9046 5325
rect 8572 5209 8606 5243
rect 8689 5209 8723 5243
rect 10313 5615 10347 5649
rect 10481 5743 10515 5777
rect 10581 5743 10615 5777
rect 10409 5615 10443 5649
rect 11010 5712 11044 5746
rect 11106 5713 11140 5747
rect 10666 5631 10700 5665
rect 10783 5631 10817 5665
rect 11274 5719 11308 5753
rect 11370 5719 11404 5753
rect 12204 5707 12238 5741
rect 11196 5608 11230 5642
rect 12303 5715 12337 5749
rect 12375 5603 12409 5637
rect 12543 5731 12577 5765
rect 12643 5731 12677 5765
rect 12471 5603 12505 5637
rect 13072 5700 13106 5734
rect 13168 5701 13202 5735
rect 12728 5619 12762 5653
rect 12845 5619 12879 5653
rect 13336 5707 13370 5741
rect 13432 5707 13466 5741
rect 14162 5715 14196 5749
rect 14261 5723 14295 5757
rect 13258 5596 13292 5630
rect 14333 5611 14367 5645
rect 14501 5739 14535 5773
rect 14601 5739 14635 5773
rect 14429 5611 14463 5645
rect 15030 5708 15064 5742
rect 15126 5709 15160 5743
rect 14686 5627 14720 5661
rect 14803 5627 14837 5661
rect 15294 5715 15328 5749
rect 15390 5715 15424 5749
rect 16156 5721 16190 5755
rect 16255 5729 16289 5763
rect 15216 5604 15250 5638
rect 16327 5617 16361 5651
rect 16495 5745 16529 5779
rect 16595 5745 16629 5779
rect 16423 5617 16457 5651
rect 17024 5714 17058 5748
rect 17120 5715 17154 5749
rect 16680 5633 16714 5667
rect 16797 5633 16831 5667
rect 17288 5721 17322 5755
rect 17384 5721 17418 5755
rect 17210 5610 17244 5644
rect 9180 5297 9214 5331
rect 9276 5297 9310 5331
rect 9102 5186 9136 5220
rect 10170 4845 10204 4879
rect 10269 4853 10303 4887
rect 10341 4741 10375 4775
rect 10509 4869 10543 4903
rect 10609 4869 10643 4903
rect 10437 4741 10471 4775
rect 11038 4838 11072 4872
rect 11134 4839 11168 4873
rect 10694 4757 10728 4791
rect 10811 4757 10845 4791
rect 11302 4845 11336 4879
rect 11398 4845 11432 4879
rect 11224 4734 11258 4768
rect 12440 4801 12474 4835
rect 12539 4809 12573 4843
rect 12611 4697 12645 4731
rect 12779 4825 12813 4859
rect 12879 4825 12913 4859
rect 12707 4697 12741 4731
rect 13308 4794 13342 4828
rect 13404 4795 13438 4829
rect 12964 4713 12998 4747
rect 13081 4713 13115 4747
rect 13572 4801 13606 4835
rect 13668 4801 13702 4835
rect 14442 4795 14476 4829
rect 13494 4690 13528 4724
rect 14541 4803 14575 4837
rect 14613 4691 14647 4725
rect 14781 4819 14815 4853
rect 14881 4819 14915 4853
rect 14709 4691 14743 4725
rect 15310 4788 15344 4822
rect 15406 4789 15440 4823
rect 14966 4707 15000 4741
rect 15083 4707 15117 4741
rect 15574 4795 15608 4829
rect 15670 4795 15704 4829
rect 15496 4684 15530 4718
rect 16464 4777 16498 4811
rect 16563 4785 16597 4819
rect 16635 4673 16669 4707
rect 16803 4801 16837 4835
rect 16903 4801 16937 4835
rect 16731 4673 16765 4707
rect 17332 4770 17366 4804
rect 17428 4771 17462 4805
rect 16988 4689 17022 4723
rect 17105 4689 17139 4723
rect 17596 4777 17630 4811
rect 17692 4777 17726 4811
rect 17518 4666 17552 4700
rect 1930 2039 1964 2073
rect 2029 2047 2063 2081
rect 2101 1935 2135 1969
rect 2269 2063 2303 2097
rect 2369 2063 2403 2097
rect 2197 1935 2231 1969
rect 2798 2032 2832 2066
rect 2894 2033 2928 2067
rect 2454 1951 2488 1985
rect 2571 1951 2605 1985
rect 3062 2039 3096 2073
rect 3158 2039 3192 2073
rect 4000 2035 4034 2069
rect 2984 1928 3018 1962
rect 4099 2043 4133 2077
rect 4171 1931 4205 1965
rect 4339 2059 4373 2093
rect 4439 2059 4473 2093
rect 4267 1931 4301 1965
rect 4868 2028 4902 2062
rect 4964 2029 4998 2063
rect 4524 1947 4558 1981
rect 4641 1947 4675 1981
rect 5132 2035 5166 2069
rect 5228 2035 5262 2069
rect 5952 2035 5986 2069
rect 6051 2043 6085 2077
rect 5054 1924 5088 1958
rect 6123 1931 6157 1965
rect 6291 2059 6325 2093
rect 6391 2059 6425 2093
rect 6219 1931 6253 1965
rect 6820 2028 6854 2062
rect 6916 2029 6950 2063
rect 6476 1947 6510 1981
rect 6593 1947 6627 1981
rect 7084 2035 7118 2069
rect 7180 2035 7214 2069
rect 7954 2041 7988 2075
rect 8053 2049 8087 2083
rect 7006 1924 7040 1958
rect 8125 1937 8159 1971
rect 8293 2065 8327 2099
rect 8393 2065 8427 2099
rect 8221 1937 8255 1971
rect 8822 2034 8856 2068
rect 8918 2035 8952 2069
rect 8478 1953 8512 1987
rect 8595 1953 8629 1987
rect 9086 2041 9120 2075
rect 9182 2041 9216 2075
rect 9906 2041 9940 2075
rect 10005 2049 10039 2083
rect 9008 1930 9042 1964
rect 10077 1937 10111 1971
rect 10245 2065 10279 2099
rect 10345 2065 10379 2099
rect 10173 1937 10207 1971
rect 10774 2034 10808 2068
rect 10870 2035 10904 2069
rect 10430 1953 10464 1987
rect 10547 1953 10581 1987
rect 11038 2041 11072 2075
rect 11134 2041 11168 2075
rect 11898 2041 11932 2075
rect 11997 2049 12031 2083
rect 10960 1930 10994 1964
rect 12069 1937 12103 1971
rect 12237 2065 12271 2099
rect 12337 2065 12371 2099
rect 12165 1937 12199 1971
rect 12766 2034 12800 2068
rect 12862 2035 12896 2069
rect 12422 1953 12456 1987
rect 12539 1953 12573 1987
rect 13030 2041 13064 2075
rect 13126 2041 13160 2075
rect 13850 2041 13884 2075
rect 13949 2049 13983 2083
rect 12952 1930 12986 1964
rect 14021 1937 14055 1971
rect 14189 2065 14223 2099
rect 14289 2065 14323 2099
rect 14117 1937 14151 1971
rect 14718 2034 14752 2068
rect 14814 2035 14848 2069
rect 14374 1953 14408 1987
rect 14491 1953 14525 1987
rect 14982 2041 15016 2075
rect 15078 2041 15112 2075
rect 15914 2041 15948 2075
rect 16013 2049 16047 2083
rect 14904 1930 14938 1964
rect 16085 1937 16119 1971
rect 16253 2065 16287 2099
rect 16353 2065 16387 2099
rect 16181 1937 16215 1971
rect 16782 2034 16816 2068
rect 16878 2035 16912 2069
rect 16438 1953 16472 1987
rect 16555 1953 16589 1987
rect 17046 2041 17080 2075
rect 17142 2041 17176 2075
rect 16968 1930 17002 1964
<< locali >>
rect 18449 35209 18483 35226
rect 18993 35209 19027 35226
rect 18449 35197 18716 35209
rect 18483 35163 18554 35197
rect 18588 35163 18647 35197
rect 18681 35163 18716 35197
rect 18449 35151 18716 35163
rect 18848 35197 19027 35209
rect 18848 35163 18865 35197
rect 18899 35163 18993 35197
rect 18848 35151 19027 35163
rect 18449 35105 18483 35151
rect 18449 35015 18483 35071
rect 18517 35106 18959 35116
rect 18517 35099 18664 35106
rect 18698 35099 18959 35106
rect 18517 35065 18525 35099
rect 18559 35065 18596 35099
rect 18630 35070 18664 35099
rect 18630 35065 18667 35070
rect 18701 35069 18879 35099
rect 18701 35065 18714 35069
rect 18828 35065 18879 35069
rect 18913 35065 18959 35099
rect 18993 35105 19027 35151
rect 18517 35049 18714 35065
rect 18449 35013 18525 35015
rect 18483 34981 18525 35013
rect 18559 34981 18593 35015
rect 18627 34981 18661 35015
rect 18695 34981 18711 35015
rect 18483 34979 18711 34981
rect 18449 34972 18711 34979
rect 18745 35001 18761 35035
rect 18795 35001 18811 35035
rect 18993 35031 19027 35071
rect 18449 34921 18483 34972
rect 18745 34934 18811 35001
rect 18901 35015 19027 35031
rect 18901 34981 18917 35015
rect 18951 35013 19027 35015
rect 18951 34981 18993 35013
rect 18901 34979 18993 34981
rect 18901 34967 19027 34979
rect 18449 34829 18483 34887
rect 18521 34920 18811 34934
rect 18993 34921 19027 34967
rect 18521 34918 18891 34920
rect 18521 34884 18525 34918
rect 18559 34884 18593 34918
rect 18627 34886 18891 34918
rect 18925 34886 18941 34920
rect 18627 34884 18941 34886
rect 18521 34880 18941 34884
rect 18521 34868 18667 34880
rect 18887 34870 18941 34880
rect 18695 34832 18862 34846
rect 18695 34830 18949 34832
rect 18449 34737 18483 34795
rect 18526 34820 18949 34830
rect 18526 34816 18868 34820
rect 18906 34816 18949 34820
rect 18526 34814 18846 34816
rect 18526 34780 18531 34814
rect 18565 34780 18599 34814
rect 18633 34780 18667 34814
rect 18701 34808 18846 34814
rect 18701 34799 18721 34808
rect 18701 34780 18711 34799
rect 18837 34797 18846 34808
rect 18526 34764 18711 34780
rect 18845 34782 18846 34797
rect 18906 34814 18914 34816
rect 18948 34782 18949 34816
rect 18745 34740 18761 34774
rect 18795 34740 18811 34774
rect 18845 34766 18949 34782
rect 18993 34829 19027 34887
rect 18483 34703 18555 34730
rect 18449 34696 18555 34703
rect 18589 34696 18635 34730
rect 18669 34696 18685 34730
rect 18449 34645 18483 34696
rect 18745 34664 18811 34740
rect 18993 34737 19027 34795
rect 18871 34698 18887 34732
rect 18921 34703 18993 34732
rect 18921 34698 19027 34703
rect 18745 34662 18950 34664
rect 18449 34553 18483 34611
rect 18517 34648 18950 34662
rect 18517 34644 18848 34648
rect 18517 34610 18525 34644
rect 18559 34610 18596 34644
rect 18630 34610 18667 34644
rect 18701 34624 18848 34644
rect 18701 34610 18704 34624
rect 18517 34594 18704 34610
rect 18845 34614 18848 34624
rect 18882 34614 18916 34648
rect 18845 34598 18950 34614
rect 18993 34645 19027 34698
rect 18483 34520 18583 34547
rect 18483 34519 18533 34520
rect 18449 34486 18533 34519
rect 18567 34486 18583 34520
rect 18449 34484 18583 34486
rect 18629 34516 18704 34594
rect 18449 34461 18483 34484
rect 18629 34482 18645 34516
rect 18679 34482 18704 34516
rect 18745 34556 18761 34590
rect 18795 34556 18811 34590
rect 18745 34448 18811 34556
rect 18993 34553 19027 34611
rect 18887 34542 18993 34545
rect 18887 34508 18903 34542
rect 18937 34519 18993 34542
rect 18937 34508 19027 34519
rect 18887 34503 19027 34508
rect 18993 34461 19027 34503
rect 18449 34369 18483 34427
rect 18449 34277 18483 34335
rect 18543 34414 18937 34448
rect 18543 34321 18577 34414
rect 18611 34346 18645 34380
rect 18679 34367 18869 34380
rect 18679 34346 18687 34367
rect 18611 34333 18687 34346
rect 18721 34333 18869 34367
rect 18611 34321 18869 34333
rect 18611 34316 18819 34321
rect 18803 34287 18819 34316
rect 18853 34287 18869 34321
rect 18903 34344 18937 34414
rect 18903 34291 18937 34310
rect 18993 34369 19027 34427
rect 18543 34271 18577 34287
rect 18617 34280 18761 34282
rect 18617 34246 18619 34280
rect 18653 34278 18761 34280
rect 18653 34246 18711 34278
rect 18617 34244 18711 34246
rect 18745 34244 18761 34278
rect 18993 34277 19027 34335
rect 18449 34185 18483 34243
rect 18903 34241 18937 34257
rect 18517 34192 18533 34226
rect 18567 34210 18583 34226
rect 18567 34207 18903 34210
rect 18567 34192 18937 34207
rect 18517 34176 18937 34192
rect 18993 34185 19027 34243
rect 18449 34142 18483 34151
rect 18449 34108 18525 34142
rect 18559 34108 18593 34142
rect 18627 34108 18643 34142
rect 18695 34108 18711 34142
rect 18745 34108 18761 34142
rect 18449 34093 18483 34108
rect 18695 34074 18747 34108
rect 18797 34084 18857 34176
rect 18993 34140 19027 34151
rect 18449 34001 18483 34059
rect 18449 33909 18483 33967
rect 18449 33817 18483 33875
rect 18538 34040 18747 34074
rect 18791 34078 18857 34084
rect 18791 34044 18807 34078
rect 18841 34044 18857 34078
rect 18893 34122 19027 34140
rect 18893 34088 18909 34122
rect 18943 34093 19027 34122
rect 18943 34088 18993 34093
rect 18893 34066 18993 34088
rect 18538 33903 18572 34040
rect 18606 33968 18679 34006
rect 18713 34002 18747 34040
rect 18713 33968 18937 34002
rect 18606 33966 18645 33968
rect 18606 33932 18619 33966
rect 18653 33932 18863 33934
rect 18606 33900 18863 33932
rect 18538 33853 18572 33869
rect 18819 33879 18863 33900
rect 18666 33863 18785 33866
rect 18666 33829 18687 33863
rect 18721 33859 18785 33863
rect 18721 33829 18723 33859
rect 18666 33825 18723 33829
rect 18757 33825 18785 33859
rect 18853 33845 18863 33879
rect 18903 33923 18937 33968
rect 18903 33867 18937 33889
rect 18993 34001 19027 34059
rect 18993 33909 19027 33967
rect 18819 33829 18863 33845
rect 18666 33818 18785 33825
rect 18903 33812 18937 33828
rect 18449 33727 18483 33783
rect 18517 33777 18533 33811
rect 18567 33784 18628 33811
rect 18849 33784 18903 33795
rect 18567 33778 18903 33784
rect 18567 33777 18937 33778
rect 18517 33761 18937 33777
rect 18993 33817 19027 33875
rect 18602 33750 18875 33761
rect 18993 33727 19027 33783
rect 18449 33725 18525 33727
rect 18483 33693 18525 33725
rect 18559 33693 18575 33727
rect 18483 33691 18575 33693
rect 18449 33674 18575 33691
rect 18677 33682 18693 33716
rect 18727 33706 18867 33716
rect 18727 33682 18816 33706
rect 18449 33633 18483 33674
rect 18677 33670 18816 33682
rect 18852 33670 18867 33706
rect 18901 33693 18917 33727
rect 18951 33725 19027 33727
rect 18951 33693 18993 33725
rect 18901 33691 18993 33693
rect 18901 33677 19027 33691
rect 18677 33660 18867 33670
rect 18993 33633 19027 33677
rect 18449 33555 18483 33599
rect 18517 33625 18941 33626
rect 18517 33623 18687 33625
rect 18517 33589 18533 33623
rect 18567 33589 18601 33623
rect 18635 33591 18687 33623
rect 18721 33623 18941 33625
rect 18721 33591 18891 33623
rect 18635 33589 18891 33591
rect 18925 33589 18941 33623
rect 18993 33555 19027 33599
rect 18449 33541 18583 33555
rect 18483 33539 18583 33541
rect 18483 33507 18549 33539
rect 18449 33505 18549 33507
rect 18449 33489 18583 33505
rect 18617 33546 18746 33554
rect 18617 33512 18619 33546
rect 18653 33520 18746 33546
rect 18780 33520 18883 33554
rect 18653 33512 18883 33520
rect 18617 33508 18883 33512
rect 18449 33449 18483 33489
rect 18617 33455 18651 33508
rect 18517 33421 18533 33455
rect 18567 33421 18601 33455
rect 18635 33421 18651 33455
rect 18685 33456 18815 33474
rect 18449 33386 18483 33415
rect 18685 33420 18748 33456
rect 18784 33452 18815 33456
rect 18685 33418 18761 33420
rect 18795 33418 18815 33452
rect 18849 33455 18883 33508
rect 18917 33541 19027 33555
rect 18917 33539 18993 33541
rect 18951 33507 18993 33539
rect 18951 33505 19027 33507
rect 18917 33489 19027 33505
rect 18849 33421 18891 33455
rect 18925 33421 18941 33455
rect 18993 33449 19027 33489
rect 18685 33404 18815 33418
rect 18993 33386 19027 33415
rect 18457 32903 18491 32920
rect 19001 32903 19035 32920
rect 18457 32891 18724 32903
rect 18491 32857 18562 32891
rect 18596 32857 18655 32891
rect 18689 32857 18724 32891
rect 18457 32845 18724 32857
rect 18856 32891 19035 32903
rect 18856 32857 18873 32891
rect 18907 32857 19001 32891
rect 18856 32845 19035 32857
rect 18457 32799 18491 32845
rect 18457 32709 18491 32765
rect 18525 32800 18967 32810
rect 18525 32793 18672 32800
rect 18706 32793 18967 32800
rect 18525 32759 18533 32793
rect 18567 32759 18604 32793
rect 18638 32764 18672 32793
rect 18638 32759 18675 32764
rect 18709 32763 18887 32793
rect 18709 32759 18722 32763
rect 18836 32759 18887 32763
rect 18921 32759 18967 32793
rect 19001 32799 19035 32845
rect 18525 32743 18722 32759
rect 18457 32707 18533 32709
rect 18491 32675 18533 32707
rect 18567 32675 18601 32709
rect 18635 32675 18669 32709
rect 18703 32675 18719 32709
rect 18491 32673 18719 32675
rect 18457 32666 18719 32673
rect 18753 32695 18769 32729
rect 18803 32695 18819 32729
rect 19001 32725 19035 32765
rect 18457 32615 18491 32666
rect 18753 32628 18819 32695
rect 18909 32709 19035 32725
rect 18909 32675 18925 32709
rect 18959 32707 19035 32709
rect 18959 32675 19001 32707
rect 18909 32673 19001 32675
rect 18909 32661 19035 32673
rect 18457 32523 18491 32581
rect 18529 32614 18819 32628
rect 19001 32615 19035 32661
rect 18529 32612 18899 32614
rect 18529 32578 18533 32612
rect 18567 32578 18601 32612
rect 18635 32580 18899 32612
rect 18933 32580 18949 32614
rect 18635 32578 18949 32580
rect 18529 32574 18949 32578
rect 18529 32562 18675 32574
rect 18895 32564 18949 32574
rect 18703 32526 18870 32540
rect 18703 32524 18957 32526
rect 18457 32431 18491 32489
rect 18534 32510 18957 32524
rect 18534 32508 18854 32510
rect 18534 32474 18539 32508
rect 18573 32474 18607 32508
rect 18641 32474 18675 32508
rect 18709 32502 18854 32508
rect 18709 32493 18729 32502
rect 18709 32474 18719 32493
rect 18845 32491 18854 32502
rect 18534 32458 18719 32474
rect 18853 32476 18854 32491
rect 18888 32476 18922 32510
rect 18956 32476 18957 32510
rect 18753 32434 18769 32468
rect 18803 32434 18819 32468
rect 18853 32460 18957 32476
rect 19001 32523 19035 32581
rect 18491 32397 18563 32424
rect 18457 32390 18563 32397
rect 18597 32390 18643 32424
rect 18677 32390 18693 32424
rect 18457 32339 18491 32390
rect 18753 32358 18819 32434
rect 19001 32431 19035 32489
rect 18879 32392 18895 32426
rect 18929 32397 19001 32426
rect 18929 32392 19035 32397
rect 18753 32356 18958 32358
rect 18457 32247 18491 32305
rect 18525 32342 18958 32356
rect 18525 32338 18856 32342
rect 18525 32304 18533 32338
rect 18567 32304 18604 32338
rect 18638 32304 18675 32338
rect 18709 32318 18856 32338
rect 18709 32304 18712 32318
rect 18525 32288 18712 32304
rect 18853 32308 18856 32318
rect 18890 32308 18924 32342
rect 18853 32292 18958 32308
rect 19001 32339 19035 32392
rect 18491 32214 18591 32241
rect 18491 32213 18541 32214
rect 18457 32180 18541 32213
rect 18575 32180 18591 32214
rect 18457 32178 18591 32180
rect 18637 32210 18712 32288
rect 18457 32155 18491 32178
rect 18637 32176 18653 32210
rect 18687 32176 18712 32210
rect 18753 32250 18769 32284
rect 18803 32250 18819 32284
rect 18753 32142 18819 32250
rect 19001 32247 19035 32305
rect 18895 32236 19001 32239
rect 18895 32202 18911 32236
rect 18945 32213 19001 32236
rect 18945 32202 19035 32213
rect 18895 32197 19035 32202
rect 19001 32155 19035 32197
rect 18457 32063 18491 32121
rect 18457 31971 18491 32029
rect 18551 32108 18945 32142
rect 18551 32015 18585 32108
rect 18619 32040 18653 32074
rect 18687 32061 18877 32074
rect 18687 32040 18695 32061
rect 18619 32027 18695 32040
rect 18729 32027 18877 32061
rect 18619 32015 18877 32027
rect 18619 32010 18827 32015
rect 18811 31981 18827 32010
rect 18861 31981 18877 32015
rect 18911 32038 18945 32108
rect 18911 31985 18945 32004
rect 19001 32063 19035 32121
rect 18551 31965 18585 31981
rect 18625 31974 18769 31976
rect 18625 31940 18627 31974
rect 18661 31972 18769 31974
rect 18661 31940 18719 31972
rect 18625 31938 18719 31940
rect 18753 31938 18769 31972
rect 19001 31971 19035 32029
rect 18457 31879 18491 31937
rect 18911 31935 18945 31951
rect 18525 31886 18541 31920
rect 18575 31904 18591 31920
rect 18575 31901 18911 31904
rect 18575 31886 18945 31901
rect 18525 31870 18945 31886
rect 19001 31879 19035 31937
rect 18457 31836 18491 31845
rect 18457 31802 18533 31836
rect 18567 31802 18601 31836
rect 18635 31802 18651 31836
rect 18703 31802 18719 31836
rect 18753 31802 18769 31836
rect 18457 31787 18491 31802
rect 18703 31768 18755 31802
rect 18805 31778 18865 31870
rect 19001 31834 19035 31845
rect 18457 31695 18491 31753
rect 18457 31603 18491 31661
rect 18457 31511 18491 31569
rect 18546 31734 18755 31768
rect 18799 31772 18865 31778
rect 18799 31738 18815 31772
rect 18849 31738 18865 31772
rect 18901 31816 19035 31834
rect 18901 31782 18917 31816
rect 18951 31787 19035 31816
rect 18951 31782 19001 31787
rect 18901 31760 19001 31782
rect 18546 31597 18580 31734
rect 18614 31662 18687 31700
rect 18721 31696 18755 31734
rect 18721 31662 18945 31696
rect 18614 31660 18653 31662
rect 18614 31626 18627 31660
rect 18661 31626 18871 31628
rect 18614 31594 18871 31626
rect 18546 31547 18580 31563
rect 18827 31573 18871 31594
rect 18674 31557 18793 31560
rect 18674 31523 18695 31557
rect 18729 31553 18793 31557
rect 18729 31523 18731 31553
rect 18674 31519 18731 31523
rect 18765 31519 18793 31553
rect 18861 31539 18871 31573
rect 18911 31617 18945 31662
rect 18911 31561 18945 31583
rect 19001 31695 19035 31753
rect 19001 31603 19035 31661
rect 18827 31523 18871 31539
rect 18674 31512 18793 31519
rect 18911 31506 18945 31522
rect 18457 31421 18491 31477
rect 18525 31471 18541 31505
rect 18575 31478 18636 31505
rect 18857 31478 18911 31489
rect 18575 31472 18911 31478
rect 18575 31471 18945 31472
rect 18525 31455 18945 31471
rect 19001 31511 19035 31569
rect 18610 31444 18883 31455
rect 19001 31421 19035 31477
rect 18457 31419 18533 31421
rect 18491 31387 18533 31419
rect 18567 31387 18583 31421
rect 18491 31385 18583 31387
rect 18457 31368 18583 31385
rect 18685 31376 18701 31410
rect 18735 31400 18875 31410
rect 18735 31376 18824 31400
rect 18457 31327 18491 31368
rect 18685 31364 18824 31376
rect 18860 31364 18875 31400
rect 18909 31387 18925 31421
rect 18959 31419 19035 31421
rect 18959 31387 19001 31419
rect 18909 31385 19001 31387
rect 18909 31371 19035 31385
rect 18685 31354 18875 31364
rect 19001 31327 19035 31371
rect 18457 31249 18491 31293
rect 18525 31319 18949 31320
rect 18525 31317 18695 31319
rect 18525 31283 18541 31317
rect 18575 31283 18609 31317
rect 18643 31285 18695 31317
rect 18729 31317 18949 31319
rect 18729 31285 18899 31317
rect 18643 31283 18899 31285
rect 18933 31283 18949 31317
rect 19001 31249 19035 31293
rect 18457 31235 18591 31249
rect 18491 31233 18591 31235
rect 18491 31201 18557 31233
rect 18457 31199 18557 31201
rect 18457 31183 18591 31199
rect 18625 31240 18754 31248
rect 18625 31206 18627 31240
rect 18661 31214 18754 31240
rect 18788 31214 18891 31248
rect 18661 31206 18891 31214
rect 18625 31202 18891 31206
rect 18457 31143 18491 31183
rect 18625 31149 18659 31202
rect 18525 31115 18541 31149
rect 18575 31115 18609 31149
rect 18643 31115 18659 31149
rect 18693 31150 18823 31168
rect 18457 31080 18491 31109
rect 18693 31114 18756 31150
rect 18792 31146 18823 31150
rect 18693 31112 18769 31114
rect 18803 31112 18823 31146
rect 18857 31149 18891 31202
rect 18925 31235 19035 31249
rect 18925 31233 19001 31235
rect 18959 31201 19001 31233
rect 18959 31199 19035 31201
rect 18925 31183 19035 31199
rect 18857 31115 18899 31149
rect 18933 31115 18949 31149
rect 19001 31143 19035 31183
rect 18693 31098 18823 31112
rect 19001 31080 19035 31109
rect 18465 30689 18499 30706
rect 19009 30689 19043 30706
rect 18465 30677 18732 30689
rect 18499 30643 18570 30677
rect 18604 30643 18663 30677
rect 18697 30643 18732 30677
rect 18465 30631 18732 30643
rect 18864 30677 19043 30689
rect 18864 30643 18881 30677
rect 18915 30643 19009 30677
rect 18864 30631 19043 30643
rect 18465 30585 18499 30631
rect 18465 30495 18499 30551
rect 18533 30586 18975 30596
rect 18533 30579 18680 30586
rect 18714 30579 18975 30586
rect 18533 30545 18541 30579
rect 18575 30545 18612 30579
rect 18646 30550 18680 30579
rect 18646 30545 18683 30550
rect 18717 30549 18895 30579
rect 18717 30545 18730 30549
rect 18844 30545 18895 30549
rect 18929 30545 18975 30579
rect 19009 30585 19043 30631
rect 18533 30529 18730 30545
rect 18465 30493 18541 30495
rect 18499 30461 18541 30493
rect 18575 30461 18609 30495
rect 18643 30461 18677 30495
rect 18711 30461 18727 30495
rect 18499 30459 18727 30461
rect 18465 30452 18727 30459
rect 18761 30481 18777 30515
rect 18811 30481 18827 30515
rect 19009 30511 19043 30551
rect 18465 30401 18499 30452
rect 18761 30414 18827 30481
rect 18917 30495 19043 30511
rect 18917 30461 18933 30495
rect 18967 30493 19043 30495
rect 18967 30461 19009 30493
rect 18917 30459 19009 30461
rect 18917 30447 19043 30459
rect 18465 30309 18499 30367
rect 18537 30400 18827 30414
rect 19009 30401 19043 30447
rect 18537 30398 18907 30400
rect 18537 30364 18541 30398
rect 18575 30364 18609 30398
rect 18643 30366 18907 30398
rect 18941 30366 18957 30400
rect 18643 30364 18957 30366
rect 18537 30360 18957 30364
rect 18537 30348 18683 30360
rect 18903 30350 18957 30360
rect 18711 30312 18878 30326
rect 18711 30310 18965 30312
rect 18465 30217 18499 30275
rect 18542 30296 18965 30310
rect 18542 30294 18862 30296
rect 18542 30260 18547 30294
rect 18581 30260 18615 30294
rect 18649 30260 18683 30294
rect 18717 30288 18862 30294
rect 18717 30279 18737 30288
rect 18717 30260 18727 30279
rect 18853 30277 18862 30288
rect 18542 30244 18727 30260
rect 18861 30262 18862 30277
rect 18896 30262 18930 30296
rect 18964 30262 18965 30296
rect 18761 30220 18777 30254
rect 18811 30220 18827 30254
rect 18861 30246 18965 30262
rect 19009 30309 19043 30367
rect 18499 30183 18571 30210
rect 18465 30176 18571 30183
rect 18605 30176 18651 30210
rect 18685 30176 18701 30210
rect 18465 30125 18499 30176
rect 18761 30144 18827 30220
rect 19009 30217 19043 30275
rect 18887 30178 18903 30212
rect 18937 30183 19009 30212
rect 18937 30178 19043 30183
rect 18761 30142 18966 30144
rect 18465 30033 18499 30091
rect 18533 30128 18966 30142
rect 18533 30124 18864 30128
rect 18533 30090 18541 30124
rect 18575 30090 18612 30124
rect 18646 30090 18683 30124
rect 18717 30104 18864 30124
rect 18717 30090 18720 30104
rect 18533 30074 18720 30090
rect 18861 30094 18864 30104
rect 18898 30094 18932 30128
rect 18861 30078 18966 30094
rect 19009 30125 19043 30178
rect 18499 30000 18599 30027
rect 18499 29999 18549 30000
rect 18465 29966 18549 29999
rect 18583 29966 18599 30000
rect 18465 29964 18599 29966
rect 18645 29996 18720 30074
rect 18465 29941 18499 29964
rect 18645 29962 18661 29996
rect 18695 29962 18720 29996
rect 18761 30036 18777 30070
rect 18811 30036 18827 30070
rect 18761 29928 18827 30036
rect 19009 30033 19043 30091
rect 18903 30022 19009 30025
rect 18903 29988 18919 30022
rect 18953 29999 19009 30022
rect 18953 29988 19043 29999
rect 18903 29983 19043 29988
rect 19009 29941 19043 29983
rect 18465 29849 18499 29907
rect 18465 29757 18499 29815
rect 18559 29894 18953 29928
rect 18559 29801 18593 29894
rect 18627 29826 18661 29860
rect 18695 29847 18885 29860
rect 18695 29826 18703 29847
rect 18627 29813 18703 29826
rect 18737 29813 18885 29847
rect 18627 29801 18885 29813
rect 18627 29796 18835 29801
rect 18819 29767 18835 29796
rect 18869 29767 18885 29801
rect 18919 29824 18953 29894
rect 18919 29771 18953 29790
rect 19009 29849 19043 29907
rect 18559 29751 18593 29767
rect 18633 29760 18777 29762
rect 18633 29726 18635 29760
rect 18669 29758 18777 29760
rect 18669 29726 18727 29758
rect 18633 29724 18727 29726
rect 18761 29724 18777 29758
rect 19009 29757 19043 29815
rect 18465 29665 18499 29723
rect 18919 29721 18953 29737
rect 18533 29672 18549 29706
rect 18583 29690 18599 29706
rect 18583 29687 18919 29690
rect 18583 29672 18953 29687
rect 18533 29656 18953 29672
rect 19009 29665 19043 29723
rect 18465 29622 18499 29631
rect 18465 29588 18541 29622
rect 18575 29588 18609 29622
rect 18643 29588 18659 29622
rect 18711 29588 18727 29622
rect 18761 29588 18777 29622
rect 18465 29573 18499 29588
rect 18711 29554 18763 29588
rect 18813 29564 18873 29656
rect 19009 29620 19043 29631
rect 18465 29481 18499 29539
rect 18465 29389 18499 29447
rect 18465 29297 18499 29355
rect 18554 29520 18763 29554
rect 18807 29558 18873 29564
rect 18807 29524 18823 29558
rect 18857 29524 18873 29558
rect 18909 29602 19043 29620
rect 18909 29568 18925 29602
rect 18959 29573 19043 29602
rect 18959 29568 19009 29573
rect 18909 29546 19009 29568
rect 18554 29383 18588 29520
rect 18622 29448 18695 29486
rect 18729 29482 18763 29520
rect 18729 29448 18953 29482
rect 18622 29446 18661 29448
rect 18622 29412 18635 29446
rect 18669 29412 18879 29414
rect 18622 29380 18879 29412
rect 18554 29333 18588 29349
rect 18835 29359 18879 29380
rect 18682 29343 18801 29346
rect 18682 29309 18703 29343
rect 18737 29339 18801 29343
rect 18737 29309 18739 29339
rect 18682 29305 18739 29309
rect 18773 29305 18801 29339
rect 18869 29325 18879 29359
rect 18919 29403 18953 29448
rect 18919 29347 18953 29369
rect 19009 29481 19043 29539
rect 19009 29389 19043 29447
rect 18835 29309 18879 29325
rect 18682 29298 18801 29305
rect 18919 29292 18953 29308
rect 18465 29207 18499 29263
rect 18533 29257 18549 29291
rect 18583 29264 18644 29291
rect 18865 29264 18919 29275
rect 18583 29258 18919 29264
rect 18583 29257 18953 29258
rect 18533 29241 18953 29257
rect 19009 29297 19043 29355
rect 18618 29230 18891 29241
rect 19009 29207 19043 29263
rect 18465 29205 18541 29207
rect 18499 29173 18541 29205
rect 18575 29173 18591 29207
rect 18499 29171 18591 29173
rect 18465 29154 18591 29171
rect 18693 29162 18709 29196
rect 18743 29186 18883 29196
rect 18743 29162 18832 29186
rect 18465 29113 18499 29154
rect 18693 29150 18832 29162
rect 18868 29150 18883 29186
rect 18917 29173 18933 29207
rect 18967 29205 19043 29207
rect 18967 29173 19009 29205
rect 18917 29171 19009 29173
rect 18917 29157 19043 29171
rect 18693 29140 18883 29150
rect 19009 29113 19043 29157
rect 18465 29035 18499 29079
rect 18533 29105 18957 29106
rect 18533 29103 18703 29105
rect 18533 29069 18549 29103
rect 18583 29069 18617 29103
rect 18651 29071 18703 29103
rect 18737 29103 18957 29105
rect 18737 29071 18907 29103
rect 18651 29069 18907 29071
rect 18941 29069 18957 29103
rect 19009 29035 19043 29079
rect 18465 29021 18599 29035
rect 18499 29019 18599 29021
rect 18499 28987 18565 29019
rect 18465 28985 18565 28987
rect 18465 28969 18599 28985
rect 18633 29026 18762 29034
rect 18633 28992 18635 29026
rect 18669 29000 18762 29026
rect 18796 29000 18899 29034
rect 18669 28992 18899 29000
rect 18633 28988 18899 28992
rect 18465 28929 18499 28969
rect 18633 28935 18667 28988
rect 18533 28901 18549 28935
rect 18583 28901 18617 28935
rect 18651 28901 18667 28935
rect 18701 28936 18831 28954
rect 18465 28866 18499 28895
rect 18701 28900 18764 28936
rect 18800 28932 18831 28936
rect 18701 28898 18777 28900
rect 18811 28898 18831 28932
rect 18865 28935 18899 28988
rect 18933 29021 19043 29035
rect 18933 29019 19009 29021
rect 18967 28987 19009 29019
rect 18967 28985 19043 28987
rect 18933 28969 19043 28985
rect 18865 28901 18907 28935
rect 18941 28901 18957 28935
rect 19009 28929 19043 28969
rect 18701 28884 18831 28898
rect 19009 28866 19043 28895
rect 18447 28489 18481 28506
rect 18991 28489 19025 28506
rect 18447 28477 18714 28489
rect 18481 28443 18552 28477
rect 18586 28443 18645 28477
rect 18679 28443 18714 28477
rect 18447 28431 18714 28443
rect 18846 28477 19025 28489
rect 18846 28443 18863 28477
rect 18897 28443 18991 28477
rect 18846 28431 19025 28443
rect 18447 28385 18481 28431
rect 18447 28295 18481 28351
rect 18515 28386 18957 28396
rect 18515 28379 18662 28386
rect 18696 28379 18957 28386
rect 18515 28345 18523 28379
rect 18557 28345 18594 28379
rect 18628 28350 18662 28379
rect 18628 28345 18665 28350
rect 18699 28349 18877 28379
rect 18699 28345 18712 28349
rect 18826 28345 18877 28349
rect 18911 28345 18957 28379
rect 18991 28385 19025 28431
rect 18515 28329 18712 28345
rect 18447 28293 18523 28295
rect 18481 28261 18523 28293
rect 18557 28261 18591 28295
rect 18625 28261 18659 28295
rect 18693 28261 18709 28295
rect 18481 28259 18709 28261
rect 18447 28252 18709 28259
rect 18743 28281 18759 28315
rect 18793 28281 18809 28315
rect 18991 28311 19025 28351
rect 18447 28201 18481 28252
rect 18743 28214 18809 28281
rect 18899 28295 19025 28311
rect 18899 28261 18915 28295
rect 18949 28293 19025 28295
rect 18949 28261 18991 28293
rect 18899 28259 18991 28261
rect 18899 28247 19025 28259
rect 18447 28109 18481 28167
rect 18519 28200 18809 28214
rect 18991 28201 19025 28247
rect 18519 28198 18889 28200
rect 18519 28164 18523 28198
rect 18557 28164 18591 28198
rect 18625 28166 18889 28198
rect 18923 28166 18939 28200
rect 18625 28164 18939 28166
rect 18519 28160 18939 28164
rect 18519 28148 18665 28160
rect 18885 28150 18939 28160
rect 18693 28112 18860 28126
rect 18693 28110 18947 28112
rect 18447 28017 18481 28075
rect 18524 28096 18947 28110
rect 18524 28094 18844 28096
rect 18524 28060 18529 28094
rect 18563 28060 18597 28094
rect 18631 28060 18665 28094
rect 18699 28088 18844 28094
rect 18699 28079 18719 28088
rect 18699 28060 18709 28079
rect 18835 28077 18844 28088
rect 18524 28044 18709 28060
rect 18843 28062 18844 28077
rect 18878 28062 18912 28096
rect 18946 28062 18947 28096
rect 18743 28020 18759 28054
rect 18793 28020 18809 28054
rect 18843 28046 18947 28062
rect 18991 28109 19025 28167
rect 18481 27983 18553 28010
rect 18447 27976 18553 27983
rect 18587 27976 18633 28010
rect 18667 27976 18683 28010
rect 18447 27925 18481 27976
rect 18743 27944 18809 28020
rect 18991 28017 19025 28075
rect 18869 27978 18885 28012
rect 18919 27983 18991 28012
rect 18919 27978 19025 27983
rect 18743 27942 18948 27944
rect 18447 27833 18481 27891
rect 18515 27928 18948 27942
rect 18515 27924 18846 27928
rect 18515 27890 18523 27924
rect 18557 27890 18594 27924
rect 18628 27890 18665 27924
rect 18699 27904 18846 27924
rect 18699 27890 18702 27904
rect 18515 27874 18702 27890
rect 18843 27894 18846 27904
rect 18880 27894 18914 27928
rect 18843 27878 18948 27894
rect 18991 27925 19025 27978
rect 18481 27800 18581 27827
rect 18481 27799 18531 27800
rect 18447 27766 18531 27799
rect 18565 27766 18581 27800
rect 18447 27764 18581 27766
rect 18627 27796 18702 27874
rect 18447 27741 18481 27764
rect 18627 27762 18643 27796
rect 18677 27762 18702 27796
rect 18743 27836 18759 27870
rect 18793 27836 18809 27870
rect 18743 27728 18809 27836
rect 18991 27833 19025 27891
rect 18885 27822 18991 27825
rect 18885 27788 18901 27822
rect 18935 27799 18991 27822
rect 18935 27788 19025 27799
rect 18885 27783 19025 27788
rect 18991 27741 19025 27783
rect 18447 27649 18481 27707
rect 18447 27557 18481 27615
rect 18541 27694 18935 27728
rect 18541 27601 18575 27694
rect 18609 27626 18643 27660
rect 18677 27647 18867 27660
rect 18677 27626 18685 27647
rect 18609 27613 18685 27626
rect 18719 27613 18867 27647
rect 18609 27601 18867 27613
rect 18609 27596 18817 27601
rect 18801 27567 18817 27596
rect 18851 27567 18867 27601
rect 18901 27624 18935 27694
rect 18901 27571 18935 27590
rect 18991 27649 19025 27707
rect 18541 27551 18575 27567
rect 18615 27560 18759 27562
rect 18615 27526 18617 27560
rect 18651 27558 18759 27560
rect 18651 27526 18709 27558
rect 18615 27524 18709 27526
rect 18743 27524 18759 27558
rect 18991 27557 19025 27615
rect 18447 27465 18481 27523
rect 18901 27521 18935 27537
rect 18515 27472 18531 27506
rect 18565 27490 18581 27506
rect 18565 27487 18901 27490
rect 18565 27472 18935 27487
rect 18515 27456 18935 27472
rect 18991 27465 19025 27523
rect 18447 27422 18481 27431
rect 18447 27388 18523 27422
rect 18557 27388 18591 27422
rect 18625 27388 18641 27422
rect 18693 27388 18709 27422
rect 18743 27388 18759 27422
rect 18447 27373 18481 27388
rect 18693 27354 18745 27388
rect 18795 27364 18855 27456
rect 18991 27420 19025 27431
rect 18447 27281 18481 27339
rect 18447 27189 18481 27247
rect 18447 27097 18481 27155
rect 18536 27320 18745 27354
rect 18789 27358 18855 27364
rect 18789 27324 18805 27358
rect 18839 27324 18855 27358
rect 18891 27402 19025 27420
rect 18891 27368 18907 27402
rect 18941 27373 19025 27402
rect 18941 27368 18991 27373
rect 18891 27346 18991 27368
rect 18536 27183 18570 27320
rect 18604 27248 18677 27286
rect 18711 27282 18745 27320
rect 18711 27248 18935 27282
rect 18604 27246 18643 27248
rect 18604 27212 18617 27246
rect 18651 27212 18861 27214
rect 18604 27180 18861 27212
rect 18536 27133 18570 27149
rect 18817 27159 18861 27180
rect 18664 27143 18783 27146
rect 18664 27109 18685 27143
rect 18719 27139 18783 27143
rect 18719 27109 18721 27139
rect 18664 27105 18721 27109
rect 18755 27105 18783 27139
rect 18851 27125 18861 27159
rect 18901 27203 18935 27248
rect 18901 27147 18935 27169
rect 18991 27281 19025 27339
rect 18991 27189 19025 27247
rect 18817 27109 18861 27125
rect 18664 27098 18783 27105
rect 18901 27092 18935 27108
rect 18447 27007 18481 27063
rect 18515 27057 18531 27091
rect 18565 27064 18626 27091
rect 18847 27064 18901 27075
rect 18565 27058 18901 27064
rect 18565 27057 18935 27058
rect 18515 27041 18935 27057
rect 18991 27097 19025 27155
rect 18600 27030 18873 27041
rect 18991 27007 19025 27063
rect 18447 27005 18523 27007
rect 18481 26973 18523 27005
rect 18557 26973 18573 27007
rect 18481 26971 18573 26973
rect 18447 26954 18573 26971
rect 18675 26962 18691 26996
rect 18725 26986 18865 26996
rect 18725 26962 18814 26986
rect 18447 26913 18481 26954
rect 18675 26950 18814 26962
rect 18850 26950 18865 26986
rect 18899 26973 18915 27007
rect 18949 27005 19025 27007
rect 18949 26973 18991 27005
rect 18899 26971 18991 26973
rect 18899 26957 19025 26971
rect 18675 26940 18865 26950
rect 18991 26913 19025 26957
rect 18447 26835 18481 26879
rect 18515 26905 18939 26906
rect 18515 26903 18685 26905
rect 18515 26869 18531 26903
rect 18565 26869 18599 26903
rect 18633 26871 18685 26903
rect 18719 26903 18939 26905
rect 18719 26871 18889 26903
rect 18633 26869 18889 26871
rect 18923 26869 18939 26903
rect 18991 26835 19025 26879
rect 18447 26821 18581 26835
rect 18481 26819 18581 26821
rect 18481 26787 18547 26819
rect 18447 26785 18547 26787
rect 18447 26769 18581 26785
rect 18615 26826 18744 26834
rect 18615 26792 18617 26826
rect 18651 26800 18744 26826
rect 18778 26800 18881 26834
rect 18651 26792 18881 26800
rect 18615 26788 18881 26792
rect 18447 26729 18481 26769
rect 18615 26735 18649 26788
rect 18515 26701 18531 26735
rect 18565 26701 18599 26735
rect 18633 26701 18649 26735
rect 18683 26736 18813 26754
rect 18447 26666 18481 26695
rect 18683 26700 18746 26736
rect 18782 26732 18813 26736
rect 18683 26698 18759 26700
rect 18793 26698 18813 26732
rect 18847 26735 18881 26788
rect 18915 26821 19025 26835
rect 18915 26819 18991 26821
rect 18949 26787 18991 26819
rect 18949 26785 19025 26787
rect 18915 26769 19025 26785
rect 18847 26701 18889 26735
rect 18923 26701 18939 26735
rect 18991 26729 19025 26769
rect 18683 26684 18813 26698
rect 18991 26666 19025 26695
rect 18455 26275 18489 26292
rect 18999 26275 19033 26292
rect 18455 26263 18722 26275
rect 18489 26229 18560 26263
rect 18594 26229 18653 26263
rect 18687 26229 18722 26263
rect 18455 26217 18722 26229
rect 18854 26263 19033 26275
rect 18854 26229 18871 26263
rect 18905 26229 18999 26263
rect 18854 26217 19033 26229
rect 18455 26171 18489 26217
rect 18455 26081 18489 26137
rect 18523 26172 18965 26182
rect 18523 26165 18670 26172
rect 18704 26165 18965 26172
rect 18523 26131 18531 26165
rect 18565 26131 18602 26165
rect 18636 26136 18670 26165
rect 18636 26131 18673 26136
rect 18707 26135 18885 26165
rect 18707 26131 18720 26135
rect 18834 26131 18885 26135
rect 18919 26131 18965 26165
rect 18999 26171 19033 26217
rect 18523 26115 18720 26131
rect 18455 26079 18531 26081
rect 18489 26047 18531 26079
rect 18565 26047 18599 26081
rect 18633 26047 18667 26081
rect 18701 26047 18717 26081
rect 18489 26045 18717 26047
rect 18455 26038 18717 26045
rect 18751 26067 18767 26101
rect 18801 26067 18817 26101
rect 18999 26097 19033 26137
rect 18455 25987 18489 26038
rect 18751 26000 18817 26067
rect 18907 26081 19033 26097
rect 18907 26047 18923 26081
rect 18957 26079 19033 26081
rect 18957 26047 18999 26079
rect 18907 26045 18999 26047
rect 18907 26033 19033 26045
rect 18455 25895 18489 25953
rect 18527 25986 18817 26000
rect 18999 25987 19033 26033
rect 18527 25984 18897 25986
rect 18527 25950 18531 25984
rect 18565 25950 18599 25984
rect 18633 25952 18897 25984
rect 18931 25952 18947 25986
rect 18633 25950 18947 25952
rect 18527 25946 18947 25950
rect 18527 25934 18673 25946
rect 18893 25936 18947 25946
rect 18701 25898 18868 25912
rect 18701 25896 18955 25898
rect 18455 25803 18489 25861
rect 18532 25882 18955 25896
rect 18532 25880 18852 25882
rect 18532 25846 18537 25880
rect 18571 25846 18605 25880
rect 18639 25846 18673 25880
rect 18707 25874 18852 25880
rect 18707 25865 18727 25874
rect 18707 25846 18717 25865
rect 18843 25863 18852 25874
rect 18532 25830 18717 25846
rect 18851 25848 18852 25863
rect 18886 25848 18920 25882
rect 18954 25848 18955 25882
rect 18751 25806 18767 25840
rect 18801 25806 18817 25840
rect 18851 25832 18955 25848
rect 18999 25895 19033 25953
rect 18489 25769 18561 25796
rect 18455 25762 18561 25769
rect 18595 25762 18641 25796
rect 18675 25762 18691 25796
rect 18455 25711 18489 25762
rect 18751 25730 18817 25806
rect 18999 25803 19033 25861
rect 18877 25764 18893 25798
rect 18927 25769 18999 25798
rect 18927 25764 19033 25769
rect 18751 25728 18956 25730
rect 18455 25619 18489 25677
rect 18523 25714 18956 25728
rect 18523 25710 18854 25714
rect 18523 25676 18531 25710
rect 18565 25676 18602 25710
rect 18636 25676 18673 25710
rect 18707 25690 18854 25710
rect 18707 25676 18710 25690
rect 18523 25660 18710 25676
rect 18851 25680 18854 25690
rect 18888 25680 18922 25714
rect 18851 25664 18956 25680
rect 18999 25711 19033 25764
rect 18489 25586 18589 25613
rect 18489 25585 18539 25586
rect 18455 25552 18539 25585
rect 18573 25552 18589 25586
rect 18455 25550 18589 25552
rect 18635 25582 18710 25660
rect 18455 25527 18489 25550
rect 18635 25548 18651 25582
rect 18685 25548 18710 25582
rect 18751 25622 18767 25656
rect 18801 25622 18817 25656
rect 18751 25514 18817 25622
rect 18999 25619 19033 25677
rect 18893 25608 18999 25611
rect 18893 25574 18909 25608
rect 18943 25585 18999 25608
rect 18943 25574 19033 25585
rect 18893 25569 19033 25574
rect 18999 25527 19033 25569
rect 18455 25435 18489 25493
rect 18455 25343 18489 25401
rect 18549 25480 18943 25514
rect 18549 25387 18583 25480
rect 18617 25412 18651 25446
rect 18685 25433 18875 25446
rect 18685 25412 18693 25433
rect 18617 25399 18693 25412
rect 18727 25399 18875 25433
rect 18617 25387 18875 25399
rect 18617 25382 18825 25387
rect 18809 25353 18825 25382
rect 18859 25353 18875 25387
rect 18909 25410 18943 25480
rect 18909 25357 18943 25376
rect 18999 25435 19033 25493
rect 18549 25337 18583 25353
rect 18623 25346 18767 25348
rect 18623 25312 18625 25346
rect 18659 25344 18767 25346
rect 18659 25312 18717 25344
rect 18623 25310 18717 25312
rect 18751 25310 18767 25344
rect 18999 25343 19033 25401
rect 18455 25251 18489 25309
rect 18909 25307 18943 25323
rect 18523 25258 18539 25292
rect 18573 25276 18589 25292
rect 18573 25273 18909 25276
rect 18573 25258 18943 25273
rect 18523 25242 18943 25258
rect 18999 25251 19033 25309
rect 18455 25208 18489 25217
rect 18455 25174 18531 25208
rect 18565 25174 18599 25208
rect 18633 25174 18649 25208
rect 18701 25174 18717 25208
rect 18751 25174 18767 25208
rect 18455 25159 18489 25174
rect 18701 25140 18753 25174
rect 18803 25150 18863 25242
rect 18999 25206 19033 25217
rect 18455 25067 18489 25125
rect 18455 24975 18489 25033
rect 18455 24883 18489 24941
rect 18544 25106 18753 25140
rect 18797 25144 18863 25150
rect 18797 25110 18813 25144
rect 18847 25110 18863 25144
rect 18899 25188 19033 25206
rect 18899 25154 18915 25188
rect 18949 25159 19033 25188
rect 18949 25154 18999 25159
rect 18899 25132 18999 25154
rect 18544 24969 18578 25106
rect 18612 25034 18685 25072
rect 18719 25068 18753 25106
rect 18719 25034 18943 25068
rect 18612 25032 18651 25034
rect 18612 24998 18625 25032
rect 18659 24998 18869 25000
rect 18612 24966 18869 24998
rect 18544 24919 18578 24935
rect 18825 24945 18869 24966
rect 18672 24929 18791 24932
rect 18672 24895 18693 24929
rect 18727 24925 18791 24929
rect 18727 24895 18729 24925
rect 18672 24891 18729 24895
rect 18763 24891 18791 24925
rect 18859 24911 18869 24945
rect 18909 24989 18943 25034
rect 18909 24933 18943 24955
rect 18999 25067 19033 25125
rect 18999 24975 19033 25033
rect 18825 24895 18869 24911
rect 18672 24884 18791 24891
rect 18909 24878 18943 24894
rect 18455 24793 18489 24849
rect 18523 24843 18539 24877
rect 18573 24850 18634 24877
rect 18855 24850 18909 24861
rect 18573 24844 18909 24850
rect 18573 24843 18943 24844
rect 18523 24827 18943 24843
rect 18999 24883 19033 24941
rect 18608 24816 18881 24827
rect 18999 24793 19033 24849
rect 18455 24791 18531 24793
rect 18489 24759 18531 24791
rect 18565 24759 18581 24793
rect 18489 24757 18581 24759
rect 18455 24740 18581 24757
rect 18683 24748 18699 24782
rect 18733 24772 18873 24782
rect 18733 24748 18822 24772
rect 18455 24699 18489 24740
rect 18683 24736 18822 24748
rect 18858 24736 18873 24772
rect 18907 24759 18923 24793
rect 18957 24791 19033 24793
rect 18957 24759 18999 24791
rect 18907 24757 18999 24759
rect 18907 24743 19033 24757
rect 18683 24726 18873 24736
rect 18999 24699 19033 24743
rect 18455 24621 18489 24665
rect 18523 24691 18947 24692
rect 18523 24689 18693 24691
rect 18523 24655 18539 24689
rect 18573 24655 18607 24689
rect 18641 24657 18693 24689
rect 18727 24689 18947 24691
rect 18727 24657 18897 24689
rect 18641 24655 18897 24657
rect 18931 24655 18947 24689
rect 18999 24621 19033 24665
rect 18455 24607 18589 24621
rect 18489 24605 18589 24607
rect 18489 24573 18555 24605
rect 18455 24571 18555 24573
rect 18455 24555 18589 24571
rect 18623 24612 18752 24620
rect 18623 24578 18625 24612
rect 18659 24586 18752 24612
rect 18786 24586 18889 24620
rect 18659 24578 18889 24586
rect 18623 24574 18889 24578
rect 18455 24515 18489 24555
rect 18623 24521 18657 24574
rect 18523 24487 18539 24521
rect 18573 24487 18607 24521
rect 18641 24487 18657 24521
rect 18691 24522 18821 24540
rect 18455 24452 18489 24481
rect 18691 24486 18754 24522
rect 18790 24518 18821 24522
rect 18691 24484 18767 24486
rect 18801 24484 18821 24518
rect 18855 24521 18889 24574
rect 18923 24607 19033 24621
rect 18923 24605 18999 24607
rect 18957 24573 18999 24605
rect 18957 24571 19033 24573
rect 18923 24555 19033 24571
rect 18855 24487 18897 24521
rect 18931 24487 18947 24521
rect 18999 24515 19033 24555
rect 18691 24470 18821 24484
rect 18999 24452 19033 24481
rect 7546 23371 7575 23405
rect 7609 23371 7667 23405
rect 7701 23371 7759 23405
rect 7793 23371 7851 23405
rect 7885 23371 7943 23405
rect 7977 23371 8035 23405
rect 8069 23371 8127 23405
rect 8161 23371 8219 23405
rect 8253 23371 8311 23405
rect 8345 23371 8403 23405
rect 8437 23371 8495 23405
rect 8529 23371 8587 23405
rect 8621 23371 8679 23405
rect 8713 23371 8771 23405
rect 8805 23371 8863 23405
rect 8897 23371 8955 23405
rect 8989 23371 9047 23405
rect 9081 23371 9139 23405
rect 9173 23371 9231 23405
rect 9265 23371 9323 23405
rect 9357 23371 9386 23405
rect 9760 23379 9789 23413
rect 9823 23379 9881 23413
rect 9915 23379 9973 23413
rect 10007 23379 10065 23413
rect 10099 23379 10157 23413
rect 10191 23379 10249 23413
rect 10283 23379 10341 23413
rect 10375 23379 10433 23413
rect 10467 23379 10525 23413
rect 10559 23379 10617 23413
rect 10651 23379 10709 23413
rect 10743 23379 10801 23413
rect 10835 23379 10893 23413
rect 10927 23379 10985 23413
rect 11019 23379 11077 23413
rect 11111 23379 11169 23413
rect 11203 23379 11261 23413
rect 11295 23379 11353 23413
rect 11387 23379 11445 23413
rect 11479 23379 11537 23413
rect 11571 23379 11600 23413
rect 7581 23321 7615 23337
rect 7581 23253 7615 23287
rect 7649 23305 7715 23371
rect 7649 23271 7665 23305
rect 7699 23271 7715 23305
rect 7749 23321 7786 23337
rect 7783 23287 7786 23321
rect 7749 23253 7786 23287
rect 7834 23329 7887 23371
rect 7834 23295 7853 23329
rect 7834 23279 7887 23295
rect 7921 23321 7971 23337
rect 7921 23287 7937 23321
rect 8268 23329 8302 23371
rect 7615 23235 7714 23237
rect 7615 23219 7672 23235
rect 7581 23203 7672 23219
rect 7668 23201 7672 23203
rect 7706 23201 7714 23235
rect 7564 23106 7634 23169
rect 7564 23093 7580 23106
rect 7564 23059 7578 23093
rect 7616 23070 7634 23106
rect 7612 23059 7634 23070
rect 7564 23039 7634 23059
rect 7668 23108 7714 23201
rect 7668 23074 7680 23108
rect 7668 23005 7714 23074
rect 7581 22971 7714 23005
rect 7783 23219 7786 23253
rect 7921 23252 7971 23287
rect 8013 23282 8029 23316
rect 8063 23282 8234 23316
rect 7749 23167 7786 23219
rect 7910 23226 7971 23252
rect 8060 23235 8166 23248
rect 7749 23133 7751 23167
rect 7785 23133 7786 23167
rect 7581 22963 7615 22971
rect 7749 22963 7786 23133
rect 7820 23161 7876 23177
rect 7820 23127 7842 23161
rect 7820 23038 7876 23127
rect 7820 23002 7830 23038
rect 7866 23002 7876 23038
rect 7820 22987 7876 23002
rect 7910 23005 7944 23226
rect 8060 23201 8092 23235
rect 8126 23209 8166 23235
rect 7978 23167 8026 23188
rect 7978 23133 7989 23167
rect 8023 23133 8026 23167
rect 7978 23131 8026 23133
rect 7978 23097 7985 23131
rect 8019 23097 8026 23131
rect 7978 23069 8026 23097
rect 8060 23035 8094 23201
rect 8128 23175 8166 23209
rect 8200 23159 8234 23282
rect 8268 23261 8302 23295
rect 8268 23211 8302 23227
rect 8336 23321 8386 23337
rect 8336 23287 8352 23321
rect 8644 23321 8707 23371
rect 8336 23271 8386 23287
rect 8431 23277 8447 23311
rect 8481 23277 8608 23311
rect 8200 23143 8302 23159
rect 8200 23141 8268 23143
rect 7910 22979 7955 23005
rect 7989 23001 8005 23035
rect 8039 23001 8094 23035
rect 7989 22991 8094 23001
rect 8128 23109 8268 23141
rect 8128 23107 8302 23109
rect 7581 22913 7615 22929
rect 7649 22903 7665 22937
rect 7699 22903 7715 22937
rect 7783 22929 7786 22963
rect 7749 22913 7786 22929
rect 7837 22937 7887 22953
rect 7649 22861 7715 22903
rect 7837 22903 7853 22937
rect 7921 22951 7955 22979
rect 8128 22951 8162 23107
rect 8268 23093 8302 23107
rect 8204 23057 8244 23063
rect 8336 23057 8370 23271
rect 8404 23235 8442 23237
rect 8404 23201 8406 23235
rect 8440 23201 8442 23235
rect 8404 23143 8442 23201
rect 8438 23109 8442 23143
rect 8404 23093 8442 23109
rect 8476 23209 8540 23243
rect 8476 23175 8506 23209
rect 8476 23167 8540 23175
rect 8476 23133 8493 23167
rect 8527 23133 8540 23167
rect 8204 23047 8370 23057
rect 8476 23051 8540 23133
rect 8238 23013 8370 23047
rect 8204 22997 8370 23013
rect 7921 22917 7938 22951
rect 7972 22917 7988 22951
rect 8027 22917 8049 22951
rect 8083 22917 8162 22951
rect 8226 22945 8300 22961
rect 7837 22861 7887 22903
rect 8226 22911 8248 22945
rect 8282 22911 8300 22945
rect 8336 22951 8370 22997
rect 8447 23035 8540 23051
rect 8481 23001 8540 23035
rect 8447 22985 8540 23001
rect 8574 23109 8608 23277
rect 8644 23287 8646 23321
rect 8680 23287 8707 23321
rect 8644 23271 8707 23287
rect 8754 23329 8822 23337
rect 8754 23295 8770 23329
rect 8804 23295 8822 23329
rect 8754 23258 8822 23295
rect 8754 23225 8770 23258
rect 8642 23224 8770 23225
rect 8804 23224 8822 23258
rect 8642 23209 8822 23224
rect 8676 23187 8822 23209
rect 8676 23175 8770 23187
rect 8642 23153 8770 23175
rect 8804 23153 8822 23187
rect 8856 23299 8890 23371
rect 9028 23329 9094 23333
rect 8856 23219 8890 23265
rect 8856 23169 8890 23185
rect 8924 23323 8990 23328
rect 8924 23289 8940 23323
rect 8974 23289 8990 23323
rect 8924 23255 8990 23289
rect 8924 23221 8940 23255
rect 8974 23221 8990 23255
rect 8924 23187 8990 23221
rect 9028 23295 9044 23329
rect 9078 23295 9094 23329
rect 9028 23261 9094 23295
rect 9028 23227 9044 23261
rect 9078 23227 9094 23261
rect 9028 23187 9094 23227
rect 8642 23150 8822 23153
rect 8784 23109 8822 23150
rect 8924 23153 8940 23187
rect 8974 23159 8990 23187
rect 8974 23153 9006 23159
rect 8924 23143 9006 23153
rect 8959 23133 9006 23143
rect 8574 23093 8750 23109
rect 8574 23059 8716 23093
rect 8574 23043 8750 23059
rect 8784 23093 8934 23109
rect 8784 23059 8900 23093
rect 8784 23043 8934 23059
rect 8574 22951 8608 23043
rect 8784 23009 8824 23043
rect 8968 23017 9006 23133
rect 8957 23009 9006 23017
rect 8758 23006 8824 23009
rect 8758 22972 8774 23006
rect 8808 22972 8824 23006
rect 8926 23008 9006 23009
rect 8336 22917 8367 22951
rect 8401 22917 8417 22951
rect 8451 22917 8470 22951
rect 8504 22917 8608 22951
rect 8663 22951 8705 22967
rect 8663 22917 8668 22951
rect 8702 22917 8705 22951
rect 8226 22861 8300 22911
rect 8663 22861 8705 22917
rect 8758 22938 8824 22972
rect 8758 22904 8774 22938
rect 8808 22904 8824 22938
rect 8858 22967 8892 22983
rect 8858 22861 8892 22933
rect 8926 22974 8942 23008
rect 8976 22992 9006 23008
rect 9040 23109 9094 23187
rect 9132 23329 9175 23371
rect 9132 23295 9141 23329
rect 9132 23261 9175 23295
rect 9132 23227 9141 23261
rect 9132 23193 9175 23227
rect 9132 23159 9141 23193
rect 9132 23143 9175 23159
rect 9209 23329 9276 23337
rect 9209 23295 9225 23329
rect 9259 23295 9276 23329
rect 9209 23258 9276 23295
rect 9209 23224 9225 23258
rect 9259 23224 9276 23258
rect 9209 23190 9276 23224
rect 9209 23187 9230 23190
rect 9209 23153 9225 23187
rect 9266 23156 9276 23190
rect 9259 23153 9276 23156
rect 9209 23140 9276 23153
rect 9040 23093 9195 23109
rect 9040 23059 9161 23093
rect 9040 23043 9195 23059
rect 8976 22974 8992 22992
rect 8926 22940 8992 22974
rect 9040 22967 9080 23043
rect 9229 23026 9276 23140
rect 9311 23300 9369 23371
rect 9311 23266 9323 23300
rect 9357 23266 9369 23300
rect 9311 23207 9369 23266
rect 9795 23329 9829 23345
rect 9795 23261 9829 23295
rect 9863 23313 9929 23379
rect 9863 23279 9879 23313
rect 9913 23279 9929 23313
rect 9963 23329 10000 23345
rect 9997 23295 10000 23329
rect 9963 23261 10000 23295
rect 10048 23337 10101 23379
rect 10048 23303 10067 23337
rect 10048 23287 10101 23303
rect 10135 23329 10185 23345
rect 10135 23295 10151 23329
rect 10482 23337 10516 23379
rect 9829 23243 9928 23245
rect 9829 23227 9886 23243
rect 9795 23211 9886 23227
rect 9311 23173 9323 23207
rect 9357 23173 9369 23207
rect 9882 23209 9886 23211
rect 9920 23209 9928 23243
rect 9311 23138 9369 23173
rect 9778 23114 9848 23177
rect 9778 23101 9794 23114
rect 9778 23067 9792 23101
rect 9830 23078 9848 23114
rect 9826 23067 9848 23078
rect 9778 23047 9848 23067
rect 9882 23116 9928 23209
rect 9882 23082 9894 23116
rect 8926 22906 8942 22940
rect 8976 22906 8992 22940
rect 9030 22963 9080 22967
rect 9030 22929 9046 22963
rect 9225 22975 9276 23026
rect 9882 23013 9928 23082
rect 9030 22913 9080 22929
rect 9127 22937 9191 22953
rect 8926 22905 8992 22906
rect 9127 22903 9141 22937
rect 9175 22903 9191 22937
rect 9127 22861 9191 22903
rect 9259 22941 9276 22975
rect 9225 22895 9276 22941
rect 9311 22989 9369 23006
rect 9311 22955 9323 22989
rect 9357 22955 9369 22989
rect 9311 22861 9369 22955
rect 9795 22979 9928 23013
rect 9997 23227 10000 23261
rect 10135 23260 10185 23295
rect 10227 23290 10243 23324
rect 10277 23290 10448 23324
rect 9963 23175 10000 23227
rect 10124 23234 10185 23260
rect 10274 23243 10380 23256
rect 9963 23141 9965 23175
rect 9999 23141 10000 23175
rect 9795 22971 9829 22979
rect 9963 22971 10000 23141
rect 10034 23169 10090 23185
rect 10034 23135 10056 23169
rect 10034 23046 10090 23135
rect 10034 23010 10044 23046
rect 10080 23010 10090 23046
rect 10034 22995 10090 23010
rect 10124 23013 10158 23234
rect 10274 23209 10306 23243
rect 10340 23217 10380 23243
rect 10192 23175 10240 23196
rect 10192 23141 10203 23175
rect 10237 23141 10240 23175
rect 10192 23139 10240 23141
rect 10192 23105 10199 23139
rect 10233 23105 10240 23139
rect 10192 23077 10240 23105
rect 10274 23043 10308 23209
rect 10342 23183 10380 23217
rect 10414 23167 10448 23290
rect 10482 23269 10516 23303
rect 10482 23219 10516 23235
rect 10550 23329 10600 23345
rect 10550 23295 10566 23329
rect 10858 23329 10921 23379
rect 10550 23279 10600 23295
rect 10645 23285 10661 23319
rect 10695 23285 10822 23319
rect 10414 23151 10516 23167
rect 10414 23149 10482 23151
rect 10124 22987 10169 23013
rect 10203 23009 10219 23043
rect 10253 23009 10308 23043
rect 10203 22999 10308 23009
rect 10342 23117 10482 23149
rect 10342 23115 10516 23117
rect 9795 22921 9829 22937
rect 9863 22911 9879 22945
rect 9913 22911 9929 22945
rect 9997 22937 10000 22971
rect 9963 22921 10000 22937
rect 10051 22945 10101 22961
rect 9863 22869 9929 22911
rect 10051 22911 10067 22945
rect 10135 22959 10169 22987
rect 10342 22959 10376 23115
rect 10482 23101 10516 23115
rect 10418 23065 10458 23071
rect 10550 23065 10584 23279
rect 10618 23243 10656 23245
rect 10618 23209 10620 23243
rect 10654 23209 10656 23243
rect 10618 23151 10656 23209
rect 10652 23117 10656 23151
rect 10618 23101 10656 23117
rect 10690 23217 10754 23251
rect 10690 23183 10720 23217
rect 10690 23175 10754 23183
rect 10690 23141 10707 23175
rect 10741 23141 10754 23175
rect 10418 23055 10584 23065
rect 10690 23059 10754 23141
rect 10452 23021 10584 23055
rect 10418 23005 10584 23021
rect 10135 22925 10152 22959
rect 10186 22925 10202 22959
rect 10241 22925 10263 22959
rect 10297 22925 10376 22959
rect 10440 22953 10514 22969
rect 10051 22869 10101 22911
rect 10440 22919 10462 22953
rect 10496 22919 10514 22953
rect 10550 22959 10584 23005
rect 10661 23043 10754 23059
rect 10695 23009 10754 23043
rect 10661 22993 10754 23009
rect 10788 23117 10822 23285
rect 10858 23295 10860 23329
rect 10894 23295 10921 23329
rect 10858 23279 10921 23295
rect 10968 23337 11036 23345
rect 10968 23303 10984 23337
rect 11018 23303 11036 23337
rect 10968 23266 11036 23303
rect 10968 23233 10984 23266
rect 10856 23232 10984 23233
rect 11018 23232 11036 23266
rect 10856 23217 11036 23232
rect 10890 23195 11036 23217
rect 10890 23183 10984 23195
rect 10856 23161 10984 23183
rect 11018 23161 11036 23195
rect 11070 23307 11104 23379
rect 11242 23337 11308 23341
rect 11070 23227 11104 23273
rect 11070 23177 11104 23193
rect 11138 23331 11204 23336
rect 11138 23297 11154 23331
rect 11188 23297 11204 23331
rect 11138 23263 11204 23297
rect 11138 23229 11154 23263
rect 11188 23229 11204 23263
rect 11138 23195 11204 23229
rect 11242 23303 11258 23337
rect 11292 23303 11308 23337
rect 11242 23269 11308 23303
rect 11242 23235 11258 23269
rect 11292 23235 11308 23269
rect 11242 23195 11308 23235
rect 10856 23158 11036 23161
rect 10998 23117 11036 23158
rect 11138 23161 11154 23195
rect 11188 23167 11204 23195
rect 11188 23161 11220 23167
rect 11138 23151 11220 23161
rect 11173 23141 11220 23151
rect 10788 23101 10964 23117
rect 10788 23067 10930 23101
rect 10788 23051 10964 23067
rect 10998 23101 11148 23117
rect 10998 23067 11114 23101
rect 10998 23051 11148 23067
rect 10788 22959 10822 23051
rect 10998 23017 11038 23051
rect 11182 23025 11220 23141
rect 11171 23017 11220 23025
rect 10972 23014 11038 23017
rect 10972 22980 10988 23014
rect 11022 22980 11038 23014
rect 11140 23016 11220 23017
rect 10550 22925 10581 22959
rect 10615 22925 10631 22959
rect 10665 22925 10684 22959
rect 10718 22925 10822 22959
rect 10877 22959 10919 22975
rect 10877 22925 10882 22959
rect 10916 22925 10919 22959
rect 10440 22869 10514 22919
rect 10877 22869 10919 22925
rect 10972 22946 11038 22980
rect 10972 22912 10988 22946
rect 11022 22912 11038 22946
rect 11072 22975 11106 22991
rect 11072 22869 11106 22941
rect 11140 22982 11156 23016
rect 11190 23000 11220 23016
rect 11254 23117 11308 23195
rect 11346 23337 11389 23379
rect 11346 23303 11355 23337
rect 11346 23269 11389 23303
rect 11346 23235 11355 23269
rect 11346 23201 11389 23235
rect 11346 23167 11355 23201
rect 11346 23151 11389 23167
rect 11423 23337 11490 23345
rect 11423 23303 11439 23337
rect 11473 23303 11490 23337
rect 11423 23266 11490 23303
rect 11423 23232 11439 23266
rect 11473 23232 11490 23266
rect 11423 23198 11490 23232
rect 11423 23195 11444 23198
rect 11423 23161 11439 23195
rect 11480 23164 11490 23198
rect 11473 23161 11490 23164
rect 11423 23148 11490 23161
rect 11254 23101 11409 23117
rect 11254 23067 11375 23101
rect 11254 23051 11409 23067
rect 11190 22982 11206 23000
rect 11140 22948 11206 22982
rect 11254 22975 11294 23051
rect 11443 23034 11490 23148
rect 11525 23308 11583 23379
rect 11960 23361 11989 23395
rect 12023 23361 12081 23395
rect 12115 23361 12173 23395
rect 12207 23361 12265 23395
rect 12299 23361 12357 23395
rect 12391 23361 12449 23395
rect 12483 23361 12541 23395
rect 12575 23361 12633 23395
rect 12667 23361 12725 23395
rect 12759 23361 12817 23395
rect 12851 23361 12909 23395
rect 12943 23361 13001 23395
rect 13035 23361 13093 23395
rect 13127 23361 13185 23395
rect 13219 23361 13277 23395
rect 13311 23361 13369 23395
rect 13403 23361 13461 23395
rect 13495 23361 13553 23395
rect 13587 23361 13645 23395
rect 13679 23361 13737 23395
rect 13771 23361 13800 23395
rect 14174 23369 14203 23403
rect 14237 23369 14295 23403
rect 14329 23369 14387 23403
rect 14421 23369 14479 23403
rect 14513 23369 14571 23403
rect 14605 23369 14663 23403
rect 14697 23369 14755 23403
rect 14789 23369 14847 23403
rect 14881 23369 14939 23403
rect 14973 23369 15031 23403
rect 15065 23369 15123 23403
rect 15157 23369 15215 23403
rect 15249 23369 15307 23403
rect 15341 23369 15399 23403
rect 15433 23369 15491 23403
rect 15525 23369 15583 23403
rect 15617 23369 15675 23403
rect 15709 23369 15767 23403
rect 15801 23369 15859 23403
rect 15893 23369 15951 23403
rect 15985 23369 16014 23403
rect 16480 23377 16509 23411
rect 16543 23377 16601 23411
rect 16635 23377 16693 23411
rect 16727 23377 16785 23411
rect 16819 23377 16877 23411
rect 16911 23377 16969 23411
rect 17003 23377 17061 23411
rect 17095 23377 17153 23411
rect 17187 23377 17245 23411
rect 17279 23377 17337 23411
rect 17371 23377 17429 23411
rect 17463 23377 17521 23411
rect 17555 23377 17613 23411
rect 17647 23377 17705 23411
rect 17739 23377 17797 23411
rect 17831 23377 17889 23411
rect 17923 23377 17981 23411
rect 18015 23377 18073 23411
rect 18107 23377 18165 23411
rect 18199 23377 18257 23411
rect 18291 23377 18320 23411
rect 11525 23274 11537 23308
rect 11571 23274 11583 23308
rect 11525 23215 11583 23274
rect 11525 23181 11537 23215
rect 11571 23181 11583 23215
rect 11995 23311 12029 23327
rect 11995 23243 12029 23277
rect 12063 23295 12129 23361
rect 12063 23261 12079 23295
rect 12113 23261 12129 23295
rect 12163 23311 12200 23327
rect 12197 23277 12200 23311
rect 12163 23243 12200 23277
rect 12248 23319 12301 23361
rect 12248 23285 12267 23319
rect 12248 23269 12301 23285
rect 12335 23311 12385 23327
rect 12335 23277 12351 23311
rect 12682 23319 12716 23361
rect 12029 23225 12128 23227
rect 12029 23209 12086 23225
rect 11995 23193 12086 23209
rect 11525 23146 11583 23181
rect 12082 23191 12086 23193
rect 12120 23191 12128 23225
rect 11140 22914 11156 22948
rect 11190 22914 11206 22948
rect 11244 22971 11294 22975
rect 11244 22937 11260 22971
rect 11439 22983 11490 23034
rect 11978 23096 12048 23159
rect 11978 23083 11994 23096
rect 11978 23049 11992 23083
rect 12030 23060 12048 23096
rect 12026 23049 12048 23060
rect 11978 23029 12048 23049
rect 12082 23098 12128 23191
rect 12082 23064 12094 23098
rect 11244 22921 11294 22937
rect 11341 22945 11405 22961
rect 11140 22913 11206 22914
rect 11341 22911 11355 22945
rect 11389 22911 11405 22945
rect 11341 22869 11405 22911
rect 11473 22949 11490 22983
rect 11439 22903 11490 22949
rect 11525 22997 11583 23014
rect 11525 22963 11537 22997
rect 11571 22963 11583 22997
rect 12082 22995 12128 23064
rect 11525 22869 11583 22963
rect 11995 22961 12128 22995
rect 12197 23209 12200 23243
rect 12335 23242 12385 23277
rect 12427 23272 12443 23306
rect 12477 23272 12648 23306
rect 12163 23157 12200 23209
rect 12324 23216 12385 23242
rect 12474 23225 12580 23238
rect 12163 23123 12165 23157
rect 12199 23123 12200 23157
rect 11995 22953 12029 22961
rect 12163 22953 12200 23123
rect 12234 23151 12290 23167
rect 12234 23117 12256 23151
rect 12234 23028 12290 23117
rect 12234 22992 12244 23028
rect 12280 22992 12290 23028
rect 12234 22977 12290 22992
rect 12324 22995 12358 23216
rect 12474 23191 12506 23225
rect 12540 23199 12580 23225
rect 12392 23157 12440 23178
rect 12392 23123 12403 23157
rect 12437 23123 12440 23157
rect 12392 23121 12440 23123
rect 12392 23087 12399 23121
rect 12433 23087 12440 23121
rect 12392 23059 12440 23087
rect 12474 23025 12508 23191
rect 12542 23165 12580 23199
rect 12614 23149 12648 23272
rect 12682 23251 12716 23285
rect 12682 23201 12716 23217
rect 12750 23311 12800 23327
rect 12750 23277 12766 23311
rect 13058 23311 13121 23361
rect 12750 23261 12800 23277
rect 12845 23267 12861 23301
rect 12895 23267 13022 23301
rect 12614 23133 12716 23149
rect 12614 23131 12682 23133
rect 12324 22969 12369 22995
rect 12403 22991 12419 23025
rect 12453 22991 12508 23025
rect 12403 22981 12508 22991
rect 12542 23099 12682 23131
rect 12542 23097 12716 23099
rect 11995 22903 12029 22919
rect 12063 22893 12079 22927
rect 12113 22893 12129 22927
rect 12197 22919 12200 22953
rect 12163 22903 12200 22919
rect 12251 22927 12301 22943
rect 7546 22827 7575 22861
rect 7609 22827 7667 22861
rect 7701 22827 7759 22861
rect 7793 22827 7851 22861
rect 7885 22827 7943 22861
rect 7977 22827 8035 22861
rect 8069 22827 8127 22861
rect 8161 22827 8219 22861
rect 8253 22827 8311 22861
rect 8345 22827 8403 22861
rect 8437 22827 8495 22861
rect 8529 22827 8587 22861
rect 8621 22827 8679 22861
rect 8713 22827 8771 22861
rect 8805 22827 8863 22861
rect 8897 22827 8955 22861
rect 8989 22827 9047 22861
rect 9081 22827 9139 22861
rect 9173 22827 9231 22861
rect 9265 22827 9323 22861
rect 9357 22827 9386 22861
rect 9760 22835 9789 22869
rect 9823 22835 9881 22869
rect 9915 22835 9973 22869
rect 10007 22835 10065 22869
rect 10099 22835 10157 22869
rect 10191 22835 10249 22869
rect 10283 22835 10341 22869
rect 10375 22835 10433 22869
rect 10467 22835 10525 22869
rect 10559 22835 10617 22869
rect 10651 22835 10709 22869
rect 10743 22835 10801 22869
rect 10835 22835 10893 22869
rect 10927 22835 10985 22869
rect 11019 22835 11077 22869
rect 11111 22835 11169 22869
rect 11203 22835 11261 22869
rect 11295 22835 11353 22869
rect 11387 22835 11445 22869
rect 11479 22835 11537 22869
rect 11571 22835 11600 22869
rect 12063 22851 12129 22893
rect 12251 22893 12267 22927
rect 12335 22941 12369 22969
rect 12542 22941 12576 23097
rect 12682 23083 12716 23097
rect 12618 23047 12658 23053
rect 12750 23047 12784 23261
rect 12818 23225 12856 23227
rect 12818 23191 12820 23225
rect 12854 23191 12856 23225
rect 12818 23133 12856 23191
rect 12852 23099 12856 23133
rect 12818 23083 12856 23099
rect 12890 23199 12954 23233
rect 12890 23165 12920 23199
rect 12890 23157 12954 23165
rect 12890 23123 12907 23157
rect 12941 23123 12954 23157
rect 12618 23037 12784 23047
rect 12890 23041 12954 23123
rect 12652 23003 12784 23037
rect 12618 22987 12784 23003
rect 12335 22907 12352 22941
rect 12386 22907 12402 22941
rect 12441 22907 12463 22941
rect 12497 22907 12576 22941
rect 12640 22935 12714 22951
rect 12251 22851 12301 22893
rect 12640 22901 12662 22935
rect 12696 22901 12714 22935
rect 12750 22941 12784 22987
rect 12861 23025 12954 23041
rect 12895 22991 12954 23025
rect 12861 22975 12954 22991
rect 12988 23099 13022 23267
rect 13058 23277 13060 23311
rect 13094 23277 13121 23311
rect 13058 23261 13121 23277
rect 13168 23319 13236 23327
rect 13168 23285 13184 23319
rect 13218 23285 13236 23319
rect 13168 23248 13236 23285
rect 13168 23215 13184 23248
rect 13056 23214 13184 23215
rect 13218 23214 13236 23248
rect 13056 23199 13236 23214
rect 13090 23177 13236 23199
rect 13090 23165 13184 23177
rect 13056 23143 13184 23165
rect 13218 23143 13236 23177
rect 13270 23289 13304 23361
rect 13442 23319 13508 23323
rect 13270 23209 13304 23255
rect 13270 23159 13304 23175
rect 13338 23313 13404 23318
rect 13338 23279 13354 23313
rect 13388 23279 13404 23313
rect 13338 23245 13404 23279
rect 13338 23211 13354 23245
rect 13388 23211 13404 23245
rect 13338 23177 13404 23211
rect 13442 23285 13458 23319
rect 13492 23285 13508 23319
rect 13442 23251 13508 23285
rect 13442 23217 13458 23251
rect 13492 23217 13508 23251
rect 13442 23177 13508 23217
rect 13056 23140 13236 23143
rect 13198 23099 13236 23140
rect 13338 23143 13354 23177
rect 13388 23149 13404 23177
rect 13388 23143 13420 23149
rect 13338 23133 13420 23143
rect 13373 23123 13420 23133
rect 12988 23083 13164 23099
rect 12988 23049 13130 23083
rect 12988 23033 13164 23049
rect 13198 23083 13348 23099
rect 13198 23049 13314 23083
rect 13198 23033 13348 23049
rect 12988 22941 13022 23033
rect 13198 22999 13238 23033
rect 13382 23007 13420 23123
rect 13371 22999 13420 23007
rect 13172 22996 13238 22999
rect 13172 22962 13188 22996
rect 13222 22962 13238 22996
rect 13340 22998 13420 22999
rect 12750 22907 12781 22941
rect 12815 22907 12831 22941
rect 12865 22907 12884 22941
rect 12918 22907 13022 22941
rect 13077 22941 13119 22957
rect 13077 22907 13082 22941
rect 13116 22907 13119 22941
rect 12640 22851 12714 22901
rect 13077 22851 13119 22907
rect 13172 22928 13238 22962
rect 13172 22894 13188 22928
rect 13222 22894 13238 22928
rect 13272 22957 13306 22973
rect 13272 22851 13306 22923
rect 13340 22964 13356 22998
rect 13390 22982 13420 22998
rect 13454 23099 13508 23177
rect 13546 23319 13589 23361
rect 13546 23285 13555 23319
rect 13546 23251 13589 23285
rect 13546 23217 13555 23251
rect 13546 23183 13589 23217
rect 13546 23149 13555 23183
rect 13546 23133 13589 23149
rect 13623 23319 13690 23327
rect 13623 23285 13639 23319
rect 13673 23285 13690 23319
rect 13623 23248 13690 23285
rect 13623 23214 13639 23248
rect 13673 23214 13690 23248
rect 13623 23180 13690 23214
rect 13623 23177 13644 23180
rect 13623 23143 13639 23177
rect 13680 23146 13690 23180
rect 13673 23143 13690 23146
rect 13623 23130 13690 23143
rect 13454 23083 13609 23099
rect 13454 23049 13575 23083
rect 13454 23033 13609 23049
rect 13390 22964 13406 22982
rect 13340 22930 13406 22964
rect 13454 22957 13494 23033
rect 13643 23016 13690 23130
rect 13725 23290 13783 23361
rect 13725 23256 13737 23290
rect 13771 23256 13783 23290
rect 13725 23197 13783 23256
rect 14209 23319 14243 23335
rect 14209 23251 14243 23285
rect 14277 23303 14343 23369
rect 14277 23269 14293 23303
rect 14327 23269 14343 23303
rect 14377 23319 14414 23335
rect 14411 23285 14414 23319
rect 14377 23251 14414 23285
rect 14462 23327 14515 23369
rect 14462 23293 14481 23327
rect 14462 23277 14515 23293
rect 14549 23319 14599 23335
rect 14549 23285 14565 23319
rect 14896 23327 14930 23369
rect 14243 23233 14342 23235
rect 14243 23217 14300 23233
rect 14209 23201 14300 23217
rect 13725 23163 13737 23197
rect 13771 23163 13783 23197
rect 14296 23199 14300 23201
rect 14334 23199 14342 23233
rect 13725 23128 13783 23163
rect 14192 23104 14262 23167
rect 14192 23091 14208 23104
rect 14192 23057 14206 23091
rect 14244 23068 14262 23104
rect 14240 23057 14262 23068
rect 14192 23037 14262 23057
rect 14296 23106 14342 23199
rect 14296 23072 14308 23106
rect 13340 22896 13356 22930
rect 13390 22896 13406 22930
rect 13444 22953 13494 22957
rect 13444 22919 13460 22953
rect 13639 22965 13690 23016
rect 14296 23003 14342 23072
rect 13444 22903 13494 22919
rect 13541 22927 13605 22943
rect 13340 22895 13406 22896
rect 13541 22893 13555 22927
rect 13589 22893 13605 22927
rect 13541 22851 13605 22893
rect 13673 22931 13690 22965
rect 13639 22885 13690 22931
rect 13725 22979 13783 22996
rect 13725 22945 13737 22979
rect 13771 22945 13783 22979
rect 13725 22851 13783 22945
rect 14209 22969 14342 23003
rect 14411 23217 14414 23251
rect 14549 23250 14599 23285
rect 14641 23280 14657 23314
rect 14691 23280 14862 23314
rect 14377 23165 14414 23217
rect 14538 23224 14599 23250
rect 14688 23233 14794 23246
rect 14377 23131 14379 23165
rect 14413 23131 14414 23165
rect 14209 22961 14243 22969
rect 14377 22961 14414 23131
rect 14448 23159 14504 23175
rect 14448 23125 14470 23159
rect 14448 23036 14504 23125
rect 14448 23000 14458 23036
rect 14494 23000 14504 23036
rect 14448 22985 14504 23000
rect 14538 23003 14572 23224
rect 14688 23199 14720 23233
rect 14754 23207 14794 23233
rect 14606 23165 14654 23186
rect 14606 23131 14617 23165
rect 14651 23131 14654 23165
rect 14606 23129 14654 23131
rect 14606 23095 14613 23129
rect 14647 23095 14654 23129
rect 14606 23067 14654 23095
rect 14688 23033 14722 23199
rect 14756 23173 14794 23207
rect 14828 23157 14862 23280
rect 14896 23259 14930 23293
rect 14896 23209 14930 23225
rect 14964 23319 15014 23335
rect 14964 23285 14980 23319
rect 15272 23319 15335 23369
rect 14964 23269 15014 23285
rect 15059 23275 15075 23309
rect 15109 23275 15236 23309
rect 14828 23141 14930 23157
rect 14828 23139 14896 23141
rect 14538 22977 14583 23003
rect 14617 22999 14633 23033
rect 14667 22999 14722 23033
rect 14617 22989 14722 22999
rect 14756 23107 14896 23139
rect 14756 23105 14930 23107
rect 14209 22911 14243 22927
rect 14277 22901 14293 22935
rect 14327 22901 14343 22935
rect 14411 22927 14414 22961
rect 14377 22911 14414 22927
rect 14465 22935 14515 22951
rect 14277 22859 14343 22901
rect 14465 22901 14481 22935
rect 14549 22949 14583 22977
rect 14756 22949 14790 23105
rect 14896 23091 14930 23105
rect 14832 23055 14872 23061
rect 14964 23055 14998 23269
rect 15032 23233 15070 23235
rect 15032 23199 15034 23233
rect 15068 23199 15070 23233
rect 15032 23141 15070 23199
rect 15066 23107 15070 23141
rect 15032 23091 15070 23107
rect 15104 23207 15168 23241
rect 15104 23173 15134 23207
rect 15104 23165 15168 23173
rect 15104 23131 15121 23165
rect 15155 23131 15168 23165
rect 14832 23045 14998 23055
rect 15104 23049 15168 23131
rect 14866 23011 14998 23045
rect 14832 22995 14998 23011
rect 14549 22915 14566 22949
rect 14600 22915 14616 22949
rect 14655 22915 14677 22949
rect 14711 22915 14790 22949
rect 14854 22943 14928 22959
rect 14465 22859 14515 22901
rect 14854 22909 14876 22943
rect 14910 22909 14928 22943
rect 14964 22949 14998 22995
rect 15075 23033 15168 23049
rect 15109 22999 15168 23033
rect 15075 22983 15168 22999
rect 15202 23107 15236 23275
rect 15272 23285 15274 23319
rect 15308 23285 15335 23319
rect 15272 23269 15335 23285
rect 15382 23327 15450 23335
rect 15382 23293 15398 23327
rect 15432 23293 15450 23327
rect 15382 23256 15450 23293
rect 15382 23223 15398 23256
rect 15270 23222 15398 23223
rect 15432 23222 15450 23256
rect 15270 23207 15450 23222
rect 15304 23185 15450 23207
rect 15304 23173 15398 23185
rect 15270 23151 15398 23173
rect 15432 23151 15450 23185
rect 15484 23297 15518 23369
rect 15656 23327 15722 23331
rect 15484 23217 15518 23263
rect 15484 23167 15518 23183
rect 15552 23321 15618 23326
rect 15552 23287 15568 23321
rect 15602 23287 15618 23321
rect 15552 23253 15618 23287
rect 15552 23219 15568 23253
rect 15602 23219 15618 23253
rect 15552 23185 15618 23219
rect 15656 23293 15672 23327
rect 15706 23293 15722 23327
rect 15656 23259 15722 23293
rect 15656 23225 15672 23259
rect 15706 23225 15722 23259
rect 15656 23185 15722 23225
rect 15270 23148 15450 23151
rect 15412 23107 15450 23148
rect 15552 23151 15568 23185
rect 15602 23157 15618 23185
rect 15602 23151 15634 23157
rect 15552 23141 15634 23151
rect 15587 23131 15634 23141
rect 15202 23091 15378 23107
rect 15202 23057 15344 23091
rect 15202 23041 15378 23057
rect 15412 23091 15562 23107
rect 15412 23057 15528 23091
rect 15412 23041 15562 23057
rect 15202 22949 15236 23041
rect 15412 23007 15452 23041
rect 15596 23015 15634 23131
rect 15585 23007 15634 23015
rect 15386 23004 15452 23007
rect 15386 22970 15402 23004
rect 15436 22970 15452 23004
rect 15554 23006 15634 23007
rect 14964 22915 14995 22949
rect 15029 22915 15045 22949
rect 15079 22915 15098 22949
rect 15132 22915 15236 22949
rect 15291 22949 15333 22965
rect 15291 22915 15296 22949
rect 15330 22915 15333 22949
rect 14854 22859 14928 22909
rect 15291 22859 15333 22915
rect 15386 22936 15452 22970
rect 15386 22902 15402 22936
rect 15436 22902 15452 22936
rect 15486 22965 15520 22981
rect 15486 22859 15520 22931
rect 15554 22972 15570 23006
rect 15604 22990 15634 23006
rect 15668 23107 15722 23185
rect 15760 23327 15803 23369
rect 15760 23293 15769 23327
rect 15760 23259 15803 23293
rect 15760 23225 15769 23259
rect 15760 23191 15803 23225
rect 15760 23157 15769 23191
rect 15760 23141 15803 23157
rect 15837 23327 15904 23335
rect 15837 23293 15853 23327
rect 15887 23293 15904 23327
rect 15837 23256 15904 23293
rect 15837 23222 15853 23256
rect 15887 23222 15904 23256
rect 15837 23188 15904 23222
rect 15837 23185 15858 23188
rect 15837 23151 15853 23185
rect 15894 23154 15904 23188
rect 15887 23151 15904 23154
rect 15837 23138 15904 23151
rect 15668 23091 15823 23107
rect 15668 23057 15789 23091
rect 15668 23041 15823 23057
rect 15604 22972 15620 22990
rect 15554 22938 15620 22972
rect 15668 22965 15708 23041
rect 15857 23024 15904 23138
rect 15939 23298 15997 23369
rect 15939 23264 15951 23298
rect 15985 23264 15997 23298
rect 15939 23205 15997 23264
rect 16515 23327 16549 23343
rect 16515 23259 16549 23293
rect 16583 23311 16649 23377
rect 16583 23277 16599 23311
rect 16633 23277 16649 23311
rect 16683 23327 16720 23343
rect 16717 23293 16720 23327
rect 16683 23259 16720 23293
rect 16768 23335 16821 23377
rect 16768 23301 16787 23335
rect 16768 23285 16821 23301
rect 16855 23327 16905 23343
rect 16855 23293 16871 23327
rect 17202 23335 17236 23377
rect 16549 23241 16648 23243
rect 16549 23225 16606 23241
rect 16515 23209 16606 23225
rect 15939 23171 15951 23205
rect 15985 23171 15997 23205
rect 16602 23207 16606 23209
rect 16640 23207 16648 23241
rect 15939 23136 15997 23171
rect 16498 23112 16568 23175
rect 16498 23099 16514 23112
rect 16498 23065 16512 23099
rect 16550 23076 16568 23112
rect 16546 23065 16568 23076
rect 16498 23045 16568 23065
rect 16602 23114 16648 23207
rect 16602 23080 16614 23114
rect 15554 22904 15570 22938
rect 15604 22904 15620 22938
rect 15658 22961 15708 22965
rect 15658 22927 15674 22961
rect 15853 22973 15904 23024
rect 16602 23011 16648 23080
rect 15658 22911 15708 22927
rect 15755 22935 15819 22951
rect 15554 22903 15620 22904
rect 15755 22901 15769 22935
rect 15803 22901 15819 22935
rect 15755 22859 15819 22901
rect 15887 22939 15904 22973
rect 15853 22893 15904 22939
rect 15939 22987 15997 23004
rect 15939 22953 15951 22987
rect 15985 22953 15997 22987
rect 15939 22859 15997 22953
rect 16515 22977 16648 23011
rect 16717 23225 16720 23259
rect 16855 23258 16905 23293
rect 16947 23288 16963 23322
rect 16997 23288 17168 23322
rect 16683 23173 16720 23225
rect 16844 23232 16905 23258
rect 16994 23241 17100 23254
rect 16683 23139 16685 23173
rect 16719 23139 16720 23173
rect 16515 22969 16549 22977
rect 16683 22969 16720 23139
rect 16754 23167 16810 23183
rect 16754 23133 16776 23167
rect 16754 23044 16810 23133
rect 16754 23008 16764 23044
rect 16800 23008 16810 23044
rect 16754 22993 16810 23008
rect 16844 23011 16878 23232
rect 16994 23207 17026 23241
rect 17060 23215 17100 23241
rect 16912 23173 16960 23194
rect 16912 23139 16923 23173
rect 16957 23139 16960 23173
rect 16912 23137 16960 23139
rect 16912 23103 16919 23137
rect 16953 23103 16960 23137
rect 16912 23075 16960 23103
rect 16994 23041 17028 23207
rect 17062 23181 17100 23215
rect 17134 23165 17168 23288
rect 17202 23267 17236 23301
rect 17202 23217 17236 23233
rect 17270 23327 17320 23343
rect 17270 23293 17286 23327
rect 17578 23327 17641 23377
rect 17270 23277 17320 23293
rect 17365 23283 17381 23317
rect 17415 23283 17542 23317
rect 17134 23149 17236 23165
rect 17134 23147 17202 23149
rect 16844 22985 16889 23011
rect 16923 23007 16939 23041
rect 16973 23007 17028 23041
rect 16923 22997 17028 23007
rect 17062 23115 17202 23147
rect 17062 23113 17236 23115
rect 16515 22919 16549 22935
rect 16583 22909 16599 22943
rect 16633 22909 16649 22943
rect 16717 22935 16720 22969
rect 16683 22919 16720 22935
rect 16771 22943 16821 22959
rect 16583 22867 16649 22909
rect 16771 22909 16787 22943
rect 16855 22957 16889 22985
rect 17062 22957 17096 23113
rect 17202 23099 17236 23113
rect 17138 23063 17178 23069
rect 17270 23063 17304 23277
rect 17338 23241 17376 23243
rect 17338 23207 17340 23241
rect 17374 23207 17376 23241
rect 17338 23149 17376 23207
rect 17372 23115 17376 23149
rect 17338 23099 17376 23115
rect 17410 23215 17474 23249
rect 17410 23181 17440 23215
rect 17410 23173 17474 23181
rect 17410 23139 17427 23173
rect 17461 23139 17474 23173
rect 17138 23053 17304 23063
rect 17410 23057 17474 23139
rect 17172 23019 17304 23053
rect 17138 23003 17304 23019
rect 16855 22923 16872 22957
rect 16906 22923 16922 22957
rect 16961 22923 16983 22957
rect 17017 22923 17096 22957
rect 17160 22951 17234 22967
rect 16771 22867 16821 22909
rect 17160 22917 17182 22951
rect 17216 22917 17234 22951
rect 17270 22957 17304 23003
rect 17381 23041 17474 23057
rect 17415 23007 17474 23041
rect 17381 22991 17474 23007
rect 17508 23115 17542 23283
rect 17578 23293 17580 23327
rect 17614 23293 17641 23327
rect 17578 23277 17641 23293
rect 17688 23335 17756 23343
rect 17688 23301 17704 23335
rect 17738 23301 17756 23335
rect 17688 23264 17756 23301
rect 17688 23231 17704 23264
rect 17576 23230 17704 23231
rect 17738 23230 17756 23264
rect 17576 23215 17756 23230
rect 17610 23193 17756 23215
rect 17610 23181 17704 23193
rect 17576 23159 17704 23181
rect 17738 23159 17756 23193
rect 17790 23305 17824 23377
rect 17962 23335 18028 23339
rect 17790 23225 17824 23271
rect 17790 23175 17824 23191
rect 17858 23329 17924 23334
rect 17858 23295 17874 23329
rect 17908 23295 17924 23329
rect 17858 23261 17924 23295
rect 17858 23227 17874 23261
rect 17908 23227 17924 23261
rect 17858 23193 17924 23227
rect 17962 23301 17978 23335
rect 18012 23301 18028 23335
rect 17962 23267 18028 23301
rect 17962 23233 17978 23267
rect 18012 23233 18028 23267
rect 17962 23193 18028 23233
rect 17576 23156 17756 23159
rect 17718 23115 17756 23156
rect 17858 23159 17874 23193
rect 17908 23165 17924 23193
rect 17908 23159 17940 23165
rect 17858 23149 17940 23159
rect 17893 23139 17940 23149
rect 17508 23099 17684 23115
rect 17508 23065 17650 23099
rect 17508 23049 17684 23065
rect 17718 23099 17868 23115
rect 17718 23065 17834 23099
rect 17718 23049 17868 23065
rect 17508 22957 17542 23049
rect 17718 23015 17758 23049
rect 17902 23023 17940 23139
rect 17891 23015 17940 23023
rect 17692 23012 17758 23015
rect 17692 22978 17708 23012
rect 17742 22978 17758 23012
rect 17860 23014 17940 23015
rect 17270 22923 17301 22957
rect 17335 22923 17351 22957
rect 17385 22923 17404 22957
rect 17438 22923 17542 22957
rect 17597 22957 17639 22973
rect 17597 22923 17602 22957
rect 17636 22923 17639 22957
rect 17160 22867 17234 22917
rect 17597 22867 17639 22923
rect 17692 22944 17758 22978
rect 17692 22910 17708 22944
rect 17742 22910 17758 22944
rect 17792 22973 17826 22989
rect 17792 22867 17826 22939
rect 17860 22980 17876 23014
rect 17910 22998 17940 23014
rect 17974 23115 18028 23193
rect 18066 23335 18109 23377
rect 18066 23301 18075 23335
rect 18066 23267 18109 23301
rect 18066 23233 18075 23267
rect 18066 23199 18109 23233
rect 18066 23165 18075 23199
rect 18066 23149 18109 23165
rect 18143 23335 18210 23343
rect 18143 23301 18159 23335
rect 18193 23301 18210 23335
rect 18143 23264 18210 23301
rect 18143 23230 18159 23264
rect 18193 23230 18210 23264
rect 18143 23196 18210 23230
rect 18143 23193 18164 23196
rect 18143 23159 18159 23193
rect 18200 23162 18210 23196
rect 18193 23159 18210 23162
rect 18143 23146 18210 23159
rect 17974 23099 18129 23115
rect 17974 23065 18095 23099
rect 17974 23049 18129 23065
rect 17910 22980 17926 22998
rect 17860 22946 17926 22980
rect 17974 22973 18014 23049
rect 18163 23032 18210 23146
rect 18245 23306 18303 23377
rect 18245 23272 18257 23306
rect 18291 23272 18303 23306
rect 18245 23213 18303 23272
rect 18245 23179 18257 23213
rect 18291 23179 18303 23213
rect 18245 23144 18303 23179
rect 17860 22912 17876 22946
rect 17910 22912 17926 22946
rect 17964 22969 18014 22973
rect 17964 22935 17980 22969
rect 18159 22981 18210 23032
rect 17964 22919 18014 22935
rect 18061 22943 18125 22959
rect 17860 22911 17926 22912
rect 18061 22909 18075 22943
rect 18109 22909 18125 22943
rect 18061 22867 18125 22909
rect 18193 22947 18210 22981
rect 18159 22901 18210 22947
rect 18245 22995 18303 23012
rect 18245 22961 18257 22995
rect 18291 22961 18303 22995
rect 18245 22867 18303 22961
rect 11960 22817 11989 22851
rect 12023 22817 12081 22851
rect 12115 22817 12173 22851
rect 12207 22817 12265 22851
rect 12299 22817 12357 22851
rect 12391 22817 12449 22851
rect 12483 22817 12541 22851
rect 12575 22817 12633 22851
rect 12667 22817 12725 22851
rect 12759 22817 12817 22851
rect 12851 22817 12909 22851
rect 12943 22817 13001 22851
rect 13035 22817 13093 22851
rect 13127 22817 13185 22851
rect 13219 22817 13277 22851
rect 13311 22817 13369 22851
rect 13403 22817 13461 22851
rect 13495 22817 13553 22851
rect 13587 22817 13645 22851
rect 13679 22817 13737 22851
rect 13771 22817 13800 22851
rect 14174 22825 14203 22859
rect 14237 22825 14295 22859
rect 14329 22825 14387 22859
rect 14421 22825 14479 22859
rect 14513 22825 14571 22859
rect 14605 22825 14663 22859
rect 14697 22825 14755 22859
rect 14789 22825 14847 22859
rect 14881 22825 14939 22859
rect 14973 22825 15031 22859
rect 15065 22825 15123 22859
rect 15157 22825 15215 22859
rect 15249 22825 15307 22859
rect 15341 22825 15399 22859
rect 15433 22825 15491 22859
rect 15525 22825 15583 22859
rect 15617 22825 15675 22859
rect 15709 22825 15767 22859
rect 15801 22825 15859 22859
rect 15893 22825 15951 22859
rect 15985 22825 16014 22859
rect 16480 22833 16509 22867
rect 16543 22833 16601 22867
rect 16635 22833 16693 22867
rect 16727 22833 16785 22867
rect 16819 22833 16877 22867
rect 16911 22833 16969 22867
rect 17003 22833 17061 22867
rect 17095 22833 17153 22867
rect 17187 22833 17245 22867
rect 17279 22833 17337 22867
rect 17371 22833 17429 22867
rect 17463 22833 17521 22867
rect 17555 22833 17613 22867
rect 17647 22833 17705 22867
rect 17739 22833 17797 22867
rect 17831 22833 17889 22867
rect 17923 22833 17981 22867
rect 18015 22833 18073 22867
rect 18107 22833 18165 22867
rect 18199 22833 18257 22867
rect 18291 22833 18320 22867
rect 16267 17667 16296 17701
rect 16330 17667 16374 17701
rect 16408 17667 16466 17701
rect 16500 17667 16558 17701
rect 16592 17667 16621 17701
rect 17133 17669 17162 17703
rect 17196 17669 17248 17703
rect 17282 17669 17340 17703
rect 17374 17669 17432 17703
rect 17466 17669 17495 17703
rect 15481 17629 15510 17663
rect 15544 17629 15596 17663
rect 15630 17629 15688 17663
rect 15722 17629 15780 17663
rect 15814 17629 15843 17663
rect 15498 17535 15556 17629
rect 15498 17501 15510 17535
rect 15544 17501 15556 17535
rect 15498 17484 15556 17501
rect 15633 17583 15699 17595
rect 15633 17549 15649 17583
rect 15683 17549 15699 17583
rect 15633 17515 15699 17549
rect 15633 17481 15649 17515
rect 15683 17481 15699 17515
rect 15633 17469 15699 17481
rect 15733 17583 15779 17629
rect 15767 17549 15779 17583
rect 15733 17515 15779 17549
rect 16284 17573 16342 17667
rect 16284 17539 16296 17573
rect 16330 17539 16342 17573
rect 16284 17522 16342 17539
rect 16411 17621 16477 17633
rect 16411 17587 16427 17621
rect 16461 17587 16477 17621
rect 16411 17553 16477 17587
rect 15767 17481 15779 17515
rect 15633 17436 15679 17469
rect 15733 17465 15779 17481
rect 16411 17519 16427 17553
rect 16461 17519 16477 17553
rect 16411 17507 16477 17519
rect 16511 17621 16557 17667
rect 16545 17587 16557 17621
rect 16511 17553 16557 17587
rect 16545 17519 16557 17553
rect 17150 17575 17208 17669
rect 17150 17541 17162 17575
rect 17196 17541 17208 17575
rect 17150 17524 17208 17541
rect 17285 17623 17351 17635
rect 17285 17589 17301 17623
rect 17335 17589 17351 17623
rect 17285 17555 17351 17589
rect 16411 17468 16457 17507
rect 16511 17503 16557 17519
rect 17285 17521 17301 17555
rect 17335 17521 17351 17555
rect 17285 17509 17351 17521
rect 17385 17623 17431 17669
rect 17911 17659 17940 17693
rect 17974 17659 18016 17693
rect 18050 17659 18108 17693
rect 18142 17659 18200 17693
rect 18234 17659 18263 17693
rect 19027 17661 19056 17695
rect 19090 17661 19138 17695
rect 19172 17661 19230 17695
rect 19264 17661 19322 17695
rect 19356 17661 19385 17695
rect 19893 17663 19922 17697
rect 19956 17663 20012 17697
rect 20046 17663 20104 17697
rect 20138 17663 20196 17697
rect 20230 17663 20259 17697
rect 17419 17589 17431 17623
rect 17385 17555 17431 17589
rect 17419 17521 17431 17555
rect 17285 17476 17331 17509
rect 17385 17505 17431 17521
rect 17928 17565 17986 17659
rect 17928 17531 17940 17565
rect 17974 17531 17986 17565
rect 17928 17514 17986 17531
rect 18053 17613 18119 17625
rect 18053 17579 18069 17613
rect 18103 17579 18119 17613
rect 18053 17545 18119 17579
rect 18053 17511 18069 17545
rect 18103 17511 18119 17545
rect 15633 17402 15635 17436
rect 15669 17402 15679 17436
rect 16411 17434 16413 17468
rect 16449 17434 16457 17468
rect 15498 17317 15556 17352
rect 15498 17283 15510 17317
rect 15544 17283 15556 17317
rect 15498 17224 15556 17283
rect 15498 17190 15510 17224
rect 15544 17190 15556 17224
rect 15498 17119 15556 17190
rect 15633 17349 15679 17402
rect 15713 17428 15729 17431
rect 15713 17394 15725 17428
rect 15763 17394 15779 17431
rect 15713 17383 15779 17394
rect 16284 17355 16342 17390
rect 15633 17331 15699 17349
rect 15633 17297 15649 17331
rect 15683 17297 15699 17331
rect 15633 17263 15699 17297
rect 15633 17229 15649 17263
rect 15683 17229 15699 17263
rect 15633 17195 15699 17229
rect 15633 17161 15649 17195
rect 15683 17161 15699 17195
rect 15633 17153 15699 17161
rect 15733 17331 15775 17347
rect 15767 17297 15775 17331
rect 15733 17263 15775 17297
rect 15767 17229 15775 17263
rect 15733 17195 15775 17229
rect 15767 17161 15775 17195
rect 15733 17119 15775 17161
rect 16284 17321 16296 17355
rect 16330 17321 16342 17355
rect 16284 17262 16342 17321
rect 16284 17228 16296 17262
rect 16330 17228 16342 17262
rect 16284 17157 16342 17228
rect 16411 17387 16457 17434
rect 16491 17435 16507 17469
rect 16541 17464 16557 17469
rect 16491 17430 16517 17435
rect 16551 17430 16557 17464
rect 16491 17421 16557 17430
rect 17285 17442 17287 17476
rect 17321 17442 17331 17476
rect 18053 17499 18119 17511
rect 18153 17613 18199 17659
rect 18187 17579 18199 17613
rect 18153 17545 18199 17579
rect 18187 17511 18199 17545
rect 19044 17567 19102 17661
rect 19044 17533 19056 17567
rect 19090 17533 19102 17567
rect 19044 17516 19102 17533
rect 19175 17615 19241 17627
rect 19175 17581 19191 17615
rect 19225 17581 19241 17615
rect 19175 17547 19241 17581
rect 18053 17472 18099 17499
rect 18153 17495 18199 17511
rect 19175 17513 19191 17547
rect 19225 17513 19241 17547
rect 19175 17501 19241 17513
rect 19275 17615 19321 17661
rect 19309 17581 19321 17615
rect 19275 17547 19321 17581
rect 19309 17513 19321 17547
rect 19910 17569 19968 17663
rect 19910 17535 19922 17569
rect 19956 17535 19968 17569
rect 19910 17518 19968 17535
rect 20049 17617 20115 17629
rect 20049 17583 20065 17617
rect 20099 17583 20115 17617
rect 20049 17549 20115 17583
rect 16411 17369 16477 17387
rect 16411 17335 16427 17369
rect 16461 17335 16477 17369
rect 16411 17301 16477 17335
rect 16411 17267 16427 17301
rect 16461 17267 16477 17301
rect 16411 17233 16477 17267
rect 16411 17199 16427 17233
rect 16461 17199 16477 17233
rect 16411 17191 16477 17199
rect 16511 17369 16553 17385
rect 16545 17335 16553 17369
rect 16511 17301 16553 17335
rect 16545 17267 16553 17301
rect 16511 17233 16553 17267
rect 16545 17199 16553 17233
rect 16511 17157 16553 17199
rect 17150 17357 17208 17392
rect 17150 17323 17162 17357
rect 17196 17323 17208 17357
rect 17150 17264 17208 17323
rect 17150 17230 17162 17264
rect 17196 17230 17208 17264
rect 17150 17159 17208 17230
rect 17285 17389 17331 17442
rect 17365 17468 17381 17471
rect 17365 17434 17377 17468
rect 17415 17434 17431 17471
rect 17365 17423 17431 17434
rect 18053 17438 18059 17472
rect 18097 17438 18099 17472
rect 19175 17462 19221 17501
rect 19275 17497 19321 17513
rect 20049 17515 20065 17549
rect 20099 17515 20115 17549
rect 20049 17503 20115 17515
rect 20149 17617 20195 17663
rect 20663 17653 20692 17687
rect 20726 17653 20780 17687
rect 20814 17653 20872 17687
rect 20906 17653 20964 17687
rect 20998 17653 21027 17687
rect 20183 17583 20195 17617
rect 20149 17549 20195 17583
rect 20183 17515 20195 17549
rect 20049 17470 20095 17503
rect 20149 17499 20195 17515
rect 20680 17559 20738 17653
rect 20680 17525 20692 17559
rect 20726 17525 20738 17559
rect 20680 17508 20738 17525
rect 20817 17607 20883 17619
rect 20817 17573 20833 17607
rect 20867 17573 20883 17607
rect 20817 17539 20883 17573
rect 20817 17505 20833 17539
rect 20867 17505 20883 17539
rect 17285 17371 17351 17389
rect 17285 17337 17301 17371
rect 17335 17337 17351 17371
rect 17285 17303 17351 17337
rect 17285 17269 17301 17303
rect 17335 17269 17351 17303
rect 17285 17235 17351 17269
rect 17285 17201 17301 17235
rect 17335 17201 17351 17235
rect 17285 17193 17351 17201
rect 17385 17371 17427 17387
rect 17419 17337 17427 17371
rect 17385 17303 17427 17337
rect 17419 17269 17427 17303
rect 17385 17235 17427 17269
rect 17419 17201 17427 17235
rect 17385 17159 17427 17201
rect 17928 17347 17986 17382
rect 17928 17313 17940 17347
rect 17974 17313 17986 17347
rect 17928 17254 17986 17313
rect 17928 17220 17940 17254
rect 17974 17220 17986 17254
rect 16267 17123 16296 17157
rect 16330 17123 16374 17157
rect 16408 17123 16466 17157
rect 16500 17123 16558 17157
rect 16592 17123 16621 17157
rect 17133 17125 17162 17159
rect 17196 17125 17248 17159
rect 17282 17125 17340 17159
rect 17374 17125 17432 17159
rect 17466 17125 17495 17159
rect 17928 17149 17986 17220
rect 18053 17379 18099 17438
rect 18133 17460 18149 17461
rect 18133 17426 18147 17460
rect 18183 17426 18199 17461
rect 18133 17413 18199 17426
rect 19175 17428 19177 17462
rect 19213 17428 19221 17462
rect 18053 17361 18119 17379
rect 18053 17327 18069 17361
rect 18103 17327 18119 17361
rect 18053 17293 18119 17327
rect 18053 17259 18069 17293
rect 18103 17259 18119 17293
rect 18053 17225 18119 17259
rect 18053 17191 18069 17225
rect 18103 17191 18119 17225
rect 18053 17183 18119 17191
rect 18153 17361 18195 17377
rect 18187 17327 18195 17361
rect 18153 17293 18195 17327
rect 18187 17259 18195 17293
rect 18153 17225 18195 17259
rect 18187 17191 18195 17225
rect 18153 17149 18195 17191
rect 19044 17349 19102 17384
rect 19044 17315 19056 17349
rect 19090 17315 19102 17349
rect 19044 17256 19102 17315
rect 19044 17222 19056 17256
rect 19090 17222 19102 17256
rect 19044 17151 19102 17222
rect 19175 17381 19221 17428
rect 19255 17429 19271 17463
rect 19305 17458 19321 17463
rect 19255 17424 19281 17429
rect 19315 17424 19321 17458
rect 19255 17415 19321 17424
rect 20049 17436 20051 17470
rect 20085 17436 20095 17470
rect 20817 17493 20883 17505
rect 20917 17607 20963 17653
rect 21365 17651 21394 17685
rect 21428 17651 21486 17685
rect 21520 17651 21578 17685
rect 21612 17651 21670 17685
rect 21704 17651 21733 17685
rect 22149 17653 22178 17687
rect 22212 17653 22268 17687
rect 22302 17653 22360 17687
rect 22394 17653 22452 17687
rect 22486 17653 22515 17687
rect 20951 17573 20963 17607
rect 20917 17539 20963 17573
rect 20951 17505 20963 17539
rect 20817 17466 20863 17493
rect 20917 17489 20963 17505
rect 21431 17605 21497 17617
rect 21431 17571 21447 17605
rect 21481 17571 21497 17605
rect 21431 17537 21497 17571
rect 21431 17503 21447 17537
rect 21481 17503 21497 17537
rect 21431 17491 21497 17503
rect 21531 17605 21577 17651
rect 21565 17571 21577 17605
rect 21531 17537 21577 17571
rect 21565 17503 21577 17537
rect 21658 17557 21716 17651
rect 21658 17523 21670 17557
rect 21704 17523 21716 17557
rect 21658 17506 21716 17523
rect 22166 17559 22224 17653
rect 22166 17525 22178 17559
rect 22212 17525 22224 17559
rect 22166 17508 22224 17525
rect 22305 17607 22371 17619
rect 22305 17573 22321 17607
rect 22355 17573 22371 17607
rect 22305 17539 22371 17573
rect 19175 17363 19241 17381
rect 19175 17329 19191 17363
rect 19225 17329 19241 17363
rect 19175 17295 19241 17329
rect 19175 17261 19191 17295
rect 19225 17261 19241 17295
rect 19175 17227 19241 17261
rect 19175 17193 19191 17227
rect 19225 17193 19241 17227
rect 19175 17185 19241 17193
rect 19275 17363 19317 17379
rect 19309 17329 19317 17363
rect 19275 17295 19317 17329
rect 19309 17261 19317 17295
rect 19275 17227 19317 17261
rect 19309 17193 19317 17227
rect 19275 17151 19317 17193
rect 19910 17351 19968 17386
rect 19910 17317 19922 17351
rect 19956 17317 19968 17351
rect 19910 17258 19968 17317
rect 19910 17224 19922 17258
rect 19956 17224 19968 17258
rect 19910 17153 19968 17224
rect 20049 17383 20095 17436
rect 20129 17462 20145 17465
rect 20129 17428 20141 17462
rect 20179 17428 20195 17465
rect 20129 17417 20195 17428
rect 20817 17432 20823 17466
rect 20861 17432 20863 17466
rect 20049 17365 20115 17383
rect 20049 17331 20065 17365
rect 20099 17331 20115 17365
rect 20049 17297 20115 17331
rect 20049 17263 20065 17297
rect 20099 17263 20115 17297
rect 20049 17229 20115 17263
rect 20049 17195 20065 17229
rect 20099 17195 20115 17229
rect 20049 17187 20115 17195
rect 20149 17365 20191 17381
rect 20183 17331 20191 17365
rect 20149 17297 20191 17331
rect 20183 17263 20191 17297
rect 20149 17229 20191 17263
rect 20183 17195 20191 17229
rect 20149 17153 20191 17195
rect 20680 17341 20738 17376
rect 20680 17307 20692 17341
rect 20726 17307 20738 17341
rect 20680 17248 20738 17307
rect 20680 17214 20692 17248
rect 20726 17214 20738 17248
rect 15481 17085 15510 17119
rect 15544 17085 15596 17119
rect 15630 17085 15688 17119
rect 15722 17085 15780 17119
rect 15814 17085 15843 17119
rect 17911 17115 17940 17149
rect 17974 17115 18016 17149
rect 18050 17115 18108 17149
rect 18142 17115 18200 17149
rect 18234 17115 18263 17149
rect 19027 17117 19056 17151
rect 19090 17117 19138 17151
rect 19172 17117 19230 17151
rect 19264 17117 19322 17151
rect 19356 17117 19385 17151
rect 19893 17119 19922 17153
rect 19956 17119 20012 17153
rect 20046 17119 20104 17153
rect 20138 17119 20196 17153
rect 20230 17119 20259 17153
rect 20680 17143 20738 17214
rect 20817 17373 20863 17432
rect 20897 17454 20913 17455
rect 20897 17420 20911 17454
rect 20947 17420 20963 17455
rect 20897 17407 20963 17420
rect 21431 17452 21477 17491
rect 21531 17487 21577 17503
rect 22305 17505 22321 17539
rect 22355 17505 22371 17539
rect 22305 17493 22371 17505
rect 22405 17607 22451 17653
rect 23007 17643 23036 17677
rect 23070 17643 23128 17677
rect 23162 17643 23220 17677
rect 23254 17643 23310 17677
rect 23344 17643 23373 17677
rect 22439 17573 22451 17607
rect 22405 17539 22451 17573
rect 22439 17505 22451 17539
rect 22305 17460 22351 17493
rect 22405 17489 22451 17505
rect 23073 17597 23139 17609
rect 23073 17563 23089 17597
rect 23123 17563 23139 17597
rect 23073 17529 23139 17563
rect 23073 17495 23089 17529
rect 23123 17495 23139 17529
rect 21431 17418 21433 17452
rect 21469 17418 21477 17452
rect 20817 17355 20883 17373
rect 21431 17371 21477 17418
rect 21511 17419 21527 17453
rect 21561 17448 21577 17453
rect 21511 17414 21537 17419
rect 21571 17414 21577 17448
rect 21511 17405 21577 17414
rect 22305 17426 22307 17460
rect 22341 17426 22351 17460
rect 23073 17483 23139 17495
rect 23173 17597 23219 17643
rect 23207 17563 23219 17597
rect 23173 17529 23219 17563
rect 23207 17495 23219 17529
rect 23298 17549 23356 17643
rect 23298 17515 23310 17549
rect 23344 17515 23356 17549
rect 23298 17498 23356 17515
rect 23073 17456 23119 17483
rect 23173 17479 23219 17495
rect 20817 17321 20833 17355
rect 20867 17321 20883 17355
rect 20817 17287 20883 17321
rect 20817 17253 20833 17287
rect 20867 17253 20883 17287
rect 20817 17219 20883 17253
rect 20817 17185 20833 17219
rect 20867 17185 20883 17219
rect 20817 17177 20883 17185
rect 20917 17355 20959 17371
rect 20951 17321 20959 17355
rect 20917 17287 20959 17321
rect 20951 17253 20959 17287
rect 20917 17219 20959 17253
rect 20951 17185 20959 17219
rect 20917 17143 20959 17185
rect 21431 17353 21497 17371
rect 21431 17319 21447 17353
rect 21481 17319 21497 17353
rect 21431 17285 21497 17319
rect 21431 17251 21447 17285
rect 21481 17251 21497 17285
rect 21431 17217 21497 17251
rect 21431 17183 21447 17217
rect 21481 17183 21497 17217
rect 21431 17175 21497 17183
rect 21531 17353 21573 17369
rect 21565 17319 21573 17353
rect 21531 17285 21573 17319
rect 21565 17251 21573 17285
rect 21531 17217 21573 17251
rect 21565 17183 21573 17217
rect 20663 17109 20692 17143
rect 20726 17109 20780 17143
rect 20814 17109 20872 17143
rect 20906 17109 20964 17143
rect 20998 17109 21027 17143
rect 21531 17141 21573 17183
rect 21658 17339 21716 17374
rect 21658 17305 21670 17339
rect 21704 17305 21716 17339
rect 21658 17246 21716 17305
rect 21658 17212 21670 17246
rect 21704 17212 21716 17246
rect 21658 17141 21716 17212
rect 22166 17341 22224 17376
rect 22166 17307 22178 17341
rect 22212 17307 22224 17341
rect 22166 17248 22224 17307
rect 22166 17214 22178 17248
rect 22212 17214 22224 17248
rect 22166 17143 22224 17214
rect 22305 17373 22351 17426
rect 22385 17452 22401 17455
rect 22385 17418 22397 17452
rect 22435 17418 22451 17455
rect 22385 17407 22451 17418
rect 23073 17422 23079 17456
rect 23117 17422 23119 17456
rect 22305 17355 22371 17373
rect 22305 17321 22321 17355
rect 22355 17321 22371 17355
rect 22305 17287 22371 17321
rect 22305 17253 22321 17287
rect 22355 17253 22371 17287
rect 22305 17219 22371 17253
rect 22305 17185 22321 17219
rect 22355 17185 22371 17219
rect 22305 17177 22371 17185
rect 22405 17355 22447 17371
rect 22439 17321 22447 17355
rect 22405 17287 22447 17321
rect 22439 17253 22447 17287
rect 22405 17219 22447 17253
rect 22439 17185 22447 17219
rect 22405 17143 22447 17185
rect 23073 17363 23119 17422
rect 23153 17444 23169 17445
rect 23153 17410 23167 17444
rect 23203 17410 23219 17445
rect 23153 17397 23219 17410
rect 23073 17345 23139 17363
rect 23073 17311 23089 17345
rect 23123 17311 23139 17345
rect 23073 17277 23139 17311
rect 23073 17243 23089 17277
rect 23123 17243 23139 17277
rect 23073 17209 23139 17243
rect 23073 17175 23089 17209
rect 23123 17175 23139 17209
rect 23073 17167 23139 17175
rect 23173 17345 23215 17361
rect 23207 17311 23215 17345
rect 23173 17277 23215 17311
rect 23207 17243 23215 17277
rect 23173 17209 23215 17243
rect 23207 17175 23215 17209
rect 21365 17107 21394 17141
rect 21428 17107 21486 17141
rect 21520 17107 21578 17141
rect 21612 17107 21670 17141
rect 21704 17107 21733 17141
rect 22149 17109 22178 17143
rect 22212 17109 22268 17143
rect 22302 17109 22360 17143
rect 22394 17109 22452 17143
rect 22486 17109 22515 17143
rect 23173 17133 23215 17175
rect 23298 17331 23356 17366
rect 23298 17297 23310 17331
rect 23344 17297 23356 17331
rect 23298 17238 23356 17297
rect 23298 17204 23310 17238
rect 23344 17204 23356 17238
rect 23298 17133 23356 17204
rect 23007 17099 23036 17133
rect 23070 17099 23128 17133
rect 23162 17099 23220 17133
rect 23254 17099 23310 17133
rect 23344 17099 23373 17133
rect 9334 16573 9363 16607
rect 9397 16573 9455 16607
rect 9489 16573 9547 16607
rect 9581 16573 9639 16607
rect 9673 16573 9731 16607
rect 9765 16573 9823 16607
rect 9857 16573 9915 16607
rect 9949 16573 9978 16607
rect 9351 16531 9427 16539
rect 9351 16497 9377 16531
rect 9411 16497 9427 16531
rect 9351 16463 9427 16497
rect 9351 16429 9377 16463
rect 9411 16429 9427 16463
rect 9351 16403 9427 16429
rect 9545 16521 9579 16573
rect 9545 16453 9579 16487
rect 9545 16403 9579 16419
rect 9613 16521 9679 16539
rect 9613 16487 9629 16521
rect 9663 16487 9679 16521
rect 9613 16453 9679 16487
rect 9713 16521 9747 16573
rect 9713 16471 9747 16487
rect 9781 16521 9861 16539
rect 9781 16487 9817 16521
rect 9851 16487 9861 16521
rect 9613 16419 9629 16453
rect 9663 16437 9679 16453
rect 9781 16453 9861 16487
rect 9781 16437 9817 16453
rect 9663 16419 9817 16437
rect 9851 16419 9861 16453
rect 9613 16403 9861 16419
rect 9897 16523 9961 16539
rect 9897 16489 9901 16523
rect 9935 16489 9961 16523
rect 9897 16455 9961 16489
rect 9897 16421 9901 16455
rect 9935 16421 9961 16455
rect 9351 16211 9385 16403
rect 9897 16394 9961 16421
rect 9897 16387 9910 16394
rect 9419 16335 9680 16369
rect 9897 16353 9901 16387
rect 9944 16356 9961 16394
rect 9935 16353 9961 16356
rect 9419 16296 9468 16335
rect 9419 16295 9420 16296
rect 9454 16262 9468 16296
rect 9453 16261 9468 16262
rect 9502 16298 9612 16301
rect 9502 16295 9540 16298
rect 9502 16261 9536 16295
rect 9574 16264 9612 16298
rect 9570 16261 9612 16264
rect 9646 16295 9680 16335
rect 9835 16319 9961 16353
rect 9755 16295 9801 16311
rect 9646 16261 9671 16295
rect 9705 16261 9721 16295
rect 9755 16261 9767 16295
rect 9419 16245 9468 16261
rect 9755 16211 9801 16261
rect 9351 16177 9801 16211
rect 9461 16163 9495 16177
rect 9361 16107 9377 16141
rect 9411 16107 9427 16141
rect 9835 16143 9869 16319
rect 9461 16113 9495 16129
rect 9361 16063 9427 16107
rect 9529 16107 9545 16141
rect 9579 16107 9595 16141
rect 9678 16109 9713 16143
rect 9747 16109 9813 16143
rect 9847 16109 9869 16143
rect 9903 16214 9961 16230
rect 9937 16180 9961 16214
rect 9903 16146 9961 16180
rect 9937 16112 9961 16146
rect 9529 16063 9595 16107
rect 9903 16063 9961 16112
rect 9334 16029 9363 16063
rect 9397 16029 9455 16063
rect 9489 16029 9547 16063
rect 9581 16029 9639 16063
rect 9673 16029 9731 16063
rect 9765 16029 9823 16063
rect 9857 16029 9915 16063
rect 9949 16029 9978 16063
rect 9432 15829 9461 15863
rect 9495 15829 9553 15863
rect 9587 15829 9645 15863
rect 9679 15829 9737 15863
rect 9771 15829 9829 15863
rect 9863 15829 9892 15863
rect 9489 15745 9545 15829
rect 9679 15787 9745 15829
rect 9489 15711 9503 15745
rect 9537 15711 9545 15745
rect 9489 15695 9545 15711
rect 9579 15745 9639 15761
rect 9579 15711 9587 15745
rect 9621 15711 9639 15745
rect 9579 15651 9639 15711
rect 9679 15753 9695 15787
rect 9729 15753 9745 15787
rect 9679 15719 9745 15753
rect 9679 15685 9695 15719
rect 9729 15685 9745 15719
rect 9783 15787 9875 15795
rect 9783 15753 9799 15787
rect 9833 15753 9875 15787
rect 9783 15719 9875 15753
rect 11474 15719 11503 15753
rect 11537 15719 11595 15753
rect 11629 15719 11687 15753
rect 11721 15719 11779 15753
rect 11813 15719 11871 15753
rect 11905 15719 11963 15753
rect 11997 15719 12055 15753
rect 12089 15719 12118 15753
rect 9783 15685 9799 15719
rect 9833 15685 9875 15719
rect 9452 15574 9505 15639
rect 9579 15617 9767 15651
rect 9452 15534 9454 15574
rect 9496 15567 9505 15574
rect 9733 15567 9767 15617
rect 9496 15551 9587 15567
rect 9496 15534 9506 15551
rect 9452 15517 9506 15534
rect 9540 15517 9587 15551
rect 9631 15564 9699 15567
rect 9631 15524 9644 15564
rect 9686 15524 9699 15564
rect 9631 15517 9647 15524
rect 9681 15517 9699 15524
rect 9733 15551 9791 15567
rect 9733 15517 9755 15551
rect 9789 15517 9791 15551
rect 9733 15501 9791 15517
rect 9733 15483 9767 15501
rect 9489 15445 9767 15483
rect 9825 15494 9875 15685
rect 11492 15677 11559 15719
rect 11492 15643 11509 15677
rect 11543 15643 11559 15677
rect 11593 15669 11643 15685
rect 11593 15635 11601 15669
rect 11635 15635 11643 15669
rect 9825 15460 9836 15494
rect 9872 15460 9875 15494
rect 9489 15423 9555 15445
rect 9489 15389 9503 15423
rect 9537 15389 9555 15423
rect 9825 15411 9875 15460
rect 9489 15373 9555 15389
rect 9679 15395 9729 15411
rect 9679 15361 9695 15395
rect 9679 15319 9729 15361
rect 9763 15395 9875 15411
rect 9763 15361 9779 15395
rect 9813 15361 9875 15395
rect 9763 15353 9875 15361
rect 11491 15441 11539 15607
rect 11593 15525 11643 15635
rect 11687 15677 11753 15719
rect 11687 15643 11703 15677
rect 11737 15643 11753 15677
rect 11687 15575 11753 15643
rect 11790 15669 11840 15685
rect 11790 15635 11798 15669
rect 11832 15635 11840 15669
rect 11790 15525 11840 15635
rect 11933 15677 11999 15719
rect 11933 15643 11949 15677
rect 11983 15643 11999 15677
rect 11933 15609 11999 15643
rect 12033 15677 12101 15685
rect 12033 15643 12049 15677
rect 12083 15643 12101 15677
rect 12033 15633 12101 15643
rect 11933 15575 11949 15609
rect 11983 15575 11999 15609
rect 11933 15559 11999 15575
rect 12049 15609 12101 15633
rect 12083 15575 12101 15609
rect 12049 15541 12101 15575
rect 11491 15407 11505 15441
rect 11491 15404 11539 15407
rect 11491 15368 11498 15404
rect 11534 15368 11539 15404
rect 11491 15345 11539 15368
rect 11573 15491 12011 15525
rect 9432 15285 9461 15319
rect 9495 15285 9553 15319
rect 9587 15285 9645 15319
rect 9679 15285 9737 15319
rect 9771 15285 9829 15319
rect 9863 15285 9892 15319
rect 11573 15309 11607 15491
rect 11948 15457 12011 15491
rect 12083 15507 12101 15541
rect 11508 15293 11607 15309
rect 11508 15259 11509 15293
rect 11543 15259 11607 15293
rect 11651 15441 11721 15457
rect 11685 15438 11721 15441
rect 11651 15402 11670 15407
rect 11704 15402 11721 15438
rect 11651 15264 11721 15402
rect 11757 15441 11817 15457
rect 11791 15407 11817 15441
rect 11757 15314 11817 15407
rect 11757 15280 11768 15314
rect 11802 15280 11817 15314
rect 11757 15263 11817 15280
rect 11853 15441 11909 15457
rect 11887 15407 11909 15441
rect 11948 15441 12014 15457
rect 11948 15407 11964 15441
rect 11998 15407 12014 15441
rect 12049 15436 12101 15507
rect 11853 15384 11909 15407
rect 11853 15348 11864 15384
rect 11898 15348 11909 15384
rect 12049 15402 12056 15436
rect 12090 15402 12101 15436
rect 11853 15263 11909 15348
rect 11945 15353 11999 15369
rect 12049 15353 12101 15402
rect 11945 15319 11950 15353
rect 11984 15319 11999 15353
rect 11945 15285 11999 15319
rect 10616 15219 10645 15253
rect 10679 15219 10737 15253
rect 10771 15219 10829 15253
rect 10863 15219 10921 15253
rect 10955 15219 11013 15253
rect 11047 15219 11076 15253
rect 11508 15243 11607 15259
rect 11945 15251 11950 15285
rect 11984 15251 11999 15285
rect 12033 15319 12049 15353
rect 12083 15319 12101 15353
rect 12033 15285 12101 15319
rect 12033 15251 12049 15285
rect 12083 15251 12101 15285
rect 10673 15135 10729 15219
rect 10863 15177 10929 15219
rect 11945 15209 11999 15251
rect 10673 15101 10687 15135
rect 10721 15101 10729 15135
rect 10673 15085 10729 15101
rect 10763 15135 10823 15151
rect 10763 15101 10771 15135
rect 10805 15101 10823 15135
rect 9344 15009 9373 15043
rect 9407 15009 9465 15043
rect 9499 15009 9557 15043
rect 9591 15009 9649 15043
rect 9683 15009 9741 15043
rect 9775 15009 9833 15043
rect 9867 15009 9925 15043
rect 9959 15009 9988 15043
rect 10763 15041 10823 15101
rect 10863 15143 10879 15177
rect 10913 15143 10929 15177
rect 10863 15109 10929 15143
rect 10863 15075 10879 15109
rect 10913 15075 10929 15109
rect 10967 15177 11059 15185
rect 10967 15143 10983 15177
rect 11017 15152 11059 15177
rect 11474 15175 11503 15209
rect 11537 15175 11595 15209
rect 11629 15175 11687 15209
rect 11721 15175 11779 15209
rect 11813 15175 11871 15209
rect 11905 15175 11963 15209
rect 11997 15175 12055 15209
rect 12089 15175 12118 15209
rect 10967 15116 11010 15143
rect 11050 15116 11059 15152
rect 10967 15109 11059 15116
rect 10967 15075 10983 15109
rect 11017 15075 11059 15109
rect 9361 14967 9437 14975
rect 9361 14933 9387 14967
rect 9421 14933 9437 14967
rect 9361 14899 9437 14933
rect 9361 14865 9387 14899
rect 9421 14865 9437 14899
rect 9361 14839 9437 14865
rect 9555 14957 9589 15009
rect 9555 14889 9589 14923
rect 9555 14839 9589 14855
rect 9623 14957 9689 14975
rect 9623 14923 9639 14957
rect 9673 14923 9689 14957
rect 9623 14889 9689 14923
rect 9723 14957 9757 15009
rect 9723 14907 9757 14923
rect 9791 14957 9871 14975
rect 9791 14923 9827 14957
rect 9861 14923 9871 14957
rect 9623 14855 9639 14889
rect 9673 14873 9689 14889
rect 9791 14889 9871 14923
rect 9791 14873 9827 14889
rect 9673 14855 9827 14873
rect 9861 14855 9871 14889
rect 9623 14839 9871 14855
rect 9907 14959 9971 14975
rect 9907 14925 9911 14959
rect 9945 14934 9971 14959
rect 9907 14900 9922 14925
rect 9956 14900 9971 14934
rect 10636 14957 10689 15029
rect 10763 15007 10951 15041
rect 10917 14957 10951 15007
rect 10636 14942 10771 14957
rect 10636 14907 10690 14942
rect 10724 14907 10771 14942
rect 10815 14942 10883 14957
rect 10815 14908 10830 14942
rect 10866 14908 10883 14942
rect 10815 14907 10831 14908
rect 10865 14907 10883 14908
rect 10917 14941 10975 14957
rect 10917 14907 10939 14941
rect 10973 14907 10975 14941
rect 9907 14891 9971 14900
rect 9907 14857 9911 14891
rect 9945 14857 9971 14891
rect 10917 14891 10975 14907
rect 10917 14873 10951 14891
rect 9361 14647 9395 14839
rect 9907 14823 9971 14857
rect 9429 14771 9690 14805
rect 9907 14789 9911 14823
rect 9945 14789 9971 14823
rect 9429 14732 9478 14771
rect 9429 14731 9430 14732
rect 9464 14698 9478 14732
rect 9463 14697 9478 14698
rect 9512 14734 9622 14737
rect 9512 14731 9550 14734
rect 9512 14697 9546 14731
rect 9584 14700 9622 14734
rect 9580 14697 9622 14700
rect 9656 14731 9690 14771
rect 9845 14755 9971 14789
rect 10673 14835 10951 14873
rect 10673 14813 10739 14835
rect 10673 14779 10687 14813
rect 10721 14779 10739 14813
rect 11009 14801 11059 15075
rect 10673 14763 10739 14779
rect 10863 14785 10913 14801
rect 9765 14731 9811 14747
rect 9656 14697 9681 14731
rect 9715 14697 9731 14731
rect 9765 14697 9777 14731
rect 9429 14681 9478 14697
rect 9765 14647 9811 14697
rect 9361 14613 9811 14647
rect 9471 14599 9505 14613
rect 9371 14543 9387 14577
rect 9421 14543 9437 14577
rect 9845 14579 9879 14755
rect 10863 14751 10879 14785
rect 10863 14709 10913 14751
rect 10947 14785 11059 14801
rect 10947 14751 10963 14785
rect 10997 14751 11059 14785
rect 10947 14743 11059 14751
rect 10616 14675 10645 14709
rect 10679 14675 10737 14709
rect 10771 14675 10829 14709
rect 10863 14675 10921 14709
rect 10955 14675 11013 14709
rect 11047 14675 11076 14709
rect 9471 14549 9505 14565
rect 9371 14499 9437 14543
rect 9539 14543 9555 14577
rect 9589 14543 9605 14577
rect 9688 14545 9723 14579
rect 9757 14545 9823 14579
rect 9857 14545 9879 14579
rect 9913 14650 9971 14666
rect 9947 14616 9971 14650
rect 9913 14582 9971 14616
rect 9947 14548 9971 14582
rect 9539 14499 9605 14543
rect 9913 14499 9971 14548
rect 9344 14465 9373 14499
rect 9407 14465 9465 14499
rect 9499 14465 9557 14499
rect 9591 14465 9649 14499
rect 9683 14465 9741 14499
rect 9775 14465 9833 14499
rect 9867 14465 9925 14499
rect 9959 14465 9988 14499
rect 9442 14265 9471 14299
rect 9505 14265 9563 14299
rect 9597 14265 9655 14299
rect 9689 14265 9747 14299
rect 9781 14265 9839 14299
rect 9873 14265 9902 14299
rect 9499 14181 9555 14265
rect 9689 14223 9755 14265
rect 10690 14253 10719 14287
rect 10753 14253 10811 14287
rect 10845 14253 10903 14287
rect 10937 14253 10995 14287
rect 11029 14253 11087 14287
rect 11121 14253 11179 14287
rect 11213 14253 11271 14287
rect 11305 14253 11334 14287
rect 9499 14147 9513 14181
rect 9547 14147 9555 14181
rect 9499 14131 9555 14147
rect 9589 14181 9649 14197
rect 9589 14147 9597 14181
rect 9631 14147 9649 14181
rect 9589 14087 9649 14147
rect 9689 14189 9705 14223
rect 9739 14189 9755 14223
rect 9689 14155 9755 14189
rect 9689 14121 9705 14155
rect 9739 14121 9755 14155
rect 9793 14223 9885 14231
rect 9793 14189 9809 14223
rect 9843 14189 9885 14223
rect 9793 14155 9885 14189
rect 10708 14211 10775 14253
rect 10708 14177 10725 14211
rect 10759 14177 10775 14211
rect 10809 14203 10859 14219
rect 9793 14121 9809 14155
rect 9843 14121 9885 14155
rect 10809 14169 10817 14203
rect 10851 14169 10859 14203
rect 9462 14010 9515 14075
rect 9589 14053 9777 14087
rect 9462 13970 9464 14010
rect 9506 14003 9515 14010
rect 9743 14003 9777 14053
rect 9506 13987 9597 14003
rect 9506 13970 9516 13987
rect 9462 13953 9516 13970
rect 9550 13953 9597 13987
rect 9641 14000 9709 14003
rect 9641 13960 9654 14000
rect 9696 13960 9709 14000
rect 9641 13953 9657 13960
rect 9691 13953 9709 13960
rect 9743 13987 9801 14003
rect 9743 13953 9765 13987
rect 9799 13953 9801 13987
rect 9743 13937 9801 13953
rect 9743 13919 9777 13937
rect 9499 13881 9777 13919
rect 9835 13888 9885 14121
rect 9499 13859 9565 13881
rect 9499 13825 9513 13859
rect 9547 13825 9565 13859
rect 9835 13854 9844 13888
rect 9880 13854 9885 13888
rect 10707 13980 10755 14141
rect 10809 14059 10859 14169
rect 10903 14211 10969 14253
rect 10903 14177 10919 14211
rect 10953 14177 10969 14211
rect 10903 14109 10969 14177
rect 11006 14203 11056 14219
rect 11006 14169 11014 14203
rect 11048 14169 11056 14203
rect 11006 14059 11056 14169
rect 11149 14211 11215 14253
rect 12588 14237 12617 14271
rect 12651 14237 12709 14271
rect 12743 14237 12801 14271
rect 12835 14237 12893 14271
rect 12927 14237 12985 14271
rect 13019 14237 13077 14271
rect 13111 14237 13140 14271
rect 11149 14177 11165 14211
rect 11199 14177 11215 14211
rect 11149 14143 11215 14177
rect 11249 14211 11317 14219
rect 11249 14177 11265 14211
rect 11299 14177 11317 14211
rect 12971 14195 13027 14237
rect 11249 14167 11317 14177
rect 11149 14109 11165 14143
rect 11199 14109 11215 14143
rect 11149 14093 11215 14109
rect 11265 14143 11317 14167
rect 11299 14109 11317 14143
rect 12606 14183 12937 14193
rect 12606 14170 12845 14183
rect 12606 14136 12762 14170
rect 12798 14149 12845 14170
rect 12879 14149 12937 14183
rect 12798 14136 12937 14149
rect 12606 14135 12937 14136
rect 12971 14161 12984 14195
rect 13018 14161 13027 14195
rect 11265 14075 11317 14109
rect 12971 14127 13027 14161
rect 10707 13946 10716 13980
rect 10750 13975 10755 13980
rect 10707 13941 10721 13946
rect 10707 13879 10755 13941
rect 10789 14025 11227 14059
rect 9835 13847 9885 13854
rect 9499 13809 9565 13825
rect 9689 13831 9739 13847
rect 9689 13797 9705 13831
rect 9689 13755 9739 13797
rect 9773 13831 9885 13847
rect 10789 13843 10823 14025
rect 11164 13991 11227 14025
rect 11299 14041 11317 14075
rect 9773 13797 9789 13831
rect 9823 13797 9885 13831
rect 9773 13789 9885 13797
rect 10724 13827 10823 13843
rect 10724 13793 10725 13827
rect 10759 13793 10823 13827
rect 10867 13975 10937 13991
rect 10901 13941 10937 13975
rect 10867 13884 10937 13941
rect 10867 13850 10886 13884
rect 10920 13850 10937 13884
rect 10867 13798 10937 13850
rect 10973 13975 11033 13991
rect 11007 13941 11033 13975
rect 10973 13924 11033 13941
rect 10973 13890 10984 13924
rect 11018 13890 11033 13924
rect 10973 13797 11033 13890
rect 11069 13975 11125 13991
rect 11103 13974 11125 13975
rect 11069 13936 11078 13941
rect 11114 13936 11125 13974
rect 11164 13975 11230 13991
rect 11164 13941 11180 13975
rect 11214 13941 11230 13975
rect 11069 13797 11125 13936
rect 11161 13887 11215 13903
rect 11265 13887 11317 14041
rect 12606 14067 12924 14101
rect 12971 14093 12984 14127
rect 13018 14093 13027 14127
rect 12971 14077 13027 14093
rect 13069 14164 13123 14203
rect 13103 14130 13123 14164
rect 13069 14096 13123 14130
rect 13103 14080 13123 14096
rect 12606 14064 12670 14067
rect 12606 14030 12623 14064
rect 12657 14030 12670 14064
rect 12890 14043 12924 14067
rect 12606 14009 12670 14030
rect 12606 13959 12676 13975
rect 12606 13942 12623 13959
rect 12657 13942 12676 13959
rect 11161 13853 11166 13887
rect 11200 13853 11215 13887
rect 11161 13819 11215 13853
rect 10724 13777 10823 13793
rect 11161 13785 11166 13819
rect 11200 13785 11215 13819
rect 11249 13856 11265 13887
rect 11249 13818 11260 13856
rect 11299 13853 11317 13887
rect 11660 13879 11689 13913
rect 11723 13879 11781 13913
rect 11815 13879 11873 13913
rect 11907 13879 11965 13913
rect 11999 13879 12057 13913
rect 12091 13879 12120 13913
rect 12606 13908 12618 13942
rect 12658 13908 12676 13942
rect 12710 13964 12852 14033
rect 12890 14009 13035 14043
rect 13069 14040 13078 14062
rect 13120 14040 13123 14080
rect 13069 14009 13123 14040
rect 13001 13975 13035 14009
rect 12710 13922 12746 13964
rect 12796 13922 12852 13964
rect 12710 13909 12852 13922
rect 12886 13960 12967 13975
rect 12886 13924 12918 13960
rect 12956 13959 12967 13960
rect 12959 13925 12967 13959
rect 12956 13924 12967 13925
rect 12886 13909 12967 13924
rect 13001 13959 13055 13975
rect 13001 13925 13021 13959
rect 13001 13909 13055 13925
rect 11298 13819 11317 13853
rect 11249 13785 11265 13818
rect 11299 13785 11317 13819
rect 11889 13821 11955 13879
rect 12606 13861 12676 13908
rect 13001 13875 13035 13909
rect 11889 13787 11905 13821
rect 11939 13787 11955 13821
rect 9442 13721 9471 13755
rect 9505 13721 9563 13755
rect 9597 13721 9655 13755
rect 9689 13721 9747 13755
rect 9781 13721 9839 13755
rect 9873 13721 9902 13755
rect 11161 13743 11215 13785
rect 11889 13753 11955 13787
rect 10690 13709 10719 13743
rect 10753 13709 10811 13743
rect 10845 13709 10903 13743
rect 10937 13709 10995 13743
rect 11029 13709 11087 13743
rect 11121 13709 11179 13743
rect 11213 13709 11271 13743
rect 11305 13709 11334 13743
rect 11714 13701 11792 13720
rect 11889 13719 11905 13753
rect 11939 13719 11955 13753
rect 11989 13837 12096 13845
rect 11989 13803 12005 13837
rect 12039 13803 12096 13837
rect 12713 13841 13035 13875
rect 13089 13862 13123 14009
rect 13069 13845 13123 13862
rect 11989 13769 12096 13803
rect 11989 13735 12005 13769
rect 12039 13768 12096 13769
rect 11989 13734 12028 13735
rect 12062 13734 12096 13768
rect 11989 13721 12096 13734
rect 12607 13793 12623 13827
rect 12657 13793 12673 13827
rect 12607 13727 12673 13793
rect 12713 13821 12747 13841
rect 12887 13821 12921 13841
rect 12713 13771 12747 13787
rect 12787 13773 12803 13807
rect 12837 13773 12853 13807
rect 12787 13727 12853 13773
rect 13103 13811 13123 13845
rect 12887 13771 12921 13787
rect 12955 13773 12981 13807
rect 13015 13773 13031 13807
rect 13069 13793 13123 13811
rect 12955 13727 13031 13773
rect 11714 13667 11736 13701
rect 11770 13685 11792 13701
rect 11770 13667 11999 13685
rect 11714 13651 11999 13667
rect 11689 13601 11760 13617
rect 11689 13567 11726 13601
rect 11689 13558 11760 13567
rect 11689 13524 11700 13558
rect 11734 13524 11760 13558
rect 11689 13505 11760 13524
rect 11794 13471 11828 13651
rect 11862 13608 11915 13617
rect 11862 13601 11878 13608
rect 11912 13574 11915 13608
rect 11896 13567 11915 13574
rect 11862 13505 11915 13567
rect 11965 13601 11999 13651
rect 11965 13551 11999 13567
rect 12033 13517 12096 13721
rect 12588 13693 12617 13727
rect 12651 13693 12709 13727
rect 12743 13693 12801 13727
rect 12835 13693 12893 13727
rect 12927 13693 12985 13727
rect 13019 13693 13077 13727
rect 13111 13693 13140 13727
rect 11973 13515 12096 13517
rect 11973 13481 11989 13515
rect 12023 13481 12096 13515
rect 11710 13455 11758 13471
rect 10814 13411 10843 13445
rect 10877 13411 10935 13445
rect 10969 13411 11027 13445
rect 11061 13411 11119 13445
rect 11153 13411 11211 13445
rect 11245 13411 11274 13445
rect 11710 13421 11724 13455
rect 9336 13341 9365 13375
rect 9399 13341 9457 13375
rect 9491 13341 9549 13375
rect 9583 13341 9641 13375
rect 9675 13341 9733 13375
rect 9767 13341 9825 13375
rect 9859 13341 9917 13375
rect 9951 13341 9980 13375
rect 9353 13299 9429 13307
rect 9353 13265 9379 13299
rect 9413 13265 9429 13299
rect 9353 13231 9429 13265
rect 9353 13197 9379 13231
rect 9413 13197 9429 13231
rect 9353 13171 9429 13197
rect 9547 13289 9581 13341
rect 9547 13221 9581 13255
rect 9547 13171 9581 13187
rect 9615 13289 9681 13307
rect 9615 13255 9631 13289
rect 9665 13255 9681 13289
rect 9615 13221 9681 13255
rect 9715 13289 9749 13341
rect 9715 13239 9749 13255
rect 9783 13289 9863 13307
rect 9783 13255 9819 13289
rect 9853 13255 9863 13289
rect 9615 13187 9631 13221
rect 9665 13205 9681 13221
rect 9783 13221 9863 13255
rect 9783 13205 9819 13221
rect 9665 13187 9819 13205
rect 9853 13187 9863 13221
rect 9615 13171 9863 13187
rect 9899 13291 9963 13307
rect 9899 13257 9903 13291
rect 9937 13257 9963 13291
rect 10831 13300 10952 13411
rect 10987 13360 11083 13377
rect 11021 13338 11083 13360
rect 10987 13309 11012 13326
rect 11048 13309 11083 13338
rect 11117 13369 11168 13411
rect 11117 13335 11121 13369
rect 11155 13335 11168 13369
rect 11117 13302 11168 13335
rect 11202 13355 11257 13377
rect 11710 13369 11758 13421
rect 11794 13455 11850 13471
rect 11794 13421 11808 13455
rect 11842 13421 11850 13455
rect 11794 13405 11850 13421
rect 11896 13455 11939 13471
rect 11896 13421 11904 13455
rect 11938 13421 11939 13455
rect 11896 13369 11939 13421
rect 11973 13447 12096 13481
rect 11973 13413 11989 13447
rect 12023 13413 12096 13447
rect 11973 13403 12096 13413
rect 11202 13321 11205 13355
rect 11239 13321 11257 13355
rect 11660 13335 11689 13369
rect 11723 13335 11781 13369
rect 11815 13335 11873 13369
rect 11907 13335 11965 13369
rect 11999 13335 12057 13369
rect 12091 13335 12120 13369
rect 10831 13280 10954 13300
rect 9899 13224 9963 13257
rect 10917 13275 10954 13280
rect 11202 13287 11257 13321
rect 10917 13260 10983 13275
rect 9899 13223 9914 13224
rect 9899 13189 9903 13223
rect 9948 13190 9963 13224
rect 9937 13189 9963 13190
rect 9353 12979 9387 13171
rect 9899 13155 9963 13189
rect 9421 13103 9682 13137
rect 9899 13121 9903 13155
rect 9937 13121 9963 13155
rect 10831 13230 10883 13246
rect 10831 13196 10849 13230
rect 10917 13226 10933 13260
rect 10967 13226 10983 13260
rect 11017 13241 11168 13261
rect 11017 13211 11026 13241
rect 11014 13207 11026 13211
rect 11060 13207 11168 13241
rect 11202 13253 11205 13287
rect 11239 13282 11257 13287
rect 11202 13244 11208 13253
rect 11246 13244 11257 13282
rect 11202 13237 11257 13244
rect 11014 13204 11168 13207
rect 11011 13202 11168 13204
rect 11010 13199 11189 13202
rect 11006 13196 11189 13199
rect 10831 13156 10883 13196
rect 11002 13194 11189 13196
rect 10997 13192 11189 13194
rect 10983 13186 11189 13192
rect 10979 13180 11189 13186
rect 10975 13174 11189 13180
rect 10969 13169 11189 13174
rect 10962 13162 11189 13169
rect 10956 13161 11189 13162
rect 10956 13160 11034 13161
rect 10956 13158 11029 13160
rect 10956 13157 11026 13158
rect 10956 13156 11023 13157
rect 10831 13155 11023 13156
rect 10831 13153 11021 13155
rect 10831 13152 11019 13153
rect 10831 13150 11017 13152
rect 10831 13148 11016 13150
rect 10831 13147 11015 13148
rect 10831 13144 11013 13147
rect 10831 13141 11012 13144
rect 10831 13136 11010 13141
rect 10831 13122 11009 13136
rect 11143 13133 11189 13161
rect 9421 13064 9470 13103
rect 9421 13063 9422 13064
rect 9456 13030 9470 13064
rect 9455 13029 9470 13030
rect 9504 13066 9614 13069
rect 9504 13063 9542 13066
rect 9504 13029 9538 13063
rect 9576 13032 9614 13066
rect 9572 13029 9614 13032
rect 9648 13063 9682 13103
rect 9837 13087 9963 13121
rect 10831 13087 10941 13088
rect 9757 13063 9803 13079
rect 9648 13029 9673 13063
rect 9707 13029 9723 13063
rect 9757 13029 9769 13063
rect 9421 13013 9470 13029
rect 9757 12979 9803 13029
rect 9353 12945 9803 12979
rect 9463 12931 9497 12945
rect 9363 12875 9379 12909
rect 9413 12875 9429 12909
rect 9837 12911 9871 13087
rect 10831 13053 10849 13087
rect 10883 13064 10941 13087
rect 10831 13030 10860 13053
rect 10894 13030 10941 13064
rect 10831 13011 10941 13030
rect 9463 12881 9497 12897
rect 9363 12831 9429 12875
rect 9531 12875 9547 12909
rect 9581 12875 9597 12909
rect 9680 12877 9715 12911
rect 9749 12877 9815 12911
rect 9849 12877 9871 12911
rect 9905 12982 9963 12998
rect 9939 12948 9963 12982
rect 10975 12977 11009 13122
rect 9905 12914 9963 12948
rect 10831 12943 10849 12977
rect 10883 12943 11009 12977
rect 11043 13093 11059 13127
rect 11093 13093 11109 13127
rect 11043 13070 11109 13093
rect 11143 13099 11155 13133
rect 11143 13082 11189 13099
rect 11043 13036 11062 13070
rect 11098 13042 11109 13070
rect 11043 12945 11087 13036
rect 11223 13031 11257 13237
rect 11121 12993 11171 13009
rect 11155 12959 11171 12993
rect 9939 12880 9963 12914
rect 11121 12901 11171 12959
rect 11205 13003 11257 13031
rect 11239 12969 11257 13003
rect 11205 12935 11257 12969
rect 9531 12831 9597 12875
rect 9905 12831 9963 12880
rect 10814 12867 10843 12901
rect 10877 12867 10935 12901
rect 10969 12867 11027 12901
rect 11061 12867 11119 12901
rect 11153 12867 11211 12901
rect 11245 12867 11274 12901
rect 9336 12797 9365 12831
rect 9399 12797 9457 12831
rect 9491 12797 9549 12831
rect 9583 12797 9641 12831
rect 9675 12797 9733 12831
rect 9767 12797 9825 12831
rect 9859 12797 9917 12831
rect 9951 12797 9980 12831
rect 9434 12597 9463 12631
rect 9497 12597 9555 12631
rect 9589 12597 9647 12631
rect 9681 12597 9739 12631
rect 9773 12597 9831 12631
rect 9865 12597 9894 12631
rect 9491 12513 9547 12597
rect 9681 12555 9747 12597
rect 9491 12479 9505 12513
rect 9539 12479 9547 12513
rect 9491 12463 9547 12479
rect 9581 12513 9641 12529
rect 9581 12479 9589 12513
rect 9623 12479 9641 12513
rect 9581 12419 9641 12479
rect 9681 12521 9697 12555
rect 9731 12521 9747 12555
rect 9681 12487 9747 12521
rect 9681 12453 9697 12487
rect 9731 12453 9747 12487
rect 9785 12555 9877 12563
rect 9785 12521 9801 12555
rect 9835 12521 9877 12555
rect 9785 12487 9877 12521
rect 9785 12453 9801 12487
rect 9835 12453 9877 12487
rect 9454 12342 9507 12407
rect 9581 12385 9769 12419
rect 9454 12302 9456 12342
rect 9498 12335 9507 12342
rect 9735 12335 9769 12385
rect 9827 12374 9877 12453
rect 10810 12391 10839 12425
rect 10873 12391 10931 12425
rect 10965 12391 11023 12425
rect 11057 12391 11115 12425
rect 11149 12391 11207 12425
rect 11241 12391 11270 12425
rect 9827 12340 9836 12374
rect 9872 12340 9877 12374
rect 9498 12319 9589 12335
rect 9498 12302 9508 12319
rect 9454 12285 9508 12302
rect 9542 12285 9589 12319
rect 9633 12332 9701 12335
rect 9633 12292 9646 12332
rect 9688 12292 9701 12332
rect 9633 12285 9649 12292
rect 9683 12285 9701 12292
rect 9735 12319 9793 12335
rect 9735 12285 9757 12319
rect 9791 12285 9793 12319
rect 9735 12269 9793 12285
rect 9735 12251 9769 12269
rect 9491 12213 9769 12251
rect 9491 12191 9557 12213
rect 9491 12157 9505 12191
rect 9539 12157 9557 12191
rect 9827 12179 9877 12340
rect 10867 12307 10923 12391
rect 11057 12349 11123 12391
rect 10867 12273 10881 12307
rect 10915 12273 10923 12307
rect 10867 12257 10923 12273
rect 10957 12307 11017 12323
rect 10957 12273 10965 12307
rect 10999 12273 11017 12307
rect 10957 12213 11017 12273
rect 11057 12315 11073 12349
rect 11107 12315 11123 12349
rect 11057 12281 11123 12315
rect 11057 12247 11073 12281
rect 11107 12247 11123 12281
rect 11161 12349 11253 12357
rect 11161 12315 11177 12349
rect 11211 12315 11253 12349
rect 11161 12281 11253 12315
rect 11161 12247 11177 12281
rect 11211 12247 11253 12281
rect 9491 12141 9557 12157
rect 9681 12163 9731 12179
rect 9681 12129 9697 12163
rect 9681 12087 9731 12129
rect 9765 12163 9877 12179
rect 9765 12129 9781 12163
rect 9815 12129 9877 12163
rect 9765 12121 9877 12129
rect 10830 12129 10883 12201
rect 10957 12179 11145 12213
rect 11111 12129 11145 12179
rect 11203 12200 11253 12247
rect 11203 12166 11212 12200
rect 11246 12166 11253 12200
rect 10830 12116 10965 12129
rect 9434 12053 9463 12087
rect 9497 12053 9555 12087
rect 9589 12053 9647 12087
rect 9681 12053 9739 12087
rect 9773 12053 9831 12087
rect 9865 12053 9894 12087
rect 10830 12079 10884 12116
rect 10920 12082 10965 12116
rect 10918 12079 10965 12082
rect 11009 12114 11077 12129
rect 11009 12080 11024 12114
rect 11060 12080 11077 12114
rect 11009 12079 11025 12080
rect 11059 12079 11077 12080
rect 11111 12113 11169 12129
rect 11111 12079 11133 12113
rect 11167 12079 11169 12113
rect 11111 12063 11169 12079
rect 11111 12045 11145 12063
rect 10867 12007 11145 12045
rect 10867 11985 10933 12007
rect 10867 11951 10881 11985
rect 10915 11951 10933 11985
rect 11203 11973 11253 12166
rect 10867 11935 10933 11951
rect 11057 11957 11107 11973
rect 11057 11923 11073 11957
rect 11057 11881 11107 11923
rect 11141 11957 11253 11973
rect 11141 11923 11157 11957
rect 11191 11923 11253 11957
rect 11141 11915 11253 11923
rect 10810 11847 10839 11881
rect 10873 11847 10931 11881
rect 10965 11847 11023 11881
rect 11057 11847 11115 11881
rect 11149 11847 11207 11881
rect 11241 11847 11270 11881
rect 9346 11777 9375 11811
rect 9409 11777 9467 11811
rect 9501 11777 9559 11811
rect 9593 11777 9651 11811
rect 9685 11777 9743 11811
rect 9777 11777 9835 11811
rect 9869 11777 9927 11811
rect 9961 11777 9990 11811
rect 9363 11735 9439 11743
rect 9363 11701 9389 11735
rect 9423 11701 9439 11735
rect 9363 11667 9439 11701
rect 9363 11633 9389 11667
rect 9423 11633 9439 11667
rect 9363 11607 9439 11633
rect 9557 11725 9591 11777
rect 9557 11657 9591 11691
rect 9557 11607 9591 11623
rect 9625 11725 9691 11743
rect 9625 11691 9641 11725
rect 9675 11691 9691 11725
rect 9625 11657 9691 11691
rect 9725 11725 9759 11777
rect 9725 11675 9759 11691
rect 9793 11725 9873 11743
rect 9793 11691 9829 11725
rect 9863 11691 9873 11725
rect 9625 11623 9641 11657
rect 9675 11641 9691 11657
rect 9793 11657 9873 11691
rect 9793 11641 9829 11657
rect 9675 11623 9829 11641
rect 9863 11623 9873 11657
rect 9625 11607 9873 11623
rect 9909 11727 9973 11743
rect 9909 11693 9913 11727
rect 9947 11693 9973 11727
rect 9909 11660 9973 11693
rect 9909 11659 9914 11660
rect 9909 11625 9913 11659
rect 9950 11626 9973 11660
rect 9947 11625 9973 11626
rect 9363 11415 9397 11607
rect 9909 11591 9973 11625
rect 9431 11539 9692 11573
rect 9909 11557 9913 11591
rect 9947 11557 9973 11591
rect 9431 11500 9480 11539
rect 9431 11499 9432 11500
rect 9466 11466 9480 11500
rect 9465 11465 9480 11466
rect 9514 11502 9624 11505
rect 9514 11499 9552 11502
rect 9514 11465 9548 11499
rect 9586 11468 9624 11502
rect 9582 11465 9624 11468
rect 9658 11499 9692 11539
rect 9847 11523 9973 11557
rect 9767 11499 9813 11515
rect 9658 11465 9683 11499
rect 9717 11465 9733 11499
rect 9767 11465 9779 11499
rect 9431 11449 9480 11465
rect 9767 11415 9813 11465
rect 9363 11381 9813 11415
rect 9473 11367 9507 11381
rect 9373 11311 9389 11345
rect 9423 11311 9439 11345
rect 9847 11347 9881 11523
rect 9473 11317 9507 11333
rect 9373 11267 9439 11311
rect 9541 11311 9557 11345
rect 9591 11311 9607 11345
rect 9690 11313 9725 11347
rect 9759 11313 9825 11347
rect 9859 11313 9881 11347
rect 9915 11418 9973 11434
rect 9949 11384 9973 11418
rect 9915 11350 9973 11384
rect 9949 11316 9973 11350
rect 9541 11267 9607 11311
rect 9915 11267 9973 11316
rect 9346 11233 9375 11267
rect 9409 11233 9467 11267
rect 9501 11233 9559 11267
rect 9593 11233 9651 11267
rect 9685 11233 9743 11267
rect 9777 11233 9835 11267
rect 9869 11233 9927 11267
rect 9961 11233 9990 11267
rect 9444 11033 9473 11067
rect 9507 11033 9565 11067
rect 9599 11033 9657 11067
rect 9691 11033 9749 11067
rect 9783 11033 9841 11067
rect 9875 11033 9904 11067
rect 9501 10949 9557 11033
rect 9691 10991 9757 11033
rect 9501 10915 9515 10949
rect 9549 10915 9557 10949
rect 9501 10899 9557 10915
rect 9591 10949 9651 10965
rect 9591 10915 9599 10949
rect 9633 10915 9651 10949
rect 9591 10855 9651 10915
rect 9691 10957 9707 10991
rect 9741 10957 9757 10991
rect 9691 10923 9757 10957
rect 9691 10889 9707 10923
rect 9741 10889 9757 10923
rect 9795 10991 9887 10999
rect 9795 10957 9811 10991
rect 9845 10957 9887 10991
rect 9795 10923 9887 10957
rect 9795 10889 9811 10923
rect 9845 10889 9887 10923
rect 9464 10778 9517 10843
rect 9591 10821 9779 10855
rect 9464 10738 9466 10778
rect 9508 10771 9517 10778
rect 9745 10771 9779 10821
rect 9508 10755 9599 10771
rect 9508 10738 9518 10755
rect 9464 10721 9518 10738
rect 9552 10721 9599 10755
rect 9643 10768 9711 10771
rect 9643 10728 9656 10768
rect 9698 10728 9711 10768
rect 9643 10721 9659 10728
rect 9693 10721 9711 10728
rect 9745 10755 9803 10771
rect 9745 10721 9767 10755
rect 9801 10721 9803 10755
rect 9745 10705 9803 10721
rect 9837 10734 9887 10889
rect 9745 10687 9779 10705
rect 9501 10649 9779 10687
rect 9837 10698 9848 10734
rect 9882 10698 9887 10734
rect 9501 10627 9567 10649
rect 9501 10593 9515 10627
rect 9549 10593 9567 10627
rect 9837 10615 9887 10698
rect 9501 10577 9567 10593
rect 9691 10599 9741 10615
rect 9691 10565 9707 10599
rect 9691 10523 9741 10565
rect 9775 10599 9887 10615
rect 9775 10565 9791 10599
rect 9825 10565 9887 10599
rect 9775 10557 9887 10565
rect 9444 10489 9473 10523
rect 9507 10489 9565 10523
rect 9599 10489 9657 10523
rect 9691 10489 9749 10523
rect 9783 10489 9841 10523
rect 9875 10489 9904 10523
rect 6112 6583 6141 6617
rect 6175 6583 6233 6617
rect 6267 6583 6325 6617
rect 6359 6583 6388 6617
rect 6178 6537 6244 6549
rect 6178 6503 6194 6537
rect 6228 6503 6244 6537
rect 6178 6469 6244 6503
rect 6178 6435 6194 6469
rect 6228 6435 6244 6469
rect 6178 6423 6244 6435
rect 6278 6537 6324 6583
rect 6312 6503 6324 6537
rect 6278 6469 6324 6503
rect 6312 6435 6324 6469
rect 6178 6382 6224 6423
rect 6278 6419 6324 6435
rect 6212 6348 6224 6382
rect 6178 6303 6224 6348
rect 6258 6350 6274 6385
rect 6308 6350 6324 6385
rect 6258 6337 6324 6350
rect 6178 6285 6244 6303
rect 6178 6251 6194 6285
rect 6228 6251 6244 6285
rect 6178 6217 6244 6251
rect 6178 6183 6194 6217
rect 6228 6183 6244 6217
rect 6178 6149 6244 6183
rect 6178 6115 6194 6149
rect 6228 6115 6244 6149
rect 6178 6107 6244 6115
rect 6278 6285 6320 6301
rect 6312 6251 6320 6285
rect 6278 6217 6320 6251
rect 6312 6183 6320 6217
rect 6278 6149 6320 6183
rect 6312 6115 6320 6149
rect 6278 6073 6320 6115
rect 6112 6039 6141 6073
rect 6175 6039 6233 6073
rect 6267 6039 6325 6073
rect 6359 6039 6388 6073
rect 10018 5951 10047 5985
rect 10081 5951 10139 5985
rect 10173 5951 10231 5985
rect 10265 5951 10323 5985
rect 10357 5951 10415 5985
rect 10449 5951 10507 5985
rect 10541 5951 10599 5985
rect 10633 5951 10691 5985
rect 10725 5951 10783 5985
rect 10817 5951 10875 5985
rect 10909 5951 10967 5985
rect 11001 5951 11059 5985
rect 11093 5951 11151 5985
rect 11185 5951 11243 5985
rect 11277 5951 11335 5985
rect 11369 5951 11427 5985
rect 11461 5951 11490 5985
rect 10042 5873 10122 5917
rect 10171 5913 10237 5951
rect 10171 5879 10187 5913
rect 10221 5879 10237 5913
rect 10271 5901 10473 5917
rect 10042 5839 10088 5873
rect 10271 5867 10439 5901
rect 10271 5845 10305 5867
rect 10439 5849 10473 5867
rect 10540 5896 10574 5917
rect 10608 5913 10674 5951
rect 10608 5879 10624 5913
rect 10658 5879 10674 5913
rect 10708 5896 10742 5917
rect 10042 5806 10122 5839
rect 10157 5811 10305 5845
rect 10540 5845 10574 5862
rect 10776 5904 10842 5951
rect 10776 5870 10792 5904
rect 10826 5870 10842 5904
rect 10896 5896 10930 5917
rect 10708 5845 10742 5862
rect 10042 5671 10108 5806
rect 10157 5769 10191 5811
rect 10142 5753 10191 5769
rect 10398 5781 10410 5815
rect 10444 5781 10497 5815
rect 10540 5811 10742 5845
rect 10964 5913 11030 5951
rect 10964 5879 10980 5913
rect 11014 5879 11030 5913
rect 11064 5896 11098 5917
rect 10896 5845 10930 5862
rect 11064 5845 11098 5862
rect 10896 5811 11098 5845
rect 11148 5896 11268 5917
rect 11182 5862 11268 5896
rect 11321 5909 11387 5951
rect 12080 5939 12109 5973
rect 12143 5939 12201 5973
rect 12235 5939 12293 5973
rect 12327 5939 12385 5973
rect 12419 5939 12477 5973
rect 12511 5939 12569 5973
rect 12603 5939 12661 5973
rect 12695 5939 12753 5973
rect 12787 5939 12845 5973
rect 12879 5939 12937 5973
rect 12971 5939 13029 5973
rect 13063 5939 13121 5973
rect 13155 5939 13213 5973
rect 13247 5939 13305 5973
rect 13339 5939 13397 5973
rect 13431 5939 13489 5973
rect 13523 5939 13552 5973
rect 14038 5947 14067 5981
rect 14101 5947 14159 5981
rect 14193 5947 14251 5981
rect 14285 5947 14343 5981
rect 14377 5947 14435 5981
rect 14469 5947 14527 5981
rect 14561 5947 14619 5981
rect 14653 5947 14711 5981
rect 14745 5947 14803 5981
rect 14837 5947 14895 5981
rect 14929 5947 14987 5981
rect 15021 5947 15079 5981
rect 15113 5947 15171 5981
rect 15205 5947 15263 5981
rect 15297 5947 15355 5981
rect 15389 5947 15447 5981
rect 15481 5947 15510 5981
rect 16032 5953 16061 5987
rect 16095 5953 16153 5987
rect 16187 5953 16245 5987
rect 16279 5953 16337 5987
rect 16371 5953 16429 5987
rect 16463 5953 16521 5987
rect 16555 5953 16613 5987
rect 16647 5953 16705 5987
rect 16739 5953 16797 5987
rect 16831 5953 16889 5987
rect 16923 5953 16981 5987
rect 17015 5953 17073 5987
rect 17107 5953 17165 5987
rect 17199 5953 17257 5987
rect 17291 5953 17349 5987
rect 17383 5953 17441 5987
rect 17475 5953 17504 5987
rect 11321 5875 11337 5909
rect 11371 5875 11387 5909
rect 11148 5841 11268 5862
rect 11421 5873 11473 5917
rect 11148 5815 11387 5841
rect 11148 5781 11150 5815
rect 11184 5807 11387 5815
rect 11184 5781 11196 5807
rect 10398 5777 10497 5781
rect 10176 5719 10191 5753
rect 10142 5703 10191 5719
rect 10225 5747 10241 5761
rect 10225 5713 10226 5747
rect 10275 5727 10313 5761
rect 10398 5743 10481 5777
rect 10515 5743 10531 5777
rect 10565 5743 10581 5777
rect 10615 5747 10640 5777
rect 10260 5713 10313 5727
rect 10565 5713 10594 5743
rect 10628 5713 10640 5747
rect 10699 5718 10932 5775
rect 11353 5769 11387 5807
rect 11455 5839 11473 5873
rect 11421 5802 11473 5839
rect 10042 5633 10122 5671
rect 10042 5599 10088 5633
rect 1836 5531 1865 5565
rect 1899 5531 1957 5565
rect 1991 5531 2049 5565
rect 2083 5531 2141 5565
rect 2175 5531 2233 5565
rect 2267 5531 2325 5565
rect 2359 5531 2417 5565
rect 2451 5531 2509 5565
rect 2543 5531 2601 5565
rect 2635 5531 2693 5565
rect 2727 5531 2785 5565
rect 2819 5531 2877 5565
rect 2911 5531 2969 5565
rect 3003 5531 3061 5565
rect 3095 5531 3153 5565
rect 3187 5531 3245 5565
rect 3279 5531 3308 5565
rect 1860 5453 1940 5497
rect 1989 5493 2055 5531
rect 1989 5459 2005 5493
rect 2039 5459 2055 5493
rect 2089 5481 2291 5497
rect 1860 5419 1906 5453
rect 2089 5447 2257 5481
rect 2089 5425 2123 5447
rect 2257 5429 2291 5447
rect 2358 5476 2392 5497
rect 2426 5493 2492 5531
rect 2426 5459 2442 5493
rect 2476 5459 2492 5493
rect 2526 5476 2560 5497
rect 1860 5386 1940 5419
rect 1975 5391 2123 5425
rect 2358 5425 2392 5442
rect 2594 5484 2660 5531
rect 2594 5450 2610 5484
rect 2644 5450 2660 5484
rect 2714 5476 2748 5497
rect 2526 5425 2560 5442
rect 1860 5251 1926 5386
rect 1975 5349 2009 5391
rect 1960 5333 2009 5349
rect 2216 5361 2228 5395
rect 2262 5361 2315 5395
rect 2358 5391 2560 5425
rect 2782 5493 2848 5531
rect 2782 5459 2798 5493
rect 2832 5459 2848 5493
rect 2882 5476 2916 5497
rect 2714 5425 2748 5442
rect 2882 5425 2916 5442
rect 2714 5391 2916 5425
rect 2966 5476 3086 5497
rect 3000 5442 3086 5476
rect 3139 5489 3205 5531
rect 3970 5523 3999 5557
rect 4033 5523 4091 5557
rect 4125 5523 4183 5557
rect 4217 5523 4275 5557
rect 4309 5523 4367 5557
rect 4401 5523 4459 5557
rect 4493 5523 4551 5557
rect 4585 5523 4643 5557
rect 4677 5523 4735 5557
rect 4769 5523 4827 5557
rect 4861 5523 4919 5557
rect 4953 5523 5011 5557
rect 5045 5523 5103 5557
rect 5137 5523 5195 5557
rect 5229 5523 5287 5557
rect 5321 5523 5379 5557
rect 5413 5523 5442 5557
rect 5922 5523 5951 5557
rect 5985 5523 6043 5557
rect 6077 5523 6135 5557
rect 6169 5523 6227 5557
rect 6261 5523 6319 5557
rect 6353 5523 6411 5557
rect 6445 5523 6503 5557
rect 6537 5523 6595 5557
rect 6629 5523 6687 5557
rect 6721 5523 6779 5557
rect 6813 5523 6871 5557
rect 6905 5523 6963 5557
rect 6997 5523 7055 5557
rect 7089 5523 7147 5557
rect 7181 5523 7239 5557
rect 7273 5523 7331 5557
rect 7365 5523 7394 5557
rect 7924 5529 7953 5563
rect 7987 5529 8045 5563
rect 8079 5529 8137 5563
rect 8171 5529 8229 5563
rect 8263 5529 8321 5563
rect 8355 5529 8413 5563
rect 8447 5529 8505 5563
rect 8539 5529 8597 5563
rect 8631 5529 8689 5563
rect 8723 5529 8781 5563
rect 8815 5529 8873 5563
rect 8907 5529 8965 5563
rect 8999 5529 9057 5563
rect 9091 5529 9149 5563
rect 9183 5529 9241 5563
rect 9275 5529 9333 5563
rect 9367 5529 9396 5563
rect 10042 5543 10122 5599
rect 10157 5581 10191 5703
rect 10279 5649 10318 5679
rect 10279 5615 10313 5649
rect 10352 5645 10363 5679
rect 10699 5665 10733 5718
rect 10347 5615 10363 5645
rect 10409 5649 10666 5665
rect 10443 5631 10666 5649
rect 10700 5631 10733 5665
rect 10778 5679 10850 5681
rect 10812 5665 10850 5679
rect 10778 5631 10783 5645
rect 10817 5631 10850 5665
rect 10443 5615 10459 5631
rect 10778 5615 10850 5631
rect 10898 5649 10932 5718
rect 10966 5747 11044 5762
rect 11242 5753 11308 5769
rect 11242 5747 11274 5753
rect 11000 5746 11044 5747
rect 11000 5713 11010 5746
rect 10966 5712 11010 5713
rect 10966 5696 11044 5712
rect 11082 5713 11106 5747
rect 11140 5713 11156 5747
rect 11276 5713 11308 5719
rect 11082 5649 11116 5713
rect 11274 5703 11308 5713
rect 11353 5753 11404 5769
rect 11353 5719 11370 5753
rect 11353 5703 11404 5719
rect 10898 5615 11116 5649
rect 11184 5645 11230 5679
rect 11150 5642 11230 5645
rect 11353 5643 11387 5703
rect 11438 5671 11473 5802
rect 10409 5614 10459 5615
rect 10157 5547 10290 5581
rect 10409 5580 10418 5614
rect 10452 5580 10459 5614
rect 11150 5608 11196 5642
rect 11150 5592 11230 5608
rect 10409 5577 10459 5580
rect 3139 5455 3155 5489
rect 3189 5455 3205 5489
rect 2966 5421 3086 5442
rect 3239 5453 3291 5497
rect 2966 5395 3205 5421
rect 2966 5361 2968 5395
rect 3002 5387 3205 5395
rect 3002 5361 3014 5387
rect 2216 5357 2315 5361
rect 1994 5299 2009 5333
rect 1960 5283 2009 5299
rect 2043 5327 2059 5341
rect 2043 5293 2044 5327
rect 2093 5307 2131 5341
rect 2216 5323 2299 5357
rect 2333 5323 2349 5357
rect 2383 5323 2399 5357
rect 2433 5327 2458 5357
rect 2078 5293 2131 5307
rect 2383 5293 2412 5323
rect 2446 5293 2458 5327
rect 2517 5298 2750 5355
rect 3171 5349 3205 5387
rect 3273 5419 3291 5453
rect 3239 5382 3291 5419
rect 1860 5213 1940 5251
rect 1860 5179 1906 5213
rect 1860 5123 1940 5179
rect 1975 5161 2009 5283
rect 2097 5229 2136 5259
rect 2097 5195 2131 5229
rect 2170 5225 2181 5259
rect 2517 5245 2551 5298
rect 2165 5195 2181 5225
rect 2227 5229 2484 5245
rect 2261 5211 2484 5229
rect 2518 5211 2551 5245
rect 2596 5259 2668 5261
rect 2630 5245 2668 5259
rect 2596 5211 2601 5225
rect 2635 5211 2668 5245
rect 2261 5195 2277 5211
rect 2596 5195 2668 5211
rect 2716 5229 2750 5298
rect 2784 5327 2862 5342
rect 3060 5333 3126 5349
rect 3060 5327 3092 5333
rect 2818 5326 2862 5327
rect 2818 5293 2828 5326
rect 2784 5292 2828 5293
rect 2784 5276 2862 5292
rect 2900 5293 2924 5327
rect 2958 5293 2974 5327
rect 3094 5293 3126 5299
rect 2900 5229 2934 5293
rect 3092 5283 3126 5293
rect 3171 5333 3222 5349
rect 3171 5299 3188 5333
rect 3171 5283 3222 5299
rect 2716 5195 2934 5229
rect 3002 5225 3048 5259
rect 2968 5222 3048 5225
rect 3171 5223 3205 5283
rect 3256 5251 3291 5382
rect 2227 5194 2277 5195
rect 1975 5127 2108 5161
rect 2227 5160 2236 5194
rect 2270 5160 2277 5194
rect 2968 5188 3014 5222
rect 2968 5172 3048 5188
rect 2227 5157 2277 5160
rect 1860 5089 1906 5123
rect 2074 5123 2108 5127
rect 2358 5127 2560 5161
rect 2074 5105 2291 5123
rect 1860 5055 1940 5089
rect 1974 5059 1990 5093
rect 2024 5059 2040 5093
rect 1974 5021 2040 5059
rect 2074 5071 2257 5105
rect 2074 5055 2291 5071
rect 2358 5110 2392 5127
rect 2526 5110 2560 5127
rect 2358 5055 2392 5076
rect 2426 5059 2442 5093
rect 2476 5059 2492 5093
rect 2426 5021 2492 5059
rect 2701 5127 2916 5161
rect 3087 5159 3205 5223
rect 3239 5210 3291 5251
rect 3273 5186 3291 5210
rect 3087 5135 3121 5159
rect 2701 5110 2748 5127
rect 2526 5055 2560 5076
rect 2594 5063 2610 5097
rect 2644 5063 2660 5097
rect 2594 5021 2660 5063
rect 2701 5076 2714 5110
rect 2882 5110 2916 5127
rect 2701 5055 2748 5076
rect 2782 5059 2798 5093
rect 2832 5059 2848 5093
rect 2782 5021 2848 5059
rect 2882 5055 2916 5076
rect 2966 5110 3121 5135
rect 3239 5150 3244 5176
rect 3284 5150 3291 5186
rect 3000 5076 3121 5110
rect 2966 5055 3121 5076
rect 3155 5101 3205 5118
rect 3189 5067 3205 5101
rect 3155 5021 3205 5067
rect 3239 5116 3291 5150
rect 3273 5082 3291 5116
rect 3239 5055 3291 5082
rect 3994 5445 4074 5489
rect 4123 5485 4189 5523
rect 4123 5451 4139 5485
rect 4173 5451 4189 5485
rect 4223 5473 4425 5489
rect 3994 5411 4040 5445
rect 4223 5439 4391 5473
rect 4223 5417 4257 5439
rect 4391 5421 4425 5439
rect 4492 5468 4526 5489
rect 4560 5485 4626 5523
rect 4560 5451 4576 5485
rect 4610 5451 4626 5485
rect 4660 5468 4694 5489
rect 3994 5378 4074 5411
rect 4109 5383 4257 5417
rect 4492 5417 4526 5434
rect 4728 5476 4794 5523
rect 4728 5442 4744 5476
rect 4778 5442 4794 5476
rect 4848 5468 4882 5489
rect 4660 5417 4694 5434
rect 3994 5243 4060 5378
rect 4109 5341 4143 5383
rect 4094 5325 4143 5341
rect 4350 5353 4362 5387
rect 4396 5353 4449 5387
rect 4492 5383 4694 5417
rect 4916 5485 4982 5523
rect 4916 5451 4932 5485
rect 4966 5451 4982 5485
rect 5016 5468 5050 5489
rect 4848 5417 4882 5434
rect 5016 5417 5050 5434
rect 4848 5383 5050 5417
rect 5100 5468 5220 5489
rect 5134 5434 5220 5468
rect 5273 5481 5339 5523
rect 5273 5447 5289 5481
rect 5323 5447 5339 5481
rect 5100 5413 5220 5434
rect 5373 5445 5425 5489
rect 5100 5387 5339 5413
rect 5100 5353 5102 5387
rect 5136 5379 5339 5387
rect 5136 5353 5148 5379
rect 4350 5349 4449 5353
rect 4128 5291 4143 5325
rect 4094 5275 4143 5291
rect 4177 5319 4193 5333
rect 4177 5285 4178 5319
rect 4227 5299 4265 5333
rect 4350 5315 4433 5349
rect 4467 5315 4483 5349
rect 4517 5315 4533 5349
rect 4567 5319 4592 5349
rect 4212 5285 4265 5299
rect 4517 5285 4546 5315
rect 4580 5285 4592 5319
rect 4651 5290 4884 5347
rect 5305 5341 5339 5379
rect 5407 5411 5425 5445
rect 5373 5374 5425 5411
rect 3994 5205 4074 5243
rect 3994 5171 4040 5205
rect 3994 5115 4074 5171
rect 4109 5153 4143 5275
rect 4231 5221 4270 5251
rect 4231 5187 4265 5221
rect 4304 5217 4315 5251
rect 4651 5237 4685 5290
rect 4299 5187 4315 5217
rect 4361 5221 4618 5237
rect 4395 5203 4618 5221
rect 4652 5203 4685 5237
rect 4730 5251 4802 5253
rect 4764 5237 4802 5251
rect 4730 5203 4735 5217
rect 4769 5203 4802 5237
rect 4395 5187 4411 5203
rect 4730 5187 4802 5203
rect 4850 5221 4884 5290
rect 4918 5319 4996 5334
rect 5194 5325 5260 5341
rect 5194 5319 5226 5325
rect 4952 5318 4996 5319
rect 4952 5285 4962 5318
rect 4918 5284 4962 5285
rect 4918 5268 4996 5284
rect 5034 5285 5058 5319
rect 5092 5285 5108 5319
rect 5228 5285 5260 5291
rect 5034 5221 5068 5285
rect 5226 5275 5260 5285
rect 5305 5325 5356 5341
rect 5305 5291 5322 5325
rect 5305 5275 5356 5291
rect 4850 5187 5068 5221
rect 5136 5217 5182 5251
rect 5102 5214 5182 5217
rect 5305 5215 5339 5275
rect 5390 5243 5425 5374
rect 4361 5184 4411 5187
rect 4109 5119 4242 5153
rect 4361 5150 4368 5184
rect 4402 5150 4411 5184
rect 5102 5180 5148 5214
rect 5102 5164 5182 5180
rect 4361 5149 4411 5150
rect 3994 5081 4040 5115
rect 4208 5115 4242 5119
rect 4492 5119 4694 5153
rect 4208 5097 4425 5115
rect 3994 5047 4074 5081
rect 4108 5051 4124 5085
rect 4158 5051 4174 5085
rect 1836 4987 1865 5021
rect 1899 4987 1957 5021
rect 1991 4987 2049 5021
rect 2083 4987 2141 5021
rect 2175 4987 2233 5021
rect 2267 4987 2325 5021
rect 2359 4987 2417 5021
rect 2451 4987 2509 5021
rect 2543 4987 2601 5021
rect 2635 4987 2693 5021
rect 2727 4987 2785 5021
rect 2819 4987 2877 5021
rect 2911 4987 2969 5021
rect 3003 4987 3061 5021
rect 3095 4987 3153 5021
rect 3187 4987 3245 5021
rect 3279 4987 3308 5021
rect 4108 5013 4174 5051
rect 4208 5063 4391 5097
rect 4208 5047 4425 5063
rect 4492 5102 4526 5119
rect 4660 5102 4694 5119
rect 4492 5047 4526 5068
rect 4560 5051 4576 5085
rect 4610 5051 4626 5085
rect 4560 5013 4626 5051
rect 4835 5119 5050 5153
rect 5221 5151 5339 5215
rect 5373 5202 5425 5243
rect 5407 5178 5425 5202
rect 5221 5127 5255 5151
rect 4835 5102 4882 5119
rect 4660 5047 4694 5068
rect 4728 5055 4744 5089
rect 4778 5055 4794 5089
rect 4728 5013 4794 5055
rect 4835 5068 4848 5102
rect 5016 5102 5050 5119
rect 4835 5047 4882 5068
rect 4916 5051 4932 5085
rect 4966 5051 4982 5085
rect 4916 5013 4982 5051
rect 5016 5047 5050 5068
rect 5100 5102 5255 5127
rect 5373 5142 5384 5168
rect 5418 5142 5425 5178
rect 5134 5068 5255 5102
rect 5100 5047 5255 5068
rect 5289 5093 5339 5110
rect 5323 5059 5339 5093
rect 5289 5013 5339 5059
rect 5373 5108 5425 5142
rect 5407 5074 5425 5108
rect 5373 5047 5425 5074
rect 5946 5445 6026 5489
rect 6075 5485 6141 5523
rect 6075 5451 6091 5485
rect 6125 5451 6141 5485
rect 6175 5473 6377 5489
rect 5946 5411 5992 5445
rect 6175 5439 6343 5473
rect 6175 5417 6209 5439
rect 6343 5421 6377 5439
rect 6444 5468 6478 5489
rect 6512 5485 6578 5523
rect 6512 5451 6528 5485
rect 6562 5451 6578 5485
rect 6612 5468 6646 5489
rect 5946 5378 6026 5411
rect 6061 5383 6209 5417
rect 6444 5417 6478 5434
rect 6680 5476 6746 5523
rect 6680 5442 6696 5476
rect 6730 5442 6746 5476
rect 6800 5468 6834 5489
rect 6612 5417 6646 5434
rect 5946 5243 6012 5378
rect 6061 5341 6095 5383
rect 6046 5325 6095 5341
rect 6302 5353 6314 5387
rect 6348 5353 6401 5387
rect 6444 5383 6646 5417
rect 6868 5485 6934 5523
rect 6868 5451 6884 5485
rect 6918 5451 6934 5485
rect 6968 5468 7002 5489
rect 6800 5417 6834 5434
rect 6968 5417 7002 5434
rect 6800 5383 7002 5417
rect 7052 5468 7172 5489
rect 7086 5434 7172 5468
rect 7225 5481 7291 5523
rect 7225 5447 7241 5481
rect 7275 5447 7291 5481
rect 7052 5413 7172 5434
rect 7325 5445 7377 5489
rect 7052 5387 7291 5413
rect 7052 5353 7054 5387
rect 7088 5379 7291 5387
rect 7088 5353 7100 5379
rect 6302 5349 6401 5353
rect 6080 5291 6095 5325
rect 6046 5275 6095 5291
rect 6129 5319 6145 5333
rect 6129 5285 6130 5319
rect 6179 5299 6217 5333
rect 6302 5315 6385 5349
rect 6419 5315 6435 5349
rect 6469 5315 6485 5349
rect 6519 5319 6544 5349
rect 6164 5285 6217 5299
rect 6469 5285 6498 5315
rect 6532 5285 6544 5319
rect 6603 5290 6836 5347
rect 7257 5341 7291 5379
rect 7359 5411 7377 5445
rect 7325 5374 7377 5411
rect 5946 5205 6026 5243
rect 5946 5171 5992 5205
rect 5946 5115 6026 5171
rect 6061 5153 6095 5275
rect 6183 5221 6222 5251
rect 6183 5187 6217 5221
rect 6256 5217 6267 5251
rect 6603 5237 6637 5290
rect 6251 5187 6267 5217
rect 6313 5221 6570 5237
rect 6347 5203 6570 5221
rect 6604 5203 6637 5237
rect 6682 5251 6754 5253
rect 6716 5237 6754 5251
rect 6682 5203 6687 5217
rect 6721 5203 6754 5237
rect 6347 5187 6363 5203
rect 6682 5187 6754 5203
rect 6802 5221 6836 5290
rect 6870 5319 6948 5334
rect 7146 5325 7212 5341
rect 7146 5319 7178 5325
rect 6904 5318 6948 5319
rect 6904 5285 6914 5318
rect 6870 5284 6914 5285
rect 6870 5268 6948 5284
rect 6986 5285 7010 5319
rect 7044 5285 7060 5319
rect 7180 5285 7212 5291
rect 6986 5221 7020 5285
rect 7178 5275 7212 5285
rect 7257 5325 7308 5341
rect 7257 5291 7274 5325
rect 7257 5275 7308 5291
rect 6802 5187 7020 5221
rect 7088 5217 7134 5251
rect 7054 5214 7134 5217
rect 7257 5215 7291 5275
rect 7342 5243 7377 5374
rect 6313 5184 6363 5187
rect 6061 5119 6194 5153
rect 6313 5150 6320 5184
rect 6354 5150 6363 5184
rect 7054 5180 7100 5214
rect 7054 5164 7134 5180
rect 6313 5149 6363 5150
rect 5946 5081 5992 5115
rect 6160 5115 6194 5119
rect 6444 5119 6646 5153
rect 6160 5097 6377 5115
rect 5946 5047 6026 5081
rect 6060 5051 6076 5085
rect 6110 5051 6126 5085
rect 6060 5013 6126 5051
rect 6160 5063 6343 5097
rect 6160 5047 6377 5063
rect 6444 5102 6478 5119
rect 6612 5102 6646 5119
rect 6444 5047 6478 5068
rect 6512 5051 6528 5085
rect 6562 5051 6578 5085
rect 6512 5013 6578 5051
rect 6787 5119 7002 5153
rect 7173 5151 7291 5215
rect 7325 5202 7377 5243
rect 7359 5178 7377 5202
rect 7173 5127 7207 5151
rect 6787 5102 6834 5119
rect 6612 5047 6646 5068
rect 6680 5055 6696 5089
rect 6730 5055 6746 5089
rect 6680 5013 6746 5055
rect 6787 5068 6800 5102
rect 6968 5102 7002 5119
rect 6787 5047 6834 5068
rect 6868 5051 6884 5085
rect 6918 5051 6934 5085
rect 6868 5013 6934 5051
rect 6968 5047 7002 5068
rect 7052 5102 7207 5127
rect 7325 5142 7336 5168
rect 7370 5142 7377 5178
rect 7086 5068 7207 5102
rect 7052 5047 7207 5068
rect 7241 5093 7291 5110
rect 7275 5059 7291 5093
rect 7241 5013 7291 5059
rect 7325 5108 7377 5142
rect 7359 5074 7377 5108
rect 7325 5047 7377 5074
rect 7948 5451 8028 5495
rect 8077 5491 8143 5529
rect 8077 5457 8093 5491
rect 8127 5457 8143 5491
rect 8177 5479 8379 5495
rect 7948 5417 7994 5451
rect 8177 5445 8345 5479
rect 8177 5423 8211 5445
rect 8345 5427 8379 5445
rect 8446 5474 8480 5495
rect 8514 5491 8580 5529
rect 8514 5457 8530 5491
rect 8564 5457 8580 5491
rect 8614 5474 8648 5495
rect 7948 5384 8028 5417
rect 8063 5389 8211 5423
rect 8446 5423 8480 5440
rect 8682 5482 8748 5529
rect 8682 5448 8698 5482
rect 8732 5448 8748 5482
rect 8802 5474 8836 5495
rect 8614 5423 8648 5440
rect 7948 5249 8014 5384
rect 8063 5347 8097 5389
rect 8048 5331 8097 5347
rect 8304 5359 8316 5393
rect 8350 5359 8403 5393
rect 8446 5389 8648 5423
rect 8870 5491 8936 5529
rect 8870 5457 8886 5491
rect 8920 5457 8936 5491
rect 8970 5474 9004 5495
rect 8802 5423 8836 5440
rect 8970 5423 9004 5440
rect 8802 5389 9004 5423
rect 9054 5474 9174 5495
rect 9088 5440 9174 5474
rect 9227 5487 9293 5529
rect 10042 5509 10088 5543
rect 10256 5543 10290 5547
rect 10540 5547 10742 5581
rect 10256 5525 10473 5543
rect 9227 5453 9243 5487
rect 9277 5453 9293 5487
rect 9054 5419 9174 5440
rect 9327 5451 9379 5495
rect 10042 5475 10122 5509
rect 10156 5479 10172 5513
rect 10206 5479 10222 5513
rect 9054 5393 9293 5419
rect 9054 5359 9056 5393
rect 9090 5385 9293 5393
rect 9090 5359 9102 5385
rect 8304 5355 8403 5359
rect 8082 5297 8097 5331
rect 8048 5281 8097 5297
rect 8131 5325 8147 5339
rect 8131 5291 8132 5325
rect 8181 5305 8219 5339
rect 8304 5321 8387 5355
rect 8421 5321 8437 5355
rect 8471 5321 8487 5355
rect 8521 5325 8546 5355
rect 8166 5291 8219 5305
rect 8471 5291 8500 5321
rect 8534 5291 8546 5325
rect 8605 5296 8838 5353
rect 9259 5347 9293 5385
rect 9361 5417 9379 5451
rect 10156 5441 10222 5479
rect 10256 5491 10439 5525
rect 10256 5475 10473 5491
rect 10540 5530 10574 5547
rect 10708 5530 10742 5547
rect 10540 5475 10574 5496
rect 10608 5479 10624 5513
rect 10658 5479 10674 5513
rect 10608 5441 10674 5479
rect 10883 5547 11098 5581
rect 11269 5579 11387 5643
rect 11421 5630 11473 5671
rect 11455 5606 11473 5630
rect 11269 5555 11303 5579
rect 10883 5530 10930 5547
rect 10708 5475 10742 5496
rect 10776 5483 10792 5517
rect 10826 5483 10842 5517
rect 10776 5441 10842 5483
rect 10883 5496 10896 5530
rect 11064 5530 11098 5547
rect 10883 5475 10930 5496
rect 10964 5479 10980 5513
rect 11014 5479 11030 5513
rect 10964 5441 11030 5479
rect 11064 5475 11098 5496
rect 11148 5530 11303 5555
rect 11421 5570 11426 5596
rect 11466 5570 11473 5606
rect 11182 5496 11303 5530
rect 11148 5475 11303 5496
rect 11337 5521 11387 5538
rect 11371 5487 11387 5521
rect 11337 5441 11387 5487
rect 11421 5536 11473 5570
rect 11455 5502 11473 5536
rect 11421 5475 11473 5502
rect 12104 5861 12184 5905
rect 12233 5901 12299 5939
rect 12233 5867 12249 5901
rect 12283 5867 12299 5901
rect 12333 5889 12535 5905
rect 12104 5827 12150 5861
rect 12333 5855 12501 5889
rect 12333 5833 12367 5855
rect 12501 5837 12535 5855
rect 12602 5884 12636 5905
rect 12670 5901 12736 5939
rect 12670 5867 12686 5901
rect 12720 5867 12736 5901
rect 12770 5884 12804 5905
rect 12104 5794 12184 5827
rect 12219 5799 12367 5833
rect 12602 5833 12636 5850
rect 12838 5892 12904 5939
rect 12838 5858 12854 5892
rect 12888 5858 12904 5892
rect 12958 5884 12992 5905
rect 12770 5833 12804 5850
rect 12104 5659 12170 5794
rect 12219 5757 12253 5799
rect 12204 5741 12253 5757
rect 12460 5769 12472 5803
rect 12506 5769 12559 5803
rect 12602 5799 12804 5833
rect 13026 5901 13092 5939
rect 13026 5867 13042 5901
rect 13076 5867 13092 5901
rect 13126 5884 13160 5905
rect 12958 5833 12992 5850
rect 13126 5833 13160 5850
rect 12958 5799 13160 5833
rect 13210 5884 13330 5905
rect 13244 5850 13330 5884
rect 13383 5897 13449 5939
rect 13383 5863 13399 5897
rect 13433 5863 13449 5897
rect 13210 5829 13330 5850
rect 13483 5861 13535 5905
rect 13210 5803 13449 5829
rect 13210 5769 13212 5803
rect 13246 5795 13449 5803
rect 13246 5769 13258 5795
rect 12460 5765 12559 5769
rect 12238 5707 12253 5741
rect 12204 5691 12253 5707
rect 12287 5735 12303 5749
rect 12287 5701 12288 5735
rect 12337 5715 12375 5749
rect 12460 5731 12543 5765
rect 12577 5731 12593 5765
rect 12627 5731 12643 5765
rect 12677 5735 12702 5765
rect 12322 5701 12375 5715
rect 12627 5701 12656 5731
rect 12690 5701 12702 5735
rect 12761 5706 12994 5763
rect 13415 5757 13449 5795
rect 13517 5827 13535 5861
rect 13483 5790 13535 5827
rect 12104 5621 12184 5659
rect 12104 5587 12150 5621
rect 12104 5531 12184 5587
rect 12219 5569 12253 5691
rect 12341 5637 12380 5667
rect 12341 5603 12375 5637
rect 12414 5633 12425 5667
rect 12761 5653 12795 5706
rect 12409 5603 12425 5633
rect 12471 5637 12728 5653
rect 12505 5619 12728 5637
rect 12762 5619 12795 5653
rect 12840 5667 12912 5669
rect 12874 5653 12912 5667
rect 12840 5619 12845 5633
rect 12879 5619 12912 5653
rect 12505 5603 12521 5619
rect 12840 5603 12912 5619
rect 12960 5637 12994 5706
rect 13028 5735 13106 5750
rect 13304 5741 13370 5757
rect 13304 5735 13336 5741
rect 13062 5734 13106 5735
rect 13062 5701 13072 5734
rect 13028 5700 13072 5701
rect 13028 5684 13106 5700
rect 13144 5701 13168 5735
rect 13202 5701 13218 5735
rect 13338 5701 13370 5707
rect 13144 5637 13178 5701
rect 13336 5691 13370 5701
rect 13415 5741 13466 5757
rect 13415 5707 13432 5741
rect 13415 5691 13466 5707
rect 12960 5603 13178 5637
rect 13246 5633 13292 5667
rect 13212 5630 13292 5633
rect 13415 5631 13449 5691
rect 13500 5659 13535 5790
rect 12471 5600 12521 5603
rect 12219 5535 12352 5569
rect 12471 5566 12478 5600
rect 12512 5566 12521 5600
rect 13212 5596 13258 5630
rect 13212 5580 13292 5596
rect 12471 5565 12521 5566
rect 12104 5497 12150 5531
rect 12318 5531 12352 5535
rect 12602 5535 12804 5569
rect 12318 5513 12535 5531
rect 12104 5463 12184 5497
rect 12218 5467 12234 5501
rect 12268 5467 12284 5501
rect 9327 5380 9379 5417
rect 10018 5407 10047 5441
rect 10081 5407 10139 5441
rect 10173 5407 10231 5441
rect 10265 5407 10323 5441
rect 10357 5407 10415 5441
rect 10449 5407 10507 5441
rect 10541 5407 10599 5441
rect 10633 5407 10691 5441
rect 10725 5407 10783 5441
rect 10817 5407 10875 5441
rect 10909 5407 10967 5441
rect 11001 5407 11059 5441
rect 11093 5407 11151 5441
rect 11185 5407 11243 5441
rect 11277 5407 11335 5441
rect 11369 5407 11427 5441
rect 11461 5407 11490 5441
rect 12218 5429 12284 5467
rect 12318 5479 12501 5513
rect 12318 5463 12535 5479
rect 12602 5518 12636 5535
rect 12770 5518 12804 5535
rect 12602 5463 12636 5484
rect 12670 5467 12686 5501
rect 12720 5467 12736 5501
rect 12670 5429 12736 5467
rect 12945 5535 13160 5569
rect 13331 5567 13449 5631
rect 13483 5618 13535 5659
rect 13517 5594 13535 5618
rect 13331 5543 13365 5567
rect 12945 5518 12992 5535
rect 12770 5463 12804 5484
rect 12838 5471 12854 5505
rect 12888 5471 12904 5505
rect 12838 5429 12904 5471
rect 12945 5484 12958 5518
rect 13126 5518 13160 5535
rect 12945 5463 12992 5484
rect 13026 5467 13042 5501
rect 13076 5467 13092 5501
rect 13026 5429 13092 5467
rect 13126 5463 13160 5484
rect 13210 5518 13365 5543
rect 13483 5558 13494 5584
rect 13528 5558 13535 5594
rect 13244 5484 13365 5518
rect 13210 5463 13365 5484
rect 13399 5509 13449 5526
rect 13433 5475 13449 5509
rect 13399 5429 13449 5475
rect 13483 5524 13535 5558
rect 13517 5490 13535 5524
rect 13483 5463 13535 5490
rect 14062 5869 14142 5913
rect 14191 5909 14257 5947
rect 14191 5875 14207 5909
rect 14241 5875 14257 5909
rect 14291 5897 14493 5913
rect 14062 5835 14108 5869
rect 14291 5863 14459 5897
rect 14291 5841 14325 5863
rect 14459 5845 14493 5863
rect 14560 5892 14594 5913
rect 14628 5909 14694 5947
rect 14628 5875 14644 5909
rect 14678 5875 14694 5909
rect 14728 5892 14762 5913
rect 14062 5802 14142 5835
rect 14177 5807 14325 5841
rect 14560 5841 14594 5858
rect 14796 5900 14862 5947
rect 14796 5866 14812 5900
rect 14846 5866 14862 5900
rect 14916 5892 14950 5913
rect 14728 5841 14762 5858
rect 14062 5667 14128 5802
rect 14177 5765 14211 5807
rect 14162 5749 14211 5765
rect 14418 5777 14430 5811
rect 14464 5777 14517 5811
rect 14560 5807 14762 5841
rect 14984 5909 15050 5947
rect 14984 5875 15000 5909
rect 15034 5875 15050 5909
rect 15084 5892 15118 5913
rect 14916 5841 14950 5858
rect 15084 5841 15118 5858
rect 14916 5807 15118 5841
rect 15168 5892 15288 5913
rect 15202 5858 15288 5892
rect 15341 5905 15407 5947
rect 15341 5871 15357 5905
rect 15391 5871 15407 5905
rect 15168 5837 15288 5858
rect 15441 5869 15493 5913
rect 15168 5811 15407 5837
rect 15168 5777 15170 5811
rect 15204 5803 15407 5811
rect 15204 5777 15216 5803
rect 14418 5773 14517 5777
rect 14196 5715 14211 5749
rect 14162 5699 14211 5715
rect 14245 5743 14261 5757
rect 14245 5709 14246 5743
rect 14295 5723 14333 5757
rect 14418 5739 14501 5773
rect 14535 5739 14551 5773
rect 14585 5739 14601 5773
rect 14635 5743 14660 5773
rect 14280 5709 14333 5723
rect 14585 5709 14614 5739
rect 14648 5709 14660 5743
rect 14719 5714 14952 5771
rect 15373 5765 15407 5803
rect 15475 5835 15493 5869
rect 15441 5798 15493 5835
rect 14062 5629 14142 5667
rect 14062 5595 14108 5629
rect 14062 5539 14142 5595
rect 14177 5577 14211 5699
rect 14299 5645 14338 5675
rect 14299 5611 14333 5645
rect 14372 5641 14383 5675
rect 14719 5661 14753 5714
rect 14367 5611 14383 5641
rect 14429 5645 14686 5661
rect 14463 5627 14686 5645
rect 14720 5627 14753 5661
rect 14798 5675 14870 5677
rect 14832 5661 14870 5675
rect 14798 5627 14803 5641
rect 14837 5627 14870 5661
rect 14463 5611 14479 5627
rect 14798 5611 14870 5627
rect 14918 5645 14952 5714
rect 14986 5743 15064 5758
rect 15262 5749 15328 5765
rect 15262 5743 15294 5749
rect 15020 5742 15064 5743
rect 15020 5709 15030 5742
rect 14986 5708 15030 5709
rect 14986 5692 15064 5708
rect 15102 5709 15126 5743
rect 15160 5709 15176 5743
rect 15296 5709 15328 5715
rect 15102 5645 15136 5709
rect 15294 5699 15328 5709
rect 15373 5749 15424 5765
rect 15373 5715 15390 5749
rect 15373 5699 15424 5715
rect 14918 5611 15136 5645
rect 15204 5641 15250 5675
rect 15170 5638 15250 5641
rect 15373 5639 15407 5699
rect 15458 5667 15493 5798
rect 14429 5608 14479 5611
rect 14177 5543 14310 5577
rect 14429 5574 14436 5608
rect 14470 5574 14479 5608
rect 15170 5604 15216 5638
rect 15170 5588 15250 5604
rect 14429 5573 14479 5574
rect 14062 5505 14108 5539
rect 14276 5539 14310 5543
rect 14560 5543 14762 5577
rect 14276 5521 14493 5539
rect 14062 5471 14142 5505
rect 14176 5475 14192 5509
rect 14226 5475 14242 5509
rect 14176 5437 14242 5475
rect 14276 5487 14459 5521
rect 14276 5471 14493 5487
rect 14560 5526 14594 5543
rect 14728 5526 14762 5543
rect 14560 5471 14594 5492
rect 14628 5475 14644 5509
rect 14678 5475 14694 5509
rect 14628 5437 14694 5475
rect 14903 5543 15118 5577
rect 15289 5575 15407 5639
rect 15441 5626 15493 5667
rect 15475 5602 15493 5626
rect 15289 5551 15323 5575
rect 14903 5526 14950 5543
rect 14728 5471 14762 5492
rect 14796 5479 14812 5513
rect 14846 5479 14862 5513
rect 14796 5437 14862 5479
rect 14903 5492 14916 5526
rect 15084 5526 15118 5543
rect 14903 5471 14950 5492
rect 14984 5475 15000 5509
rect 15034 5475 15050 5509
rect 14984 5437 15050 5475
rect 15084 5471 15118 5492
rect 15168 5526 15323 5551
rect 15441 5566 15452 5592
rect 15486 5566 15493 5602
rect 15202 5492 15323 5526
rect 15168 5471 15323 5492
rect 15357 5517 15407 5534
rect 15391 5483 15407 5517
rect 15357 5437 15407 5483
rect 15441 5532 15493 5566
rect 15475 5498 15493 5532
rect 15441 5471 15493 5498
rect 16056 5875 16136 5919
rect 16185 5915 16251 5953
rect 16185 5881 16201 5915
rect 16235 5881 16251 5915
rect 16285 5903 16487 5919
rect 16056 5841 16102 5875
rect 16285 5869 16453 5903
rect 16285 5847 16319 5869
rect 16453 5851 16487 5869
rect 16554 5898 16588 5919
rect 16622 5915 16688 5953
rect 16622 5881 16638 5915
rect 16672 5881 16688 5915
rect 16722 5898 16756 5919
rect 16056 5808 16136 5841
rect 16171 5813 16319 5847
rect 16554 5847 16588 5864
rect 16790 5906 16856 5953
rect 16790 5872 16806 5906
rect 16840 5872 16856 5906
rect 16910 5898 16944 5919
rect 16722 5847 16756 5864
rect 16056 5673 16122 5808
rect 16171 5771 16205 5813
rect 16156 5755 16205 5771
rect 16412 5783 16424 5817
rect 16458 5783 16511 5817
rect 16554 5813 16756 5847
rect 16978 5915 17044 5953
rect 16978 5881 16994 5915
rect 17028 5881 17044 5915
rect 17078 5898 17112 5919
rect 16910 5847 16944 5864
rect 17078 5847 17112 5864
rect 16910 5813 17112 5847
rect 17162 5898 17282 5919
rect 17196 5864 17282 5898
rect 17335 5911 17401 5953
rect 17335 5877 17351 5911
rect 17385 5877 17401 5911
rect 17162 5843 17282 5864
rect 17435 5875 17487 5919
rect 17162 5817 17401 5843
rect 17162 5783 17164 5817
rect 17198 5809 17401 5817
rect 17198 5783 17210 5809
rect 16412 5779 16511 5783
rect 16190 5721 16205 5755
rect 16156 5705 16205 5721
rect 16239 5749 16255 5763
rect 16239 5715 16240 5749
rect 16289 5729 16327 5763
rect 16412 5745 16495 5779
rect 16529 5745 16545 5779
rect 16579 5745 16595 5779
rect 16629 5749 16654 5779
rect 16274 5715 16327 5729
rect 16579 5715 16608 5745
rect 16642 5715 16654 5749
rect 16713 5720 16946 5777
rect 17367 5771 17401 5809
rect 17469 5841 17487 5875
rect 17435 5804 17487 5841
rect 16056 5635 16136 5673
rect 16056 5601 16102 5635
rect 16056 5545 16136 5601
rect 16171 5583 16205 5705
rect 16293 5651 16332 5681
rect 16293 5617 16327 5651
rect 16366 5647 16377 5681
rect 16713 5667 16747 5720
rect 16361 5617 16377 5647
rect 16423 5651 16680 5667
rect 16457 5633 16680 5651
rect 16714 5633 16747 5667
rect 16792 5681 16864 5683
rect 16826 5667 16864 5681
rect 16792 5633 16797 5647
rect 16831 5633 16864 5667
rect 16457 5617 16473 5633
rect 16792 5617 16864 5633
rect 16912 5651 16946 5720
rect 16980 5749 17058 5764
rect 17256 5755 17322 5771
rect 17256 5749 17288 5755
rect 17014 5748 17058 5749
rect 17014 5715 17024 5748
rect 16980 5714 17024 5715
rect 16980 5698 17058 5714
rect 17096 5715 17120 5749
rect 17154 5715 17170 5749
rect 17290 5715 17322 5721
rect 17096 5651 17130 5715
rect 17288 5705 17322 5715
rect 17367 5755 17418 5771
rect 17367 5721 17384 5755
rect 17367 5705 17418 5721
rect 16912 5617 17130 5651
rect 17198 5647 17244 5681
rect 17164 5644 17244 5647
rect 17367 5645 17401 5705
rect 17452 5673 17487 5804
rect 16423 5614 16473 5617
rect 16171 5549 16304 5583
rect 16423 5580 16430 5614
rect 16464 5580 16473 5614
rect 17164 5610 17210 5644
rect 17164 5594 17244 5610
rect 16423 5579 16473 5580
rect 16056 5511 16102 5545
rect 16270 5545 16304 5549
rect 16554 5549 16756 5583
rect 16270 5527 16487 5545
rect 16056 5477 16136 5511
rect 16170 5481 16186 5515
rect 16220 5481 16236 5515
rect 16170 5443 16236 5481
rect 16270 5493 16453 5527
rect 16270 5477 16487 5493
rect 16554 5532 16588 5549
rect 16722 5532 16756 5549
rect 16554 5477 16588 5498
rect 16622 5481 16638 5515
rect 16672 5481 16688 5515
rect 16622 5443 16688 5481
rect 16897 5549 17112 5583
rect 17283 5581 17401 5645
rect 17435 5632 17487 5673
rect 17469 5608 17487 5632
rect 17283 5557 17317 5581
rect 16897 5532 16944 5549
rect 16722 5477 16756 5498
rect 16790 5485 16806 5519
rect 16840 5485 16856 5519
rect 16790 5443 16856 5485
rect 16897 5498 16910 5532
rect 17078 5532 17112 5549
rect 16897 5477 16944 5498
rect 16978 5481 16994 5515
rect 17028 5481 17044 5515
rect 16978 5443 17044 5481
rect 17078 5477 17112 5498
rect 17162 5532 17317 5557
rect 17435 5572 17446 5598
rect 17480 5572 17487 5608
rect 17196 5498 17317 5532
rect 17162 5477 17317 5498
rect 17351 5523 17401 5540
rect 17385 5489 17401 5523
rect 17351 5443 17401 5489
rect 17435 5538 17487 5572
rect 17469 5504 17487 5538
rect 17435 5477 17487 5504
rect 12080 5395 12109 5429
rect 12143 5395 12201 5429
rect 12235 5395 12293 5429
rect 12327 5395 12385 5429
rect 12419 5395 12477 5429
rect 12511 5395 12569 5429
rect 12603 5395 12661 5429
rect 12695 5395 12753 5429
rect 12787 5395 12845 5429
rect 12879 5395 12937 5429
rect 12971 5395 13029 5429
rect 13063 5395 13121 5429
rect 13155 5395 13213 5429
rect 13247 5395 13305 5429
rect 13339 5395 13397 5429
rect 13431 5395 13489 5429
rect 13523 5395 13552 5429
rect 14038 5403 14067 5437
rect 14101 5403 14159 5437
rect 14193 5403 14251 5437
rect 14285 5403 14343 5437
rect 14377 5403 14435 5437
rect 14469 5403 14527 5437
rect 14561 5403 14619 5437
rect 14653 5403 14711 5437
rect 14745 5403 14803 5437
rect 14837 5403 14895 5437
rect 14929 5403 14987 5437
rect 15021 5403 15079 5437
rect 15113 5403 15171 5437
rect 15205 5403 15263 5437
rect 15297 5403 15355 5437
rect 15389 5403 15447 5437
rect 15481 5403 15510 5437
rect 16032 5409 16061 5443
rect 16095 5409 16153 5443
rect 16187 5409 16245 5443
rect 16279 5409 16337 5443
rect 16371 5409 16429 5443
rect 16463 5409 16521 5443
rect 16555 5409 16613 5443
rect 16647 5409 16705 5443
rect 16739 5409 16797 5443
rect 16831 5409 16889 5443
rect 16923 5409 16981 5443
rect 17015 5409 17073 5443
rect 17107 5409 17165 5443
rect 17199 5409 17257 5443
rect 17291 5409 17349 5443
rect 17383 5409 17441 5443
rect 17475 5409 17504 5443
rect 7948 5211 8028 5249
rect 7948 5177 7994 5211
rect 7948 5121 8028 5177
rect 8063 5159 8097 5281
rect 8185 5227 8224 5257
rect 8185 5193 8219 5227
rect 8258 5223 8269 5257
rect 8605 5243 8639 5296
rect 8253 5193 8269 5223
rect 8315 5227 8572 5243
rect 8349 5209 8572 5227
rect 8606 5209 8639 5243
rect 8684 5257 8756 5259
rect 8718 5243 8756 5257
rect 8684 5209 8689 5223
rect 8723 5209 8756 5243
rect 8349 5193 8365 5209
rect 8684 5193 8756 5209
rect 8804 5227 8838 5296
rect 8872 5325 8950 5340
rect 9148 5331 9214 5347
rect 9148 5325 9180 5331
rect 8906 5324 8950 5325
rect 8906 5291 8916 5324
rect 8872 5290 8916 5291
rect 8872 5274 8950 5290
rect 8988 5291 9012 5325
rect 9046 5291 9062 5325
rect 9182 5291 9214 5297
rect 8988 5227 9022 5291
rect 9180 5281 9214 5291
rect 9259 5331 9310 5347
rect 9259 5297 9276 5331
rect 9259 5281 9310 5297
rect 8804 5193 9022 5227
rect 9090 5223 9136 5257
rect 9056 5220 9136 5223
rect 9259 5221 9293 5281
rect 9344 5249 9379 5380
rect 8315 5190 8365 5193
rect 8063 5125 8196 5159
rect 8315 5156 8322 5190
rect 8356 5156 8365 5190
rect 9056 5186 9102 5220
rect 9056 5170 9136 5186
rect 8315 5155 8365 5156
rect 7948 5087 7994 5121
rect 8162 5121 8196 5125
rect 8446 5125 8648 5159
rect 8162 5103 8379 5121
rect 7948 5053 8028 5087
rect 8062 5057 8078 5091
rect 8112 5057 8128 5091
rect 8062 5019 8128 5057
rect 8162 5069 8345 5103
rect 8162 5053 8379 5069
rect 8446 5108 8480 5125
rect 8614 5108 8648 5125
rect 8446 5053 8480 5074
rect 8514 5057 8530 5091
rect 8564 5057 8580 5091
rect 8514 5019 8580 5057
rect 8789 5125 9004 5159
rect 9175 5157 9293 5221
rect 9327 5208 9379 5249
rect 9361 5184 9379 5208
rect 9175 5133 9209 5157
rect 8789 5108 8836 5125
rect 8614 5053 8648 5074
rect 8682 5061 8698 5095
rect 8732 5061 8748 5095
rect 8682 5019 8748 5061
rect 8789 5074 8802 5108
rect 8970 5108 9004 5125
rect 8789 5053 8836 5074
rect 8870 5057 8886 5091
rect 8920 5057 8936 5091
rect 8870 5019 8936 5057
rect 8970 5053 9004 5074
rect 9054 5108 9209 5133
rect 9327 5148 9338 5174
rect 9372 5148 9379 5184
rect 9088 5074 9209 5108
rect 9054 5053 9209 5074
rect 9243 5099 9293 5116
rect 9277 5065 9293 5099
rect 9243 5019 9293 5065
rect 9327 5114 9379 5148
rect 9361 5080 9379 5114
rect 9327 5053 9379 5080
rect 10046 5077 10075 5111
rect 10109 5077 10167 5111
rect 10201 5077 10259 5111
rect 10293 5077 10351 5111
rect 10385 5077 10443 5111
rect 10477 5077 10535 5111
rect 10569 5077 10627 5111
rect 10661 5077 10719 5111
rect 10753 5077 10811 5111
rect 10845 5077 10903 5111
rect 10937 5077 10995 5111
rect 11029 5077 11087 5111
rect 11121 5077 11179 5111
rect 11213 5077 11271 5111
rect 11305 5077 11363 5111
rect 11397 5077 11455 5111
rect 11489 5077 11518 5111
rect 3970 4979 3999 5013
rect 4033 4979 4091 5013
rect 4125 4979 4183 5013
rect 4217 4979 4275 5013
rect 4309 4979 4367 5013
rect 4401 4979 4459 5013
rect 4493 4979 4551 5013
rect 4585 4979 4643 5013
rect 4677 4979 4735 5013
rect 4769 4979 4827 5013
rect 4861 4979 4919 5013
rect 4953 4979 5011 5013
rect 5045 4979 5103 5013
rect 5137 4979 5195 5013
rect 5229 4979 5287 5013
rect 5321 4979 5379 5013
rect 5413 4979 5442 5013
rect 5922 4979 5951 5013
rect 5985 4979 6043 5013
rect 6077 4979 6135 5013
rect 6169 4979 6227 5013
rect 6261 4979 6319 5013
rect 6353 4979 6411 5013
rect 6445 4979 6503 5013
rect 6537 4979 6595 5013
rect 6629 4979 6687 5013
rect 6721 4979 6779 5013
rect 6813 4979 6871 5013
rect 6905 4979 6963 5013
rect 6997 4979 7055 5013
rect 7089 4979 7147 5013
rect 7181 4979 7239 5013
rect 7273 4979 7331 5013
rect 7365 4979 7394 5013
rect 7924 4985 7953 5019
rect 7987 4985 8045 5019
rect 8079 4985 8137 5019
rect 8171 4985 8229 5019
rect 8263 4985 8321 5019
rect 8355 4985 8413 5019
rect 8447 4985 8505 5019
rect 8539 4985 8597 5019
rect 8631 4985 8689 5019
rect 8723 4985 8781 5019
rect 8815 4985 8873 5019
rect 8907 4985 8965 5019
rect 8999 4985 9057 5019
rect 9091 4985 9149 5019
rect 9183 4985 9241 5019
rect 9275 4985 9333 5019
rect 9367 4985 9396 5019
rect 10070 4999 10150 5043
rect 10199 5039 10265 5077
rect 10199 5005 10215 5039
rect 10249 5005 10265 5039
rect 10299 5027 10501 5043
rect 10070 4965 10116 4999
rect 10299 4993 10467 5027
rect 10299 4971 10333 4993
rect 10467 4975 10501 4993
rect 10568 5022 10602 5043
rect 10636 5039 10702 5077
rect 10636 5005 10652 5039
rect 10686 5005 10702 5039
rect 10736 5022 10770 5043
rect 10070 4932 10150 4965
rect 10185 4937 10333 4971
rect 10568 4971 10602 4988
rect 10804 5030 10870 5077
rect 10804 4996 10820 5030
rect 10854 4996 10870 5030
rect 10924 5022 10958 5043
rect 10736 4971 10770 4988
rect 10070 4797 10136 4932
rect 10185 4895 10219 4937
rect 10170 4879 10219 4895
rect 10426 4907 10438 4941
rect 10472 4907 10525 4941
rect 10568 4937 10770 4971
rect 10992 5039 11058 5077
rect 10992 5005 11008 5039
rect 11042 5005 11058 5039
rect 11092 5022 11126 5043
rect 10924 4971 10958 4988
rect 11092 4971 11126 4988
rect 10924 4937 11126 4971
rect 11176 5022 11296 5043
rect 11210 4988 11296 5022
rect 11349 5035 11415 5077
rect 11349 5001 11365 5035
rect 11399 5001 11415 5035
rect 11176 4967 11296 4988
rect 11449 4999 11501 5043
rect 12316 5033 12345 5067
rect 12379 5033 12437 5067
rect 12471 5033 12529 5067
rect 12563 5033 12621 5067
rect 12655 5033 12713 5067
rect 12747 5033 12805 5067
rect 12839 5033 12897 5067
rect 12931 5033 12989 5067
rect 13023 5033 13081 5067
rect 13115 5033 13173 5067
rect 13207 5033 13265 5067
rect 13299 5033 13357 5067
rect 13391 5033 13449 5067
rect 13483 5033 13541 5067
rect 13575 5033 13633 5067
rect 13667 5033 13725 5067
rect 13759 5033 13788 5067
rect 11176 4941 11415 4967
rect 11176 4907 11178 4941
rect 11212 4933 11415 4941
rect 11212 4907 11224 4933
rect 10426 4903 10525 4907
rect 10204 4845 10219 4879
rect 10170 4829 10219 4845
rect 10253 4873 10269 4887
rect 10253 4839 10254 4873
rect 10303 4853 10341 4887
rect 10426 4869 10509 4903
rect 10543 4869 10559 4903
rect 10593 4869 10609 4903
rect 10643 4873 10668 4903
rect 10288 4839 10341 4853
rect 10593 4839 10622 4869
rect 10656 4839 10668 4873
rect 10727 4844 10960 4901
rect 11381 4895 11415 4933
rect 11483 4965 11501 4999
rect 11449 4928 11501 4965
rect 10070 4759 10150 4797
rect 10070 4725 10116 4759
rect 10070 4669 10150 4725
rect 10185 4707 10219 4829
rect 10307 4775 10346 4805
rect 10307 4741 10341 4775
rect 10380 4771 10391 4805
rect 10727 4791 10761 4844
rect 10375 4741 10391 4771
rect 10437 4775 10694 4791
rect 10471 4757 10694 4775
rect 10728 4757 10761 4791
rect 10806 4805 10878 4807
rect 10840 4791 10878 4805
rect 10806 4757 10811 4771
rect 10845 4757 10878 4791
rect 10471 4741 10487 4757
rect 10806 4741 10878 4757
rect 10926 4775 10960 4844
rect 10994 4873 11072 4888
rect 11270 4879 11336 4895
rect 11270 4873 11302 4879
rect 11028 4872 11072 4873
rect 11028 4839 11038 4872
rect 10994 4838 11038 4839
rect 10994 4822 11072 4838
rect 11110 4839 11134 4873
rect 11168 4839 11184 4873
rect 11304 4839 11336 4845
rect 11110 4775 11144 4839
rect 11302 4829 11336 4839
rect 11381 4879 11432 4895
rect 11381 4845 11398 4879
rect 11381 4829 11432 4845
rect 10926 4741 11144 4775
rect 11212 4771 11258 4805
rect 11178 4768 11258 4771
rect 11381 4769 11415 4829
rect 11466 4797 11501 4928
rect 10437 4740 10487 4741
rect 10185 4673 10318 4707
rect 10437 4706 10446 4740
rect 10480 4706 10487 4740
rect 11178 4734 11224 4768
rect 11178 4718 11258 4734
rect 10437 4703 10487 4706
rect 10070 4635 10116 4669
rect 10284 4669 10318 4673
rect 10568 4673 10770 4707
rect 10284 4651 10501 4669
rect 10070 4601 10150 4635
rect 10184 4605 10200 4639
rect 10234 4605 10250 4639
rect 10184 4567 10250 4605
rect 10284 4617 10467 4651
rect 10284 4601 10501 4617
rect 10568 4656 10602 4673
rect 10736 4656 10770 4673
rect 10568 4601 10602 4622
rect 10636 4605 10652 4639
rect 10686 4605 10702 4639
rect 10636 4567 10702 4605
rect 10911 4673 11126 4707
rect 11297 4705 11415 4769
rect 11449 4756 11501 4797
rect 11483 4732 11501 4756
rect 11297 4681 11331 4705
rect 10911 4656 10958 4673
rect 10736 4601 10770 4622
rect 10804 4609 10820 4643
rect 10854 4609 10870 4643
rect 10804 4567 10870 4609
rect 10911 4622 10924 4656
rect 11092 4656 11126 4673
rect 10911 4601 10958 4622
rect 10992 4605 11008 4639
rect 11042 4605 11058 4639
rect 10992 4567 11058 4605
rect 11092 4601 11126 4622
rect 11176 4656 11331 4681
rect 11449 4696 11454 4722
rect 11494 4696 11501 4732
rect 11210 4622 11331 4656
rect 11176 4601 11331 4622
rect 11365 4647 11415 4664
rect 11399 4613 11415 4647
rect 11365 4567 11415 4613
rect 11449 4662 11501 4696
rect 11483 4628 11501 4662
rect 11449 4601 11501 4628
rect 12340 4955 12420 4999
rect 12469 4995 12535 5033
rect 12469 4961 12485 4995
rect 12519 4961 12535 4995
rect 12569 4983 12771 4999
rect 12340 4921 12386 4955
rect 12569 4949 12737 4983
rect 12569 4927 12603 4949
rect 12737 4931 12771 4949
rect 12838 4978 12872 4999
rect 12906 4995 12972 5033
rect 12906 4961 12922 4995
rect 12956 4961 12972 4995
rect 13006 4978 13040 4999
rect 12340 4888 12420 4921
rect 12455 4893 12603 4927
rect 12838 4927 12872 4944
rect 13074 4986 13140 5033
rect 13074 4952 13090 4986
rect 13124 4952 13140 4986
rect 13194 4978 13228 4999
rect 13006 4927 13040 4944
rect 12340 4753 12406 4888
rect 12455 4851 12489 4893
rect 12440 4835 12489 4851
rect 12696 4863 12708 4897
rect 12742 4863 12795 4897
rect 12838 4893 13040 4927
rect 13262 4995 13328 5033
rect 13262 4961 13278 4995
rect 13312 4961 13328 4995
rect 13362 4978 13396 4999
rect 13194 4927 13228 4944
rect 13362 4927 13396 4944
rect 13194 4893 13396 4927
rect 13446 4978 13566 4999
rect 13480 4944 13566 4978
rect 13619 4991 13685 5033
rect 14318 5027 14347 5061
rect 14381 5027 14439 5061
rect 14473 5027 14531 5061
rect 14565 5027 14623 5061
rect 14657 5027 14715 5061
rect 14749 5027 14807 5061
rect 14841 5027 14899 5061
rect 14933 5027 14991 5061
rect 15025 5027 15083 5061
rect 15117 5027 15175 5061
rect 15209 5027 15267 5061
rect 15301 5027 15359 5061
rect 15393 5027 15451 5061
rect 15485 5027 15543 5061
rect 15577 5027 15635 5061
rect 15669 5027 15727 5061
rect 15761 5027 15790 5061
rect 13619 4957 13635 4991
rect 13669 4957 13685 4991
rect 13446 4923 13566 4944
rect 13719 4955 13771 4999
rect 13446 4897 13685 4923
rect 13446 4863 13448 4897
rect 13482 4889 13685 4897
rect 13482 4863 13494 4889
rect 12696 4859 12795 4863
rect 12474 4801 12489 4835
rect 12440 4785 12489 4801
rect 12523 4829 12539 4843
rect 12523 4795 12524 4829
rect 12573 4809 12611 4843
rect 12696 4825 12779 4859
rect 12813 4825 12829 4859
rect 12863 4825 12879 4859
rect 12913 4829 12938 4859
rect 12558 4795 12611 4809
rect 12863 4795 12892 4825
rect 12926 4795 12938 4829
rect 12997 4800 13230 4857
rect 13651 4851 13685 4889
rect 13753 4921 13771 4955
rect 13719 4884 13771 4921
rect 12340 4715 12420 4753
rect 12340 4681 12386 4715
rect 12340 4625 12420 4681
rect 12455 4663 12489 4785
rect 12577 4731 12616 4761
rect 12577 4697 12611 4731
rect 12650 4727 12661 4761
rect 12997 4747 13031 4800
rect 12645 4697 12661 4727
rect 12707 4731 12964 4747
rect 12741 4713 12964 4731
rect 12998 4713 13031 4747
rect 13076 4761 13148 4763
rect 13110 4747 13148 4761
rect 13076 4713 13081 4727
rect 13115 4713 13148 4747
rect 12741 4697 12757 4713
rect 13076 4697 13148 4713
rect 13196 4731 13230 4800
rect 13264 4829 13342 4844
rect 13540 4835 13606 4851
rect 13540 4829 13572 4835
rect 13298 4828 13342 4829
rect 13298 4795 13308 4828
rect 13264 4794 13308 4795
rect 13264 4778 13342 4794
rect 13380 4795 13404 4829
rect 13438 4795 13454 4829
rect 13574 4795 13606 4801
rect 13380 4731 13414 4795
rect 13572 4785 13606 4795
rect 13651 4835 13702 4851
rect 13651 4801 13668 4835
rect 13651 4785 13702 4801
rect 13196 4697 13414 4731
rect 13482 4727 13528 4761
rect 13448 4724 13528 4727
rect 13651 4725 13685 4785
rect 13736 4753 13771 4884
rect 12707 4694 12757 4697
rect 12455 4629 12588 4663
rect 12707 4660 12714 4694
rect 12748 4660 12757 4694
rect 13448 4690 13494 4724
rect 13448 4674 13528 4690
rect 12707 4659 12757 4660
rect 12340 4591 12386 4625
rect 12554 4625 12588 4629
rect 12838 4629 13040 4663
rect 12554 4607 12771 4625
rect 10046 4533 10075 4567
rect 10109 4533 10167 4567
rect 10201 4533 10259 4567
rect 10293 4533 10351 4567
rect 10385 4533 10443 4567
rect 10477 4533 10535 4567
rect 10569 4533 10627 4567
rect 10661 4533 10719 4567
rect 10753 4533 10811 4567
rect 10845 4533 10903 4567
rect 10937 4533 10995 4567
rect 11029 4533 11087 4567
rect 11121 4533 11179 4567
rect 11213 4533 11271 4567
rect 11305 4533 11363 4567
rect 11397 4533 11455 4567
rect 11489 4533 11518 4567
rect 12340 4557 12420 4591
rect 12454 4561 12470 4595
rect 12504 4561 12520 4595
rect 12454 4523 12520 4561
rect 12554 4573 12737 4607
rect 12554 4557 12771 4573
rect 12838 4612 12872 4629
rect 13006 4612 13040 4629
rect 12838 4557 12872 4578
rect 12906 4561 12922 4595
rect 12956 4561 12972 4595
rect 12906 4523 12972 4561
rect 13181 4629 13396 4663
rect 13567 4661 13685 4725
rect 13719 4712 13771 4753
rect 13753 4688 13771 4712
rect 13567 4637 13601 4661
rect 13181 4612 13228 4629
rect 13006 4557 13040 4578
rect 13074 4565 13090 4599
rect 13124 4565 13140 4599
rect 13074 4523 13140 4565
rect 13181 4578 13194 4612
rect 13362 4612 13396 4629
rect 13181 4557 13228 4578
rect 13262 4561 13278 4595
rect 13312 4561 13328 4595
rect 13262 4523 13328 4561
rect 13362 4557 13396 4578
rect 13446 4612 13601 4637
rect 13719 4652 13730 4678
rect 13764 4652 13771 4688
rect 13480 4578 13601 4612
rect 13446 4557 13601 4578
rect 13635 4603 13685 4620
rect 13669 4569 13685 4603
rect 13635 4523 13685 4569
rect 13719 4618 13771 4652
rect 13753 4584 13771 4618
rect 13719 4557 13771 4584
rect 14342 4949 14422 4993
rect 14471 4989 14537 5027
rect 14471 4955 14487 4989
rect 14521 4955 14537 4989
rect 14571 4977 14773 4993
rect 14342 4915 14388 4949
rect 14571 4943 14739 4977
rect 14571 4921 14605 4943
rect 14739 4925 14773 4943
rect 14840 4972 14874 4993
rect 14908 4989 14974 5027
rect 14908 4955 14924 4989
rect 14958 4955 14974 4989
rect 15008 4972 15042 4993
rect 14342 4882 14422 4915
rect 14457 4887 14605 4921
rect 14840 4921 14874 4938
rect 15076 4980 15142 5027
rect 15076 4946 15092 4980
rect 15126 4946 15142 4980
rect 15196 4972 15230 4993
rect 15008 4921 15042 4938
rect 14342 4747 14408 4882
rect 14457 4845 14491 4887
rect 14442 4829 14491 4845
rect 14698 4857 14710 4891
rect 14744 4857 14797 4891
rect 14840 4887 15042 4921
rect 15264 4989 15330 5027
rect 15264 4955 15280 4989
rect 15314 4955 15330 4989
rect 15364 4972 15398 4993
rect 15196 4921 15230 4938
rect 15364 4921 15398 4938
rect 15196 4887 15398 4921
rect 15448 4972 15568 4993
rect 15482 4938 15568 4972
rect 15621 4985 15687 5027
rect 16340 5009 16369 5043
rect 16403 5009 16461 5043
rect 16495 5009 16553 5043
rect 16587 5009 16645 5043
rect 16679 5009 16737 5043
rect 16771 5009 16829 5043
rect 16863 5009 16921 5043
rect 16955 5009 17013 5043
rect 17047 5009 17105 5043
rect 17139 5009 17197 5043
rect 17231 5009 17289 5043
rect 17323 5009 17381 5043
rect 17415 5009 17473 5043
rect 17507 5009 17565 5043
rect 17599 5009 17657 5043
rect 17691 5009 17749 5043
rect 17783 5009 17812 5043
rect 15621 4951 15637 4985
rect 15671 4951 15687 4985
rect 15448 4917 15568 4938
rect 15721 4949 15773 4993
rect 15448 4891 15687 4917
rect 15448 4857 15450 4891
rect 15484 4883 15687 4891
rect 15484 4857 15496 4883
rect 14698 4853 14797 4857
rect 14476 4795 14491 4829
rect 14442 4779 14491 4795
rect 14525 4823 14541 4837
rect 14525 4789 14526 4823
rect 14575 4803 14613 4837
rect 14698 4819 14781 4853
rect 14815 4819 14831 4853
rect 14865 4819 14881 4853
rect 14915 4823 14940 4853
rect 14560 4789 14613 4803
rect 14865 4789 14894 4819
rect 14928 4789 14940 4823
rect 14999 4794 15232 4851
rect 15653 4845 15687 4883
rect 15755 4915 15773 4949
rect 15721 4878 15773 4915
rect 14342 4709 14422 4747
rect 14342 4675 14388 4709
rect 14342 4619 14422 4675
rect 14457 4657 14491 4779
rect 14579 4725 14618 4755
rect 14579 4691 14613 4725
rect 14652 4721 14663 4755
rect 14999 4741 15033 4794
rect 14647 4691 14663 4721
rect 14709 4725 14966 4741
rect 14743 4707 14966 4725
rect 15000 4707 15033 4741
rect 15078 4755 15150 4757
rect 15112 4741 15150 4755
rect 15078 4707 15083 4721
rect 15117 4707 15150 4741
rect 14743 4691 14759 4707
rect 15078 4691 15150 4707
rect 15198 4725 15232 4794
rect 15266 4823 15344 4838
rect 15542 4829 15608 4845
rect 15542 4823 15574 4829
rect 15300 4822 15344 4823
rect 15300 4789 15310 4822
rect 15266 4788 15310 4789
rect 15266 4772 15344 4788
rect 15382 4789 15406 4823
rect 15440 4789 15456 4823
rect 15576 4789 15608 4795
rect 15382 4725 15416 4789
rect 15574 4779 15608 4789
rect 15653 4829 15704 4845
rect 15653 4795 15670 4829
rect 15653 4779 15704 4795
rect 15198 4691 15416 4725
rect 15484 4721 15530 4755
rect 15450 4718 15530 4721
rect 15653 4719 15687 4779
rect 15738 4747 15773 4878
rect 14709 4688 14759 4691
rect 14457 4623 14590 4657
rect 14709 4654 14716 4688
rect 14750 4654 14759 4688
rect 15450 4684 15496 4718
rect 15450 4668 15530 4684
rect 14709 4653 14759 4654
rect 14342 4585 14388 4619
rect 14556 4619 14590 4623
rect 14840 4623 15042 4657
rect 14556 4601 14773 4619
rect 14342 4551 14422 4585
rect 14456 4555 14472 4589
rect 14506 4555 14522 4589
rect 12316 4489 12345 4523
rect 12379 4489 12437 4523
rect 12471 4489 12529 4523
rect 12563 4489 12621 4523
rect 12655 4489 12713 4523
rect 12747 4489 12805 4523
rect 12839 4489 12897 4523
rect 12931 4489 12989 4523
rect 13023 4489 13081 4523
rect 13115 4489 13173 4523
rect 13207 4489 13265 4523
rect 13299 4489 13357 4523
rect 13391 4489 13449 4523
rect 13483 4489 13541 4523
rect 13575 4489 13633 4523
rect 13667 4489 13725 4523
rect 13759 4489 13788 4523
rect 14456 4517 14522 4555
rect 14556 4567 14739 4601
rect 14556 4551 14773 4567
rect 14840 4606 14874 4623
rect 15008 4606 15042 4623
rect 14840 4551 14874 4572
rect 14908 4555 14924 4589
rect 14958 4555 14974 4589
rect 14908 4517 14974 4555
rect 15183 4623 15398 4657
rect 15569 4655 15687 4719
rect 15721 4706 15773 4747
rect 15755 4682 15773 4706
rect 15569 4631 15603 4655
rect 15183 4606 15230 4623
rect 15008 4551 15042 4572
rect 15076 4559 15092 4593
rect 15126 4559 15142 4593
rect 15076 4517 15142 4559
rect 15183 4572 15196 4606
rect 15364 4606 15398 4623
rect 15183 4551 15230 4572
rect 15264 4555 15280 4589
rect 15314 4555 15330 4589
rect 15264 4517 15330 4555
rect 15364 4551 15398 4572
rect 15448 4606 15603 4631
rect 15721 4646 15732 4672
rect 15766 4646 15773 4682
rect 15482 4572 15603 4606
rect 15448 4551 15603 4572
rect 15637 4597 15687 4614
rect 15671 4563 15687 4597
rect 15637 4517 15687 4563
rect 15721 4612 15773 4646
rect 15755 4578 15773 4612
rect 15721 4551 15773 4578
rect 16364 4931 16444 4975
rect 16493 4971 16559 5009
rect 16493 4937 16509 4971
rect 16543 4937 16559 4971
rect 16593 4959 16795 4975
rect 16364 4897 16410 4931
rect 16593 4925 16761 4959
rect 16593 4903 16627 4925
rect 16761 4907 16795 4925
rect 16862 4954 16896 4975
rect 16930 4971 16996 5009
rect 16930 4937 16946 4971
rect 16980 4937 16996 4971
rect 17030 4954 17064 4975
rect 16364 4864 16444 4897
rect 16479 4869 16627 4903
rect 16862 4903 16896 4920
rect 17098 4962 17164 5009
rect 17098 4928 17114 4962
rect 17148 4928 17164 4962
rect 17218 4954 17252 4975
rect 17030 4903 17064 4920
rect 16364 4729 16430 4864
rect 16479 4827 16513 4869
rect 16464 4811 16513 4827
rect 16720 4839 16732 4873
rect 16766 4839 16819 4873
rect 16862 4869 17064 4903
rect 17286 4971 17352 5009
rect 17286 4937 17302 4971
rect 17336 4937 17352 4971
rect 17386 4954 17420 4975
rect 17218 4903 17252 4920
rect 17386 4903 17420 4920
rect 17218 4869 17420 4903
rect 17470 4954 17590 4975
rect 17504 4920 17590 4954
rect 17643 4967 17709 5009
rect 17643 4933 17659 4967
rect 17693 4933 17709 4967
rect 17470 4899 17590 4920
rect 17743 4931 17795 4975
rect 17470 4873 17709 4899
rect 17470 4839 17472 4873
rect 17506 4865 17709 4873
rect 17506 4839 17518 4865
rect 16720 4835 16819 4839
rect 16498 4777 16513 4811
rect 16464 4761 16513 4777
rect 16547 4805 16563 4819
rect 16547 4771 16548 4805
rect 16597 4785 16635 4819
rect 16720 4801 16803 4835
rect 16837 4801 16853 4835
rect 16887 4801 16903 4835
rect 16937 4805 16962 4835
rect 16582 4771 16635 4785
rect 16887 4771 16916 4801
rect 16950 4771 16962 4805
rect 17021 4776 17254 4833
rect 17675 4827 17709 4865
rect 17777 4897 17795 4931
rect 17743 4860 17795 4897
rect 16364 4691 16444 4729
rect 16364 4657 16410 4691
rect 16364 4601 16444 4657
rect 16479 4639 16513 4761
rect 16601 4707 16640 4737
rect 16601 4673 16635 4707
rect 16674 4703 16685 4737
rect 17021 4723 17055 4776
rect 16669 4673 16685 4703
rect 16731 4707 16988 4723
rect 16765 4689 16988 4707
rect 17022 4689 17055 4723
rect 17100 4737 17172 4739
rect 17134 4723 17172 4737
rect 17100 4689 17105 4703
rect 17139 4689 17172 4723
rect 16765 4673 16781 4689
rect 17100 4673 17172 4689
rect 17220 4707 17254 4776
rect 17288 4805 17366 4820
rect 17564 4811 17630 4827
rect 17564 4805 17596 4811
rect 17322 4804 17366 4805
rect 17322 4771 17332 4804
rect 17288 4770 17332 4771
rect 17288 4754 17366 4770
rect 17404 4771 17428 4805
rect 17462 4771 17478 4805
rect 17598 4771 17630 4777
rect 17404 4707 17438 4771
rect 17596 4761 17630 4771
rect 17675 4811 17726 4827
rect 17675 4777 17692 4811
rect 17675 4761 17726 4777
rect 17220 4673 17438 4707
rect 17506 4703 17552 4737
rect 17472 4700 17552 4703
rect 17675 4701 17709 4761
rect 17760 4729 17795 4860
rect 16731 4670 16781 4673
rect 16479 4605 16612 4639
rect 16731 4636 16738 4670
rect 16772 4636 16781 4670
rect 17472 4666 17518 4700
rect 17472 4650 17552 4666
rect 16731 4635 16781 4636
rect 16364 4567 16410 4601
rect 16578 4601 16612 4605
rect 16862 4605 17064 4639
rect 16578 4583 16795 4601
rect 16364 4533 16444 4567
rect 16478 4537 16494 4571
rect 16528 4537 16544 4571
rect 14318 4483 14347 4517
rect 14381 4483 14439 4517
rect 14473 4483 14531 4517
rect 14565 4483 14623 4517
rect 14657 4483 14715 4517
rect 14749 4483 14807 4517
rect 14841 4483 14899 4517
rect 14933 4483 14991 4517
rect 15025 4483 15083 4517
rect 15117 4483 15175 4517
rect 15209 4483 15267 4517
rect 15301 4483 15359 4517
rect 15393 4483 15451 4517
rect 15485 4483 15543 4517
rect 15577 4483 15635 4517
rect 15669 4483 15727 4517
rect 15761 4483 15790 4517
rect 16478 4499 16544 4537
rect 16578 4549 16761 4583
rect 16578 4533 16795 4549
rect 16862 4588 16896 4605
rect 17030 4588 17064 4605
rect 16862 4533 16896 4554
rect 16930 4537 16946 4571
rect 16980 4537 16996 4571
rect 16930 4499 16996 4537
rect 17205 4605 17420 4639
rect 17591 4637 17709 4701
rect 17743 4688 17795 4729
rect 17777 4664 17795 4688
rect 17591 4613 17625 4637
rect 17205 4588 17252 4605
rect 17030 4533 17064 4554
rect 17098 4541 17114 4575
rect 17148 4541 17164 4575
rect 17098 4499 17164 4541
rect 17205 4554 17218 4588
rect 17386 4588 17420 4605
rect 17205 4533 17252 4554
rect 17286 4537 17302 4571
rect 17336 4537 17352 4571
rect 17286 4499 17352 4537
rect 17386 4533 17420 4554
rect 17470 4588 17625 4613
rect 17743 4628 17754 4654
rect 17788 4628 17795 4664
rect 17504 4554 17625 4588
rect 17470 4533 17625 4554
rect 17659 4579 17709 4596
rect 17693 4545 17709 4579
rect 17659 4499 17709 4545
rect 17743 4594 17795 4628
rect 17777 4560 17795 4594
rect 17743 4533 17795 4560
rect 16340 4465 16369 4499
rect 16403 4465 16461 4499
rect 16495 4465 16553 4499
rect 16587 4465 16645 4499
rect 16679 4465 16737 4499
rect 16771 4465 16829 4499
rect 16863 4465 16921 4499
rect 16955 4465 17013 4499
rect 17047 4465 17105 4499
rect 17139 4465 17197 4499
rect 17231 4465 17289 4499
rect 17323 4465 17381 4499
rect 17415 4465 17473 4499
rect 17507 4465 17565 4499
rect 17599 4465 17657 4499
rect 17691 4465 17749 4499
rect 17783 4465 17812 4499
rect 1806 2271 1835 2305
rect 1869 2271 1927 2305
rect 1961 2271 2019 2305
rect 2053 2271 2111 2305
rect 2145 2271 2203 2305
rect 2237 2271 2295 2305
rect 2329 2271 2387 2305
rect 2421 2271 2479 2305
rect 2513 2271 2571 2305
rect 2605 2271 2663 2305
rect 2697 2271 2755 2305
rect 2789 2271 2847 2305
rect 2881 2271 2939 2305
rect 2973 2271 3031 2305
rect 3065 2271 3123 2305
rect 3157 2271 3215 2305
rect 3249 2271 3278 2305
rect 1830 2193 1910 2237
rect 1959 2233 2025 2271
rect 1959 2199 1975 2233
rect 2009 2199 2025 2233
rect 2059 2221 2261 2237
rect 1830 2159 1876 2193
rect 2059 2187 2227 2221
rect 2059 2165 2093 2187
rect 2227 2169 2261 2187
rect 2328 2216 2362 2237
rect 2396 2233 2462 2271
rect 2396 2199 2412 2233
rect 2446 2199 2462 2233
rect 2496 2216 2530 2237
rect 1830 2126 1910 2159
rect 1945 2131 2093 2165
rect 2328 2165 2362 2182
rect 2564 2224 2630 2271
rect 2564 2190 2580 2224
rect 2614 2190 2630 2224
rect 2684 2216 2718 2237
rect 2496 2165 2530 2182
rect 1830 1991 1896 2126
rect 1945 2089 1979 2131
rect 1930 2073 1979 2089
rect 2186 2101 2198 2135
rect 2232 2101 2285 2135
rect 2328 2131 2530 2165
rect 2752 2233 2818 2271
rect 2752 2199 2768 2233
rect 2802 2199 2818 2233
rect 2852 2216 2886 2237
rect 2684 2165 2718 2182
rect 2852 2165 2886 2182
rect 2684 2131 2886 2165
rect 2936 2216 3056 2237
rect 2970 2182 3056 2216
rect 3109 2229 3175 2271
rect 3876 2267 3905 2301
rect 3939 2267 3997 2301
rect 4031 2267 4089 2301
rect 4123 2267 4181 2301
rect 4215 2267 4273 2301
rect 4307 2267 4365 2301
rect 4399 2267 4457 2301
rect 4491 2267 4549 2301
rect 4583 2267 4641 2301
rect 4675 2267 4733 2301
rect 4767 2267 4825 2301
rect 4859 2267 4917 2301
rect 4951 2267 5009 2301
rect 5043 2267 5101 2301
rect 5135 2267 5193 2301
rect 5227 2267 5285 2301
rect 5319 2267 5348 2301
rect 5828 2267 5857 2301
rect 5891 2267 5949 2301
rect 5983 2267 6041 2301
rect 6075 2267 6133 2301
rect 6167 2267 6225 2301
rect 6259 2267 6317 2301
rect 6351 2267 6409 2301
rect 6443 2267 6501 2301
rect 6535 2267 6593 2301
rect 6627 2267 6685 2301
rect 6719 2267 6777 2301
rect 6811 2267 6869 2301
rect 6903 2267 6961 2301
rect 6995 2267 7053 2301
rect 7087 2267 7145 2301
rect 7179 2267 7237 2301
rect 7271 2267 7300 2301
rect 7830 2273 7859 2307
rect 7893 2273 7951 2307
rect 7985 2273 8043 2307
rect 8077 2273 8135 2307
rect 8169 2273 8227 2307
rect 8261 2273 8319 2307
rect 8353 2273 8411 2307
rect 8445 2273 8503 2307
rect 8537 2273 8595 2307
rect 8629 2273 8687 2307
rect 8721 2273 8779 2307
rect 8813 2273 8871 2307
rect 8905 2273 8963 2307
rect 8997 2273 9055 2307
rect 9089 2273 9147 2307
rect 9181 2273 9239 2307
rect 9273 2273 9302 2307
rect 9782 2273 9811 2307
rect 9845 2273 9903 2307
rect 9937 2273 9995 2307
rect 10029 2273 10087 2307
rect 10121 2273 10179 2307
rect 10213 2273 10271 2307
rect 10305 2273 10363 2307
rect 10397 2273 10455 2307
rect 10489 2273 10547 2307
rect 10581 2273 10639 2307
rect 10673 2273 10731 2307
rect 10765 2273 10823 2307
rect 10857 2273 10915 2307
rect 10949 2273 11007 2307
rect 11041 2273 11099 2307
rect 11133 2273 11191 2307
rect 11225 2273 11254 2307
rect 11774 2273 11803 2307
rect 11837 2273 11895 2307
rect 11929 2273 11987 2307
rect 12021 2273 12079 2307
rect 12113 2273 12171 2307
rect 12205 2273 12263 2307
rect 12297 2273 12355 2307
rect 12389 2273 12447 2307
rect 12481 2273 12539 2307
rect 12573 2273 12631 2307
rect 12665 2273 12723 2307
rect 12757 2273 12815 2307
rect 12849 2273 12907 2307
rect 12941 2273 12999 2307
rect 13033 2273 13091 2307
rect 13125 2273 13183 2307
rect 13217 2273 13246 2307
rect 13726 2273 13755 2307
rect 13789 2273 13847 2307
rect 13881 2273 13939 2307
rect 13973 2273 14031 2307
rect 14065 2273 14123 2307
rect 14157 2273 14215 2307
rect 14249 2273 14307 2307
rect 14341 2273 14399 2307
rect 14433 2273 14491 2307
rect 14525 2273 14583 2307
rect 14617 2273 14675 2307
rect 14709 2273 14767 2307
rect 14801 2273 14859 2307
rect 14893 2273 14951 2307
rect 14985 2273 15043 2307
rect 15077 2273 15135 2307
rect 15169 2273 15198 2307
rect 15790 2273 15819 2307
rect 15853 2273 15911 2307
rect 15945 2273 16003 2307
rect 16037 2273 16095 2307
rect 16129 2273 16187 2307
rect 16221 2273 16279 2307
rect 16313 2273 16371 2307
rect 16405 2273 16463 2307
rect 16497 2273 16555 2307
rect 16589 2273 16647 2307
rect 16681 2273 16739 2307
rect 16773 2273 16831 2307
rect 16865 2273 16923 2307
rect 16957 2273 17015 2307
rect 17049 2273 17107 2307
rect 17141 2273 17199 2307
rect 17233 2273 17262 2307
rect 3109 2195 3125 2229
rect 3159 2195 3175 2229
rect 2936 2161 3056 2182
rect 3209 2193 3261 2237
rect 2936 2135 3175 2161
rect 2936 2101 2938 2135
rect 2972 2127 3175 2135
rect 2972 2101 2984 2127
rect 2186 2097 2285 2101
rect 1964 2039 1979 2073
rect 1930 2023 1979 2039
rect 2013 2067 2029 2081
rect 2013 2033 2014 2067
rect 2063 2047 2101 2081
rect 2186 2063 2269 2097
rect 2303 2063 2319 2097
rect 2353 2063 2369 2097
rect 2403 2067 2428 2097
rect 2048 2033 2101 2047
rect 2353 2033 2382 2063
rect 2416 2033 2428 2067
rect 2487 2038 2720 2095
rect 3141 2089 3175 2127
rect 3243 2159 3261 2193
rect 3209 2122 3261 2159
rect 1830 1953 1910 1991
rect 1830 1919 1876 1953
rect 1830 1863 1910 1919
rect 1945 1901 1979 2023
rect 2067 1969 2106 1999
rect 2067 1935 2101 1969
rect 2140 1965 2151 1999
rect 2487 1985 2521 2038
rect 2135 1935 2151 1965
rect 2197 1969 2454 1985
rect 2231 1951 2454 1969
rect 2488 1951 2521 1985
rect 2566 1999 2638 2001
rect 2600 1985 2638 1999
rect 2566 1951 2571 1965
rect 2605 1951 2638 1985
rect 2231 1935 2247 1951
rect 2566 1935 2638 1951
rect 2686 1969 2720 2038
rect 2754 2067 2832 2082
rect 3030 2073 3096 2089
rect 3030 2067 3062 2073
rect 2788 2066 2832 2067
rect 2788 2033 2798 2066
rect 2754 2032 2798 2033
rect 2754 2016 2832 2032
rect 2870 2033 2894 2067
rect 2928 2033 2944 2067
rect 3064 2033 3096 2039
rect 2870 1969 2904 2033
rect 3062 2023 3096 2033
rect 3141 2073 3192 2089
rect 3141 2039 3158 2073
rect 3141 2023 3192 2039
rect 2686 1935 2904 1969
rect 2972 1965 3018 1999
rect 2938 1962 3018 1965
rect 3141 1963 3175 2023
rect 3226 1991 3261 2122
rect 2197 1934 2247 1935
rect 1945 1867 2078 1901
rect 2197 1900 2206 1934
rect 2240 1900 2247 1934
rect 2938 1928 2984 1962
rect 2938 1912 3018 1928
rect 2197 1897 2247 1900
rect 1830 1829 1876 1863
rect 2044 1863 2078 1867
rect 2328 1867 2530 1901
rect 2044 1845 2261 1863
rect 1830 1795 1910 1829
rect 1944 1799 1960 1833
rect 1994 1799 2010 1833
rect 1944 1761 2010 1799
rect 2044 1811 2227 1845
rect 2044 1795 2261 1811
rect 2328 1850 2362 1867
rect 2496 1850 2530 1867
rect 2328 1795 2362 1816
rect 2396 1799 2412 1833
rect 2446 1799 2462 1833
rect 2396 1761 2462 1799
rect 2671 1867 2886 1901
rect 3057 1899 3175 1963
rect 3209 1950 3261 1991
rect 3243 1926 3261 1950
rect 3057 1875 3091 1899
rect 2671 1850 2718 1867
rect 2496 1795 2530 1816
rect 2564 1803 2580 1837
rect 2614 1803 2630 1837
rect 2564 1761 2630 1803
rect 2671 1816 2684 1850
rect 2852 1850 2886 1867
rect 2671 1795 2718 1816
rect 2752 1799 2768 1833
rect 2802 1799 2818 1833
rect 2752 1761 2818 1799
rect 2852 1795 2886 1816
rect 2936 1850 3091 1875
rect 3209 1890 3214 1916
rect 3254 1890 3261 1926
rect 2970 1816 3091 1850
rect 2936 1795 3091 1816
rect 3125 1841 3175 1858
rect 3159 1807 3175 1841
rect 3125 1761 3175 1807
rect 3209 1856 3261 1890
rect 3243 1822 3261 1856
rect 3209 1795 3261 1822
rect 3900 2189 3980 2233
rect 4029 2229 4095 2267
rect 4029 2195 4045 2229
rect 4079 2195 4095 2229
rect 4129 2217 4331 2233
rect 3900 2155 3946 2189
rect 4129 2183 4297 2217
rect 4129 2161 4163 2183
rect 4297 2165 4331 2183
rect 4398 2212 4432 2233
rect 4466 2229 4532 2267
rect 4466 2195 4482 2229
rect 4516 2195 4532 2229
rect 4566 2212 4600 2233
rect 3900 2122 3980 2155
rect 4015 2127 4163 2161
rect 4398 2161 4432 2178
rect 4634 2220 4700 2267
rect 4634 2186 4650 2220
rect 4684 2186 4700 2220
rect 4754 2212 4788 2233
rect 4566 2161 4600 2178
rect 3900 1987 3966 2122
rect 4015 2085 4049 2127
rect 4000 2069 4049 2085
rect 4256 2097 4268 2131
rect 4302 2097 4355 2131
rect 4398 2127 4600 2161
rect 4822 2229 4888 2267
rect 4822 2195 4838 2229
rect 4872 2195 4888 2229
rect 4922 2212 4956 2233
rect 4754 2161 4788 2178
rect 4922 2161 4956 2178
rect 4754 2127 4956 2161
rect 5006 2212 5126 2233
rect 5040 2178 5126 2212
rect 5179 2225 5245 2267
rect 5179 2191 5195 2225
rect 5229 2191 5245 2225
rect 5006 2157 5126 2178
rect 5279 2189 5331 2233
rect 5006 2131 5245 2157
rect 5006 2097 5008 2131
rect 5042 2123 5245 2131
rect 5042 2097 5054 2123
rect 4256 2093 4355 2097
rect 4034 2035 4049 2069
rect 4000 2019 4049 2035
rect 4083 2063 4099 2077
rect 4083 2029 4084 2063
rect 4133 2043 4171 2077
rect 4256 2059 4339 2093
rect 4373 2059 4389 2093
rect 4423 2059 4439 2093
rect 4473 2063 4498 2093
rect 4118 2029 4171 2043
rect 4423 2029 4452 2059
rect 4486 2029 4498 2063
rect 4557 2034 4790 2091
rect 5211 2085 5245 2123
rect 5313 2155 5331 2189
rect 5279 2118 5331 2155
rect 3900 1949 3980 1987
rect 3900 1915 3946 1949
rect 3900 1859 3980 1915
rect 4015 1897 4049 2019
rect 4137 1965 4176 1995
rect 4137 1931 4171 1965
rect 4210 1961 4221 1995
rect 4557 1981 4591 2034
rect 4205 1931 4221 1961
rect 4267 1965 4524 1981
rect 4301 1947 4524 1965
rect 4558 1947 4591 1981
rect 4636 1995 4708 1997
rect 4670 1981 4708 1995
rect 4636 1947 4641 1961
rect 4675 1947 4708 1981
rect 4301 1931 4317 1947
rect 4636 1931 4708 1947
rect 4756 1965 4790 2034
rect 4824 2063 4902 2078
rect 5100 2069 5166 2085
rect 5100 2063 5132 2069
rect 4858 2062 4902 2063
rect 4858 2029 4868 2062
rect 4824 2028 4868 2029
rect 4824 2012 4902 2028
rect 4940 2029 4964 2063
rect 4998 2029 5014 2063
rect 5134 2029 5166 2035
rect 4940 1965 4974 2029
rect 5132 2019 5166 2029
rect 5211 2069 5262 2085
rect 5211 2035 5228 2069
rect 5211 2019 5262 2035
rect 4756 1931 4974 1965
rect 5042 1961 5088 1995
rect 5008 1958 5088 1961
rect 5211 1959 5245 2019
rect 5296 1987 5331 2118
rect 4267 1928 4317 1931
rect 4015 1863 4148 1897
rect 4267 1894 4274 1928
rect 4308 1894 4317 1928
rect 5008 1924 5054 1958
rect 5008 1908 5088 1924
rect 4267 1893 4317 1894
rect 3900 1825 3946 1859
rect 4114 1859 4148 1863
rect 4398 1863 4600 1897
rect 4114 1841 4331 1859
rect 3900 1791 3980 1825
rect 4014 1795 4030 1829
rect 4064 1795 4080 1829
rect 1806 1727 1835 1761
rect 1869 1727 1927 1761
rect 1961 1727 2019 1761
rect 2053 1727 2111 1761
rect 2145 1727 2203 1761
rect 2237 1727 2295 1761
rect 2329 1727 2387 1761
rect 2421 1727 2479 1761
rect 2513 1727 2571 1761
rect 2605 1727 2663 1761
rect 2697 1727 2755 1761
rect 2789 1727 2847 1761
rect 2881 1727 2939 1761
rect 2973 1727 3031 1761
rect 3065 1727 3123 1761
rect 3157 1727 3215 1761
rect 3249 1727 3278 1761
rect 4014 1757 4080 1795
rect 4114 1807 4297 1841
rect 4114 1791 4331 1807
rect 4398 1846 4432 1863
rect 4566 1846 4600 1863
rect 4398 1791 4432 1812
rect 4466 1795 4482 1829
rect 4516 1795 4532 1829
rect 4466 1757 4532 1795
rect 4741 1863 4956 1897
rect 5127 1895 5245 1959
rect 5279 1946 5331 1987
rect 5313 1922 5331 1946
rect 5127 1871 5161 1895
rect 4741 1846 4788 1863
rect 4566 1791 4600 1812
rect 4634 1799 4650 1833
rect 4684 1799 4700 1833
rect 4634 1757 4700 1799
rect 4741 1812 4754 1846
rect 4922 1846 4956 1863
rect 4741 1791 4788 1812
rect 4822 1795 4838 1829
rect 4872 1795 4888 1829
rect 4822 1757 4888 1795
rect 4922 1791 4956 1812
rect 5006 1846 5161 1871
rect 5279 1886 5290 1912
rect 5324 1886 5331 1922
rect 5040 1812 5161 1846
rect 5006 1791 5161 1812
rect 5195 1837 5245 1854
rect 5229 1803 5245 1837
rect 5195 1757 5245 1803
rect 5279 1852 5331 1886
rect 5313 1818 5331 1852
rect 5279 1791 5331 1818
rect 5852 2189 5932 2233
rect 5981 2229 6047 2267
rect 5981 2195 5997 2229
rect 6031 2195 6047 2229
rect 6081 2217 6283 2233
rect 5852 2155 5898 2189
rect 6081 2183 6249 2217
rect 6081 2161 6115 2183
rect 6249 2165 6283 2183
rect 6350 2212 6384 2233
rect 6418 2229 6484 2267
rect 6418 2195 6434 2229
rect 6468 2195 6484 2229
rect 6518 2212 6552 2233
rect 5852 2122 5932 2155
rect 5967 2127 6115 2161
rect 6350 2161 6384 2178
rect 6586 2220 6652 2267
rect 6586 2186 6602 2220
rect 6636 2186 6652 2220
rect 6706 2212 6740 2233
rect 6518 2161 6552 2178
rect 5852 1987 5918 2122
rect 5967 2085 6001 2127
rect 5952 2069 6001 2085
rect 6208 2097 6220 2131
rect 6254 2097 6307 2131
rect 6350 2127 6552 2161
rect 6774 2229 6840 2267
rect 6774 2195 6790 2229
rect 6824 2195 6840 2229
rect 6874 2212 6908 2233
rect 6706 2161 6740 2178
rect 6874 2161 6908 2178
rect 6706 2127 6908 2161
rect 6958 2212 7078 2233
rect 6992 2178 7078 2212
rect 7131 2225 7197 2267
rect 7131 2191 7147 2225
rect 7181 2191 7197 2225
rect 6958 2157 7078 2178
rect 7231 2189 7283 2233
rect 6958 2131 7197 2157
rect 6958 2097 6960 2131
rect 6994 2123 7197 2131
rect 6994 2097 7006 2123
rect 6208 2093 6307 2097
rect 5986 2035 6001 2069
rect 5952 2019 6001 2035
rect 6035 2063 6051 2077
rect 6035 2029 6036 2063
rect 6085 2043 6123 2077
rect 6208 2059 6291 2093
rect 6325 2059 6341 2093
rect 6375 2059 6391 2093
rect 6425 2063 6450 2093
rect 6070 2029 6123 2043
rect 6375 2029 6404 2059
rect 6438 2029 6450 2063
rect 6509 2034 6742 2091
rect 7163 2085 7197 2123
rect 7265 2155 7283 2189
rect 7231 2118 7283 2155
rect 5852 1949 5932 1987
rect 5852 1915 5898 1949
rect 5852 1859 5932 1915
rect 5967 1897 6001 2019
rect 6089 1965 6128 1995
rect 6089 1931 6123 1965
rect 6162 1961 6173 1995
rect 6509 1981 6543 2034
rect 6157 1931 6173 1961
rect 6219 1965 6476 1981
rect 6253 1947 6476 1965
rect 6510 1947 6543 1981
rect 6588 1995 6660 1997
rect 6622 1981 6660 1995
rect 6588 1947 6593 1961
rect 6627 1947 6660 1981
rect 6253 1931 6269 1947
rect 6588 1931 6660 1947
rect 6708 1965 6742 2034
rect 6776 2063 6854 2078
rect 7052 2069 7118 2085
rect 7052 2063 7084 2069
rect 6810 2062 6854 2063
rect 6810 2029 6820 2062
rect 6776 2028 6820 2029
rect 6776 2012 6854 2028
rect 6892 2029 6916 2063
rect 6950 2029 6966 2063
rect 7086 2029 7118 2035
rect 6892 1965 6926 2029
rect 7084 2019 7118 2029
rect 7163 2069 7214 2085
rect 7163 2035 7180 2069
rect 7163 2019 7214 2035
rect 6708 1931 6926 1965
rect 6994 1961 7040 1995
rect 6960 1958 7040 1961
rect 7163 1959 7197 2019
rect 7248 1987 7283 2118
rect 6219 1928 6269 1931
rect 5967 1863 6100 1897
rect 6219 1894 6226 1928
rect 6260 1894 6269 1928
rect 6960 1924 7006 1958
rect 6960 1908 7040 1924
rect 6219 1893 6269 1894
rect 5852 1825 5898 1859
rect 6066 1859 6100 1863
rect 6350 1863 6552 1897
rect 6066 1841 6283 1859
rect 5852 1791 5932 1825
rect 5966 1795 5982 1829
rect 6016 1795 6032 1829
rect 5966 1757 6032 1795
rect 6066 1807 6249 1841
rect 6066 1791 6283 1807
rect 6350 1846 6384 1863
rect 6518 1846 6552 1863
rect 6350 1791 6384 1812
rect 6418 1795 6434 1829
rect 6468 1795 6484 1829
rect 6418 1757 6484 1795
rect 6693 1863 6908 1897
rect 7079 1895 7197 1959
rect 7231 1946 7283 1987
rect 7265 1922 7283 1946
rect 7079 1871 7113 1895
rect 6693 1846 6740 1863
rect 6518 1791 6552 1812
rect 6586 1799 6602 1833
rect 6636 1799 6652 1833
rect 6586 1757 6652 1799
rect 6693 1812 6706 1846
rect 6874 1846 6908 1863
rect 6693 1791 6740 1812
rect 6774 1795 6790 1829
rect 6824 1795 6840 1829
rect 6774 1757 6840 1795
rect 6874 1791 6908 1812
rect 6958 1846 7113 1871
rect 7231 1886 7242 1912
rect 7276 1886 7283 1922
rect 6992 1812 7113 1846
rect 6958 1791 7113 1812
rect 7147 1837 7197 1854
rect 7181 1803 7197 1837
rect 7147 1757 7197 1803
rect 7231 1852 7283 1886
rect 7265 1818 7283 1852
rect 7231 1791 7283 1818
rect 7854 2195 7934 2239
rect 7983 2235 8049 2273
rect 7983 2201 7999 2235
rect 8033 2201 8049 2235
rect 8083 2223 8285 2239
rect 7854 2161 7900 2195
rect 8083 2189 8251 2223
rect 8083 2167 8117 2189
rect 8251 2171 8285 2189
rect 8352 2218 8386 2239
rect 8420 2235 8486 2273
rect 8420 2201 8436 2235
rect 8470 2201 8486 2235
rect 8520 2218 8554 2239
rect 7854 2128 7934 2161
rect 7969 2133 8117 2167
rect 8352 2167 8386 2184
rect 8588 2226 8654 2273
rect 8588 2192 8604 2226
rect 8638 2192 8654 2226
rect 8708 2218 8742 2239
rect 8520 2167 8554 2184
rect 7854 1993 7920 2128
rect 7969 2091 8003 2133
rect 7954 2075 8003 2091
rect 8210 2103 8222 2137
rect 8256 2103 8309 2137
rect 8352 2133 8554 2167
rect 8776 2235 8842 2273
rect 8776 2201 8792 2235
rect 8826 2201 8842 2235
rect 8876 2218 8910 2239
rect 8708 2167 8742 2184
rect 8876 2167 8910 2184
rect 8708 2133 8910 2167
rect 8960 2218 9080 2239
rect 8994 2184 9080 2218
rect 9133 2231 9199 2273
rect 9133 2197 9149 2231
rect 9183 2197 9199 2231
rect 8960 2163 9080 2184
rect 9233 2195 9285 2239
rect 8960 2137 9199 2163
rect 8960 2103 8962 2137
rect 8996 2129 9199 2137
rect 8996 2103 9008 2129
rect 8210 2099 8309 2103
rect 7988 2041 8003 2075
rect 7954 2025 8003 2041
rect 8037 2069 8053 2083
rect 8037 2035 8038 2069
rect 8087 2049 8125 2083
rect 8210 2065 8293 2099
rect 8327 2065 8343 2099
rect 8377 2065 8393 2099
rect 8427 2069 8452 2099
rect 8072 2035 8125 2049
rect 8377 2035 8406 2065
rect 8440 2035 8452 2069
rect 8511 2040 8744 2097
rect 9165 2091 9199 2129
rect 9267 2161 9285 2195
rect 9233 2124 9285 2161
rect 7854 1955 7934 1993
rect 7854 1921 7900 1955
rect 7854 1865 7934 1921
rect 7969 1903 8003 2025
rect 8091 1971 8130 2001
rect 8091 1937 8125 1971
rect 8164 1967 8175 2001
rect 8511 1987 8545 2040
rect 8159 1937 8175 1967
rect 8221 1971 8478 1987
rect 8255 1953 8478 1971
rect 8512 1953 8545 1987
rect 8590 2001 8662 2003
rect 8624 1987 8662 2001
rect 8590 1953 8595 1967
rect 8629 1953 8662 1987
rect 8255 1937 8271 1953
rect 8590 1937 8662 1953
rect 8710 1971 8744 2040
rect 8778 2069 8856 2084
rect 9054 2075 9120 2091
rect 9054 2069 9086 2075
rect 8812 2068 8856 2069
rect 8812 2035 8822 2068
rect 8778 2034 8822 2035
rect 8778 2018 8856 2034
rect 8894 2035 8918 2069
rect 8952 2035 8968 2069
rect 9088 2035 9120 2041
rect 8894 1971 8928 2035
rect 9086 2025 9120 2035
rect 9165 2075 9216 2091
rect 9165 2041 9182 2075
rect 9165 2025 9216 2041
rect 8710 1937 8928 1971
rect 8996 1967 9042 2001
rect 8962 1964 9042 1967
rect 9165 1965 9199 2025
rect 9250 1993 9285 2124
rect 8221 1934 8271 1937
rect 7969 1869 8102 1903
rect 8221 1900 8228 1934
rect 8262 1900 8271 1934
rect 8962 1930 9008 1964
rect 8962 1914 9042 1930
rect 8221 1899 8271 1900
rect 7854 1831 7900 1865
rect 8068 1865 8102 1869
rect 8352 1869 8554 1903
rect 8068 1847 8285 1865
rect 7854 1797 7934 1831
rect 7968 1801 7984 1835
rect 8018 1801 8034 1835
rect 7968 1763 8034 1801
rect 8068 1813 8251 1847
rect 8068 1797 8285 1813
rect 8352 1852 8386 1869
rect 8520 1852 8554 1869
rect 8352 1797 8386 1818
rect 8420 1801 8436 1835
rect 8470 1801 8486 1835
rect 8420 1763 8486 1801
rect 8695 1869 8910 1903
rect 9081 1901 9199 1965
rect 9233 1952 9285 1993
rect 9267 1928 9285 1952
rect 9081 1877 9115 1901
rect 8695 1852 8742 1869
rect 8520 1797 8554 1818
rect 8588 1805 8604 1839
rect 8638 1805 8654 1839
rect 8588 1763 8654 1805
rect 8695 1818 8708 1852
rect 8876 1852 8910 1869
rect 8695 1797 8742 1818
rect 8776 1801 8792 1835
rect 8826 1801 8842 1835
rect 8776 1763 8842 1801
rect 8876 1797 8910 1818
rect 8960 1852 9115 1877
rect 9233 1892 9244 1918
rect 9278 1892 9285 1928
rect 8994 1818 9115 1852
rect 8960 1797 9115 1818
rect 9149 1843 9199 1860
rect 9183 1809 9199 1843
rect 9149 1763 9199 1809
rect 9233 1858 9285 1892
rect 9267 1824 9285 1858
rect 9233 1797 9285 1824
rect 9806 2195 9886 2239
rect 9935 2235 10001 2273
rect 9935 2201 9951 2235
rect 9985 2201 10001 2235
rect 10035 2223 10237 2239
rect 9806 2161 9852 2195
rect 10035 2189 10203 2223
rect 10035 2167 10069 2189
rect 10203 2171 10237 2189
rect 10304 2218 10338 2239
rect 10372 2235 10438 2273
rect 10372 2201 10388 2235
rect 10422 2201 10438 2235
rect 10472 2218 10506 2239
rect 9806 2128 9886 2161
rect 9921 2133 10069 2167
rect 10304 2167 10338 2184
rect 10540 2226 10606 2273
rect 10540 2192 10556 2226
rect 10590 2192 10606 2226
rect 10660 2218 10694 2239
rect 10472 2167 10506 2184
rect 9806 1993 9872 2128
rect 9921 2091 9955 2133
rect 9906 2075 9955 2091
rect 10162 2103 10174 2137
rect 10208 2103 10261 2137
rect 10304 2133 10506 2167
rect 10728 2235 10794 2273
rect 10728 2201 10744 2235
rect 10778 2201 10794 2235
rect 10828 2218 10862 2239
rect 10660 2167 10694 2184
rect 10828 2167 10862 2184
rect 10660 2133 10862 2167
rect 10912 2218 11032 2239
rect 10946 2184 11032 2218
rect 11085 2231 11151 2273
rect 11085 2197 11101 2231
rect 11135 2197 11151 2231
rect 10912 2163 11032 2184
rect 11185 2195 11237 2239
rect 10912 2137 11151 2163
rect 10912 2103 10914 2137
rect 10948 2129 11151 2137
rect 10948 2103 10960 2129
rect 10162 2099 10261 2103
rect 9940 2041 9955 2075
rect 9906 2025 9955 2041
rect 9989 2069 10005 2083
rect 9989 2035 9990 2069
rect 10039 2049 10077 2083
rect 10162 2065 10245 2099
rect 10279 2065 10295 2099
rect 10329 2065 10345 2099
rect 10379 2069 10404 2099
rect 10024 2035 10077 2049
rect 10329 2035 10358 2065
rect 10392 2035 10404 2069
rect 10463 2040 10696 2097
rect 11117 2091 11151 2129
rect 11219 2161 11237 2195
rect 11185 2124 11237 2161
rect 9806 1955 9886 1993
rect 9806 1921 9852 1955
rect 9806 1865 9886 1921
rect 9921 1903 9955 2025
rect 10043 1971 10082 2001
rect 10043 1937 10077 1971
rect 10116 1967 10127 2001
rect 10463 1987 10497 2040
rect 10111 1937 10127 1967
rect 10173 1971 10430 1987
rect 10207 1953 10430 1971
rect 10464 1953 10497 1987
rect 10542 2001 10614 2003
rect 10576 1987 10614 2001
rect 10542 1953 10547 1967
rect 10581 1953 10614 1987
rect 10207 1937 10223 1953
rect 10542 1937 10614 1953
rect 10662 1971 10696 2040
rect 10730 2069 10808 2084
rect 11006 2075 11072 2091
rect 11006 2069 11038 2075
rect 10764 2068 10808 2069
rect 10764 2035 10774 2068
rect 10730 2034 10774 2035
rect 10730 2018 10808 2034
rect 10846 2035 10870 2069
rect 10904 2035 10920 2069
rect 11040 2035 11072 2041
rect 10846 1971 10880 2035
rect 11038 2025 11072 2035
rect 11117 2075 11168 2091
rect 11117 2041 11134 2075
rect 11117 2025 11168 2041
rect 10662 1937 10880 1971
rect 10948 1967 10994 2001
rect 10914 1964 10994 1967
rect 11117 1965 11151 2025
rect 11202 1993 11237 2124
rect 10173 1934 10223 1937
rect 9921 1869 10054 1903
rect 10173 1900 10180 1934
rect 10214 1900 10223 1934
rect 10914 1930 10960 1964
rect 10914 1914 10994 1930
rect 10173 1899 10223 1900
rect 9806 1831 9852 1865
rect 10020 1865 10054 1869
rect 10304 1869 10506 1903
rect 10020 1847 10237 1865
rect 9806 1797 9886 1831
rect 9920 1801 9936 1835
rect 9970 1801 9986 1835
rect 9920 1763 9986 1801
rect 10020 1813 10203 1847
rect 10020 1797 10237 1813
rect 10304 1852 10338 1869
rect 10472 1852 10506 1869
rect 10304 1797 10338 1818
rect 10372 1801 10388 1835
rect 10422 1801 10438 1835
rect 10372 1763 10438 1801
rect 10647 1869 10862 1903
rect 11033 1901 11151 1965
rect 11185 1952 11237 1993
rect 11219 1928 11237 1952
rect 11033 1877 11067 1901
rect 10647 1852 10694 1869
rect 10472 1797 10506 1818
rect 10540 1805 10556 1839
rect 10590 1805 10606 1839
rect 10540 1763 10606 1805
rect 10647 1818 10660 1852
rect 10828 1852 10862 1869
rect 10647 1797 10694 1818
rect 10728 1801 10744 1835
rect 10778 1801 10794 1835
rect 10728 1763 10794 1801
rect 10828 1797 10862 1818
rect 10912 1852 11067 1877
rect 11185 1892 11196 1918
rect 11230 1892 11237 1928
rect 10946 1818 11067 1852
rect 10912 1797 11067 1818
rect 11101 1843 11151 1860
rect 11135 1809 11151 1843
rect 11101 1763 11151 1809
rect 11185 1858 11237 1892
rect 11219 1824 11237 1858
rect 11185 1797 11237 1824
rect 11798 2195 11878 2239
rect 11927 2235 11993 2273
rect 11927 2201 11943 2235
rect 11977 2201 11993 2235
rect 12027 2223 12229 2239
rect 11798 2161 11844 2195
rect 12027 2189 12195 2223
rect 12027 2167 12061 2189
rect 12195 2171 12229 2189
rect 12296 2218 12330 2239
rect 12364 2235 12430 2273
rect 12364 2201 12380 2235
rect 12414 2201 12430 2235
rect 12464 2218 12498 2239
rect 11798 2128 11878 2161
rect 11913 2133 12061 2167
rect 12296 2167 12330 2184
rect 12532 2226 12598 2273
rect 12532 2192 12548 2226
rect 12582 2192 12598 2226
rect 12652 2218 12686 2239
rect 12464 2167 12498 2184
rect 11798 1993 11864 2128
rect 11913 2091 11947 2133
rect 11898 2075 11947 2091
rect 12154 2103 12166 2137
rect 12200 2103 12253 2137
rect 12296 2133 12498 2167
rect 12720 2235 12786 2273
rect 12720 2201 12736 2235
rect 12770 2201 12786 2235
rect 12820 2218 12854 2239
rect 12652 2167 12686 2184
rect 12820 2167 12854 2184
rect 12652 2133 12854 2167
rect 12904 2218 13024 2239
rect 12938 2184 13024 2218
rect 13077 2231 13143 2273
rect 13077 2197 13093 2231
rect 13127 2197 13143 2231
rect 12904 2163 13024 2184
rect 13177 2195 13229 2239
rect 12904 2137 13143 2163
rect 12904 2103 12906 2137
rect 12940 2129 13143 2137
rect 12940 2103 12952 2129
rect 12154 2099 12253 2103
rect 11932 2041 11947 2075
rect 11898 2025 11947 2041
rect 11981 2069 11997 2083
rect 11981 2035 11982 2069
rect 12031 2049 12069 2083
rect 12154 2065 12237 2099
rect 12271 2065 12287 2099
rect 12321 2065 12337 2099
rect 12371 2069 12396 2099
rect 12016 2035 12069 2049
rect 12321 2035 12350 2065
rect 12384 2035 12396 2069
rect 12455 2040 12688 2097
rect 13109 2091 13143 2129
rect 13211 2161 13229 2195
rect 13177 2124 13229 2161
rect 11798 1955 11878 1993
rect 11798 1921 11844 1955
rect 11798 1865 11878 1921
rect 11913 1903 11947 2025
rect 12035 1971 12074 2001
rect 12035 1937 12069 1971
rect 12108 1967 12119 2001
rect 12455 1987 12489 2040
rect 12103 1937 12119 1967
rect 12165 1971 12422 1987
rect 12199 1953 12422 1971
rect 12456 1953 12489 1987
rect 12534 2001 12606 2003
rect 12568 1987 12606 2001
rect 12534 1953 12539 1967
rect 12573 1953 12606 1987
rect 12199 1937 12215 1953
rect 12534 1937 12606 1953
rect 12654 1971 12688 2040
rect 12722 2069 12800 2084
rect 12998 2075 13064 2091
rect 12998 2069 13030 2075
rect 12756 2068 12800 2069
rect 12756 2035 12766 2068
rect 12722 2034 12766 2035
rect 12722 2018 12800 2034
rect 12838 2035 12862 2069
rect 12896 2035 12912 2069
rect 13032 2035 13064 2041
rect 12838 1971 12872 2035
rect 13030 2025 13064 2035
rect 13109 2075 13160 2091
rect 13109 2041 13126 2075
rect 13109 2025 13160 2041
rect 12654 1937 12872 1971
rect 12940 1967 12986 2001
rect 12906 1964 12986 1967
rect 13109 1965 13143 2025
rect 13194 1993 13229 2124
rect 12165 1934 12215 1937
rect 11913 1869 12046 1903
rect 12165 1900 12172 1934
rect 12206 1900 12215 1934
rect 12906 1930 12952 1964
rect 12906 1914 12986 1930
rect 12165 1899 12215 1900
rect 11798 1831 11844 1865
rect 12012 1865 12046 1869
rect 12296 1869 12498 1903
rect 12012 1847 12229 1865
rect 11798 1797 11878 1831
rect 11912 1801 11928 1835
rect 11962 1801 11978 1835
rect 11912 1763 11978 1801
rect 12012 1813 12195 1847
rect 12012 1797 12229 1813
rect 12296 1852 12330 1869
rect 12464 1852 12498 1869
rect 12296 1797 12330 1818
rect 12364 1801 12380 1835
rect 12414 1801 12430 1835
rect 12364 1763 12430 1801
rect 12639 1869 12854 1903
rect 13025 1901 13143 1965
rect 13177 1952 13229 1993
rect 13211 1928 13229 1952
rect 13025 1877 13059 1901
rect 12639 1852 12686 1869
rect 12464 1797 12498 1818
rect 12532 1805 12548 1839
rect 12582 1805 12598 1839
rect 12532 1763 12598 1805
rect 12639 1818 12652 1852
rect 12820 1852 12854 1869
rect 12639 1797 12686 1818
rect 12720 1801 12736 1835
rect 12770 1801 12786 1835
rect 12720 1763 12786 1801
rect 12820 1797 12854 1818
rect 12904 1852 13059 1877
rect 13177 1892 13188 1918
rect 13222 1892 13229 1928
rect 12938 1818 13059 1852
rect 12904 1797 13059 1818
rect 13093 1843 13143 1860
rect 13127 1809 13143 1843
rect 13093 1763 13143 1809
rect 13177 1858 13229 1892
rect 13211 1824 13229 1858
rect 13177 1797 13229 1824
rect 13750 2195 13830 2239
rect 13879 2235 13945 2273
rect 13879 2201 13895 2235
rect 13929 2201 13945 2235
rect 13979 2223 14181 2239
rect 13750 2161 13796 2195
rect 13979 2189 14147 2223
rect 13979 2167 14013 2189
rect 14147 2171 14181 2189
rect 14248 2218 14282 2239
rect 14316 2235 14382 2273
rect 14316 2201 14332 2235
rect 14366 2201 14382 2235
rect 14416 2218 14450 2239
rect 13750 2128 13830 2161
rect 13865 2133 14013 2167
rect 14248 2167 14282 2184
rect 14484 2226 14550 2273
rect 14484 2192 14500 2226
rect 14534 2192 14550 2226
rect 14604 2218 14638 2239
rect 14416 2167 14450 2184
rect 13750 1993 13816 2128
rect 13865 2091 13899 2133
rect 13850 2075 13899 2091
rect 14106 2103 14118 2137
rect 14152 2103 14205 2137
rect 14248 2133 14450 2167
rect 14672 2235 14738 2273
rect 14672 2201 14688 2235
rect 14722 2201 14738 2235
rect 14772 2218 14806 2239
rect 14604 2167 14638 2184
rect 14772 2167 14806 2184
rect 14604 2133 14806 2167
rect 14856 2218 14976 2239
rect 14890 2184 14976 2218
rect 15029 2231 15095 2273
rect 15029 2197 15045 2231
rect 15079 2197 15095 2231
rect 14856 2163 14976 2184
rect 15129 2195 15181 2239
rect 14856 2137 15095 2163
rect 14856 2103 14858 2137
rect 14892 2129 15095 2137
rect 14892 2103 14904 2129
rect 14106 2099 14205 2103
rect 13884 2041 13899 2075
rect 13850 2025 13899 2041
rect 13933 2069 13949 2083
rect 13933 2035 13934 2069
rect 13983 2049 14021 2083
rect 14106 2065 14189 2099
rect 14223 2065 14239 2099
rect 14273 2065 14289 2099
rect 14323 2069 14348 2099
rect 13968 2035 14021 2049
rect 14273 2035 14302 2065
rect 14336 2035 14348 2069
rect 14407 2040 14640 2097
rect 15061 2091 15095 2129
rect 15163 2161 15181 2195
rect 15129 2124 15181 2161
rect 13750 1955 13830 1993
rect 13750 1921 13796 1955
rect 13750 1865 13830 1921
rect 13865 1903 13899 2025
rect 13987 1971 14026 2001
rect 13987 1937 14021 1971
rect 14060 1967 14071 2001
rect 14407 1987 14441 2040
rect 14055 1937 14071 1967
rect 14117 1971 14374 1987
rect 14151 1953 14374 1971
rect 14408 1953 14441 1987
rect 14486 2001 14558 2003
rect 14520 1987 14558 2001
rect 14486 1953 14491 1967
rect 14525 1953 14558 1987
rect 14151 1937 14167 1953
rect 14486 1937 14558 1953
rect 14606 1971 14640 2040
rect 14674 2069 14752 2084
rect 14950 2075 15016 2091
rect 14950 2069 14982 2075
rect 14708 2068 14752 2069
rect 14708 2035 14718 2068
rect 14674 2034 14718 2035
rect 14674 2018 14752 2034
rect 14790 2035 14814 2069
rect 14848 2035 14864 2069
rect 14984 2035 15016 2041
rect 14790 1971 14824 2035
rect 14982 2025 15016 2035
rect 15061 2075 15112 2091
rect 15061 2041 15078 2075
rect 15061 2025 15112 2041
rect 14606 1937 14824 1971
rect 14892 1967 14938 2001
rect 14858 1964 14938 1967
rect 15061 1965 15095 2025
rect 15146 1993 15181 2124
rect 14117 1934 14167 1937
rect 13865 1869 13998 1903
rect 14117 1900 14124 1934
rect 14158 1900 14167 1934
rect 14858 1930 14904 1964
rect 14858 1914 14938 1930
rect 14117 1899 14167 1900
rect 13750 1831 13796 1865
rect 13964 1865 13998 1869
rect 14248 1869 14450 1903
rect 13964 1847 14181 1865
rect 13750 1797 13830 1831
rect 13864 1801 13880 1835
rect 13914 1801 13930 1835
rect 13864 1763 13930 1801
rect 13964 1813 14147 1847
rect 13964 1797 14181 1813
rect 14248 1852 14282 1869
rect 14416 1852 14450 1869
rect 14248 1797 14282 1818
rect 14316 1801 14332 1835
rect 14366 1801 14382 1835
rect 14316 1763 14382 1801
rect 14591 1869 14806 1903
rect 14977 1901 15095 1965
rect 15129 1952 15181 1993
rect 15163 1928 15181 1952
rect 14977 1877 15011 1901
rect 14591 1852 14638 1869
rect 14416 1797 14450 1818
rect 14484 1805 14500 1839
rect 14534 1805 14550 1839
rect 14484 1763 14550 1805
rect 14591 1818 14604 1852
rect 14772 1852 14806 1869
rect 14591 1797 14638 1818
rect 14672 1801 14688 1835
rect 14722 1801 14738 1835
rect 14672 1763 14738 1801
rect 14772 1797 14806 1818
rect 14856 1852 15011 1877
rect 15129 1892 15140 1918
rect 15174 1892 15181 1928
rect 14890 1818 15011 1852
rect 14856 1797 15011 1818
rect 15045 1843 15095 1860
rect 15079 1809 15095 1843
rect 15045 1763 15095 1809
rect 15129 1858 15181 1892
rect 15163 1824 15181 1858
rect 15129 1797 15181 1824
rect 15814 2195 15894 2239
rect 15943 2235 16009 2273
rect 15943 2201 15959 2235
rect 15993 2201 16009 2235
rect 16043 2223 16245 2239
rect 15814 2161 15860 2195
rect 16043 2189 16211 2223
rect 16043 2167 16077 2189
rect 16211 2171 16245 2189
rect 16312 2218 16346 2239
rect 16380 2235 16446 2273
rect 16380 2201 16396 2235
rect 16430 2201 16446 2235
rect 16480 2218 16514 2239
rect 15814 2128 15894 2161
rect 15929 2133 16077 2167
rect 16312 2167 16346 2184
rect 16548 2226 16614 2273
rect 16548 2192 16564 2226
rect 16598 2192 16614 2226
rect 16668 2218 16702 2239
rect 16480 2167 16514 2184
rect 15814 1993 15880 2128
rect 15929 2091 15963 2133
rect 15914 2075 15963 2091
rect 16170 2103 16182 2137
rect 16216 2103 16269 2137
rect 16312 2133 16514 2167
rect 16736 2235 16802 2273
rect 16736 2201 16752 2235
rect 16786 2201 16802 2235
rect 16836 2218 16870 2239
rect 16668 2167 16702 2184
rect 16836 2167 16870 2184
rect 16668 2133 16870 2167
rect 16920 2218 17040 2239
rect 16954 2184 17040 2218
rect 17093 2231 17159 2273
rect 17093 2197 17109 2231
rect 17143 2197 17159 2231
rect 16920 2163 17040 2184
rect 17193 2195 17245 2239
rect 16920 2137 17159 2163
rect 16920 2103 16922 2137
rect 16956 2129 17159 2137
rect 16956 2103 16968 2129
rect 16170 2099 16269 2103
rect 15948 2041 15963 2075
rect 15914 2025 15963 2041
rect 15997 2069 16013 2083
rect 15997 2035 15998 2069
rect 16047 2049 16085 2083
rect 16170 2065 16253 2099
rect 16287 2065 16303 2099
rect 16337 2065 16353 2099
rect 16387 2069 16412 2099
rect 16032 2035 16085 2049
rect 16337 2035 16366 2065
rect 16400 2035 16412 2069
rect 16471 2040 16704 2097
rect 17125 2091 17159 2129
rect 17227 2161 17245 2195
rect 17193 2124 17245 2161
rect 15814 1955 15894 1993
rect 15814 1921 15860 1955
rect 15814 1865 15894 1921
rect 15929 1903 15963 2025
rect 16051 1971 16090 2001
rect 16051 1937 16085 1971
rect 16124 1967 16135 2001
rect 16471 1987 16505 2040
rect 16119 1937 16135 1967
rect 16181 1971 16438 1987
rect 16215 1953 16438 1971
rect 16472 1953 16505 1987
rect 16550 2001 16622 2003
rect 16584 1987 16622 2001
rect 16550 1953 16555 1967
rect 16589 1953 16622 1987
rect 16215 1937 16231 1953
rect 16550 1937 16622 1953
rect 16670 1971 16704 2040
rect 16738 2069 16816 2084
rect 17014 2075 17080 2091
rect 17014 2069 17046 2075
rect 16772 2068 16816 2069
rect 16772 2035 16782 2068
rect 16738 2034 16782 2035
rect 16738 2018 16816 2034
rect 16854 2035 16878 2069
rect 16912 2035 16928 2069
rect 17048 2035 17080 2041
rect 16854 1971 16888 2035
rect 17046 2025 17080 2035
rect 17125 2075 17176 2091
rect 17125 2041 17142 2075
rect 17125 2025 17176 2041
rect 16670 1937 16888 1971
rect 16956 1967 17002 2001
rect 16922 1964 17002 1967
rect 17125 1965 17159 2025
rect 17210 1993 17245 2124
rect 16181 1934 16231 1937
rect 15929 1869 16062 1903
rect 16181 1900 16188 1934
rect 16222 1900 16231 1934
rect 16922 1930 16968 1964
rect 16922 1914 17002 1930
rect 16181 1899 16231 1900
rect 15814 1831 15860 1865
rect 16028 1865 16062 1869
rect 16312 1869 16514 1903
rect 16028 1847 16245 1865
rect 15814 1797 15894 1831
rect 15928 1801 15944 1835
rect 15978 1801 15994 1835
rect 15928 1763 15994 1801
rect 16028 1813 16211 1847
rect 16028 1797 16245 1813
rect 16312 1852 16346 1869
rect 16480 1852 16514 1869
rect 16312 1797 16346 1818
rect 16380 1801 16396 1835
rect 16430 1801 16446 1835
rect 16380 1763 16446 1801
rect 16655 1869 16870 1903
rect 17041 1901 17159 1965
rect 17193 1952 17245 1993
rect 17227 1928 17245 1952
rect 17041 1877 17075 1901
rect 16655 1852 16702 1869
rect 16480 1797 16514 1818
rect 16548 1805 16564 1839
rect 16598 1805 16614 1839
rect 16548 1763 16614 1805
rect 16655 1818 16668 1852
rect 16836 1852 16870 1869
rect 16655 1797 16702 1818
rect 16736 1801 16752 1835
rect 16786 1801 16802 1835
rect 16736 1763 16802 1801
rect 16836 1797 16870 1818
rect 16920 1852 17075 1877
rect 17193 1892 17204 1918
rect 17238 1892 17245 1928
rect 16954 1818 17075 1852
rect 16920 1797 17075 1818
rect 17109 1843 17159 1860
rect 17143 1809 17159 1843
rect 17109 1763 17159 1809
rect 17193 1858 17245 1892
rect 17227 1824 17245 1858
rect 17193 1797 17245 1824
rect 3876 1723 3905 1757
rect 3939 1723 3997 1757
rect 4031 1723 4089 1757
rect 4123 1723 4181 1757
rect 4215 1723 4273 1757
rect 4307 1723 4365 1757
rect 4399 1723 4457 1757
rect 4491 1723 4549 1757
rect 4583 1723 4641 1757
rect 4675 1723 4733 1757
rect 4767 1723 4825 1757
rect 4859 1723 4917 1757
rect 4951 1723 5009 1757
rect 5043 1723 5101 1757
rect 5135 1723 5193 1757
rect 5227 1723 5285 1757
rect 5319 1723 5348 1757
rect 5828 1723 5857 1757
rect 5891 1723 5949 1757
rect 5983 1723 6041 1757
rect 6075 1723 6133 1757
rect 6167 1723 6225 1757
rect 6259 1723 6317 1757
rect 6351 1723 6409 1757
rect 6443 1723 6501 1757
rect 6535 1723 6593 1757
rect 6627 1723 6685 1757
rect 6719 1723 6777 1757
rect 6811 1723 6869 1757
rect 6903 1723 6961 1757
rect 6995 1723 7053 1757
rect 7087 1723 7145 1757
rect 7179 1723 7237 1757
rect 7271 1723 7300 1757
rect 7830 1729 7859 1763
rect 7893 1729 7951 1763
rect 7985 1729 8043 1763
rect 8077 1729 8135 1763
rect 8169 1729 8227 1763
rect 8261 1729 8319 1763
rect 8353 1729 8411 1763
rect 8445 1729 8503 1763
rect 8537 1729 8595 1763
rect 8629 1729 8687 1763
rect 8721 1729 8779 1763
rect 8813 1729 8871 1763
rect 8905 1729 8963 1763
rect 8997 1729 9055 1763
rect 9089 1729 9147 1763
rect 9181 1729 9239 1763
rect 9273 1729 9302 1763
rect 9782 1729 9811 1763
rect 9845 1729 9903 1763
rect 9937 1729 9995 1763
rect 10029 1729 10087 1763
rect 10121 1729 10179 1763
rect 10213 1729 10271 1763
rect 10305 1729 10363 1763
rect 10397 1729 10455 1763
rect 10489 1729 10547 1763
rect 10581 1729 10639 1763
rect 10673 1729 10731 1763
rect 10765 1729 10823 1763
rect 10857 1729 10915 1763
rect 10949 1729 11007 1763
rect 11041 1729 11099 1763
rect 11133 1729 11191 1763
rect 11225 1729 11254 1763
rect 11774 1729 11803 1763
rect 11837 1729 11895 1763
rect 11929 1729 11987 1763
rect 12021 1729 12079 1763
rect 12113 1729 12171 1763
rect 12205 1729 12263 1763
rect 12297 1729 12355 1763
rect 12389 1729 12447 1763
rect 12481 1729 12539 1763
rect 12573 1729 12631 1763
rect 12665 1729 12723 1763
rect 12757 1729 12815 1763
rect 12849 1729 12907 1763
rect 12941 1729 12999 1763
rect 13033 1729 13091 1763
rect 13125 1729 13183 1763
rect 13217 1729 13246 1763
rect 13726 1729 13755 1763
rect 13789 1729 13847 1763
rect 13881 1729 13939 1763
rect 13973 1729 14031 1763
rect 14065 1729 14123 1763
rect 14157 1729 14215 1763
rect 14249 1729 14307 1763
rect 14341 1729 14399 1763
rect 14433 1729 14491 1763
rect 14525 1729 14583 1763
rect 14617 1729 14675 1763
rect 14709 1729 14767 1763
rect 14801 1729 14859 1763
rect 14893 1729 14951 1763
rect 14985 1729 15043 1763
rect 15077 1729 15135 1763
rect 15169 1729 15198 1763
rect 15790 1729 15819 1763
rect 15853 1729 15911 1763
rect 15945 1729 16003 1763
rect 16037 1729 16095 1763
rect 16129 1729 16187 1763
rect 16221 1729 16279 1763
rect 16313 1729 16371 1763
rect 16405 1729 16463 1763
rect 16497 1729 16555 1763
rect 16589 1729 16647 1763
rect 16681 1729 16739 1763
rect 16773 1729 16831 1763
rect 16865 1729 16923 1763
rect 16957 1729 17015 1763
rect 17049 1729 17107 1763
rect 17141 1729 17199 1763
rect 17233 1729 17262 1763
<< viali >>
rect 18882 43258 18916 43294
rect 18886 41990 18920 42024
rect 18868 41364 18902 41398
rect 18870 40434 18904 40468
rect 18862 39570 18896 39606
rect 18876 39056 18910 39090
rect 18886 38306 18920 38340
rect 18888 37760 18922 37794
rect 18892 37158 18926 37192
rect 18900 36884 18934 36920
rect 18904 36190 18940 36226
rect 18904 36094 18948 36130
rect 18449 35163 18483 35197
rect 18993 35163 19027 35197
rect 18449 35071 18483 35105
rect 18664 35099 18698 35106
rect 18664 35070 18667 35099
rect 18667 35070 18698 35099
rect 18993 35071 19027 35105
rect 18449 34979 18483 35013
rect 18993 34979 19027 35013
rect 18449 34887 18483 34921
rect 18993 34887 19027 34921
rect 18449 34795 18483 34829
rect 18868 34816 18906 34820
rect 18868 34782 18880 34816
rect 18880 34782 18906 34816
rect 18449 34703 18483 34737
rect 18993 34795 19027 34829
rect 18993 34703 19027 34737
rect 18449 34611 18483 34645
rect 18993 34611 19027 34645
rect 18449 34519 18483 34553
rect 18449 34427 18483 34461
rect 18993 34519 19027 34553
rect 18449 34335 18483 34369
rect 18449 34243 18483 34277
rect 18687 34333 18721 34367
rect 18993 34427 19027 34461
rect 18993 34335 19027 34369
rect 18619 34246 18653 34280
rect 18449 34151 18483 34185
rect 18993 34243 19027 34277
rect 18449 34059 18483 34093
rect 18993 34151 19027 34185
rect 18449 33967 18483 34001
rect 18449 33875 18483 33909
rect 18993 34059 19027 34093
rect 18619 33934 18645 33966
rect 18645 33934 18653 33966
rect 18619 33932 18653 33934
rect 18687 33829 18721 33863
rect 18993 33967 19027 34001
rect 18993 33875 19027 33909
rect 18449 33783 18483 33817
rect 18993 33783 19027 33817
rect 18449 33691 18483 33725
rect 18816 33670 18852 33706
rect 18993 33691 19027 33725
rect 18449 33599 18483 33633
rect 18687 33591 18721 33625
rect 18993 33599 19027 33633
rect 18449 33507 18483 33541
rect 18619 33512 18653 33546
rect 18449 33415 18483 33449
rect 18748 33452 18784 33456
rect 18748 33420 18761 33452
rect 18761 33420 18784 33452
rect 18993 33507 19027 33541
rect 18993 33415 19027 33449
rect 18457 32857 18491 32891
rect 19001 32857 19035 32891
rect 18457 32765 18491 32799
rect 18672 32793 18706 32800
rect 18672 32764 18675 32793
rect 18675 32764 18706 32793
rect 19001 32765 19035 32799
rect 18457 32673 18491 32707
rect 19001 32673 19035 32707
rect 18457 32581 18491 32615
rect 19001 32581 19035 32615
rect 18457 32489 18491 32523
rect 18457 32397 18491 32431
rect 19001 32489 19035 32523
rect 19001 32397 19035 32431
rect 18457 32305 18491 32339
rect 19001 32305 19035 32339
rect 18457 32213 18491 32247
rect 18457 32121 18491 32155
rect 19001 32213 19035 32247
rect 18457 32029 18491 32063
rect 18457 31937 18491 31971
rect 18695 32027 18729 32061
rect 19001 32121 19035 32155
rect 19001 32029 19035 32063
rect 18627 31940 18661 31974
rect 18457 31845 18491 31879
rect 19001 31937 19035 31971
rect 18457 31753 18491 31787
rect 19001 31845 19035 31879
rect 18457 31661 18491 31695
rect 18457 31569 18491 31603
rect 19001 31753 19035 31787
rect 18627 31628 18653 31660
rect 18653 31628 18661 31660
rect 18627 31626 18661 31628
rect 18695 31523 18729 31557
rect 19001 31661 19035 31695
rect 19001 31569 19035 31603
rect 18457 31477 18491 31511
rect 19001 31477 19035 31511
rect 18457 31385 18491 31419
rect 18824 31364 18860 31400
rect 19001 31385 19035 31419
rect 18457 31293 18491 31327
rect 18695 31285 18729 31319
rect 19001 31293 19035 31327
rect 18457 31201 18491 31235
rect 18627 31206 18661 31240
rect 18457 31109 18491 31143
rect 18756 31146 18792 31150
rect 18756 31114 18769 31146
rect 18769 31114 18792 31146
rect 19001 31201 19035 31235
rect 19001 31109 19035 31143
rect 18465 30643 18499 30677
rect 19009 30643 19043 30677
rect 18465 30551 18499 30585
rect 18680 30579 18714 30586
rect 18680 30550 18683 30579
rect 18683 30550 18714 30579
rect 19009 30551 19043 30585
rect 18465 30459 18499 30493
rect 19009 30459 19043 30493
rect 18465 30367 18499 30401
rect 19009 30367 19043 30401
rect 18465 30275 18499 30309
rect 18465 30183 18499 30217
rect 19009 30275 19043 30309
rect 19009 30183 19043 30217
rect 18465 30091 18499 30125
rect 19009 30091 19043 30125
rect 18465 29999 18499 30033
rect 18465 29907 18499 29941
rect 19009 29999 19043 30033
rect 18465 29815 18499 29849
rect 18465 29723 18499 29757
rect 18703 29813 18737 29847
rect 19009 29907 19043 29941
rect 19009 29815 19043 29849
rect 18635 29726 18669 29760
rect 18465 29631 18499 29665
rect 19009 29723 19043 29757
rect 18465 29539 18499 29573
rect 19009 29631 19043 29665
rect 18465 29447 18499 29481
rect 18465 29355 18499 29389
rect 19009 29539 19043 29573
rect 18635 29414 18661 29446
rect 18661 29414 18669 29446
rect 18635 29412 18669 29414
rect 18703 29309 18737 29343
rect 19009 29447 19043 29481
rect 19009 29355 19043 29389
rect 18465 29263 18499 29297
rect 19009 29263 19043 29297
rect 18465 29171 18499 29205
rect 18832 29150 18868 29186
rect 19009 29171 19043 29205
rect 18465 29079 18499 29113
rect 18703 29071 18737 29105
rect 19009 29079 19043 29113
rect 18465 28987 18499 29021
rect 18635 28992 18669 29026
rect 18465 28895 18499 28929
rect 18764 28932 18800 28936
rect 18764 28900 18777 28932
rect 18777 28900 18800 28932
rect 19009 28987 19043 29021
rect 19009 28895 19043 28929
rect 18447 28443 18481 28477
rect 18991 28443 19025 28477
rect 18447 28351 18481 28385
rect 18662 28379 18696 28386
rect 18662 28350 18665 28379
rect 18665 28350 18696 28379
rect 18991 28351 19025 28385
rect 18447 28259 18481 28293
rect 18991 28259 19025 28293
rect 18447 28167 18481 28201
rect 18991 28167 19025 28201
rect 18447 28075 18481 28109
rect 18447 27983 18481 28017
rect 18991 28075 19025 28109
rect 18991 27983 19025 28017
rect 18447 27891 18481 27925
rect 18991 27891 19025 27925
rect 18447 27799 18481 27833
rect 18447 27707 18481 27741
rect 18991 27799 19025 27833
rect 18447 27615 18481 27649
rect 18447 27523 18481 27557
rect 18685 27613 18719 27647
rect 18991 27707 19025 27741
rect 18991 27615 19025 27649
rect 18617 27526 18651 27560
rect 18447 27431 18481 27465
rect 18991 27523 19025 27557
rect 18447 27339 18481 27373
rect 18991 27431 19025 27465
rect 18447 27247 18481 27281
rect 18447 27155 18481 27189
rect 18991 27339 19025 27373
rect 18617 27214 18643 27246
rect 18643 27214 18651 27246
rect 18617 27212 18651 27214
rect 18685 27109 18719 27143
rect 18991 27247 19025 27281
rect 18991 27155 19025 27189
rect 18447 27063 18481 27097
rect 18991 27063 19025 27097
rect 18447 26971 18481 27005
rect 18814 26950 18850 26986
rect 18991 26971 19025 27005
rect 18447 26879 18481 26913
rect 18685 26871 18719 26905
rect 18991 26879 19025 26913
rect 18447 26787 18481 26821
rect 18617 26792 18651 26826
rect 18447 26695 18481 26729
rect 18746 26732 18782 26736
rect 18746 26700 18759 26732
rect 18759 26700 18782 26732
rect 18991 26787 19025 26821
rect 18991 26695 19025 26729
rect 18455 26229 18489 26263
rect 18999 26229 19033 26263
rect 18455 26137 18489 26171
rect 18670 26165 18704 26172
rect 18670 26136 18673 26165
rect 18673 26136 18704 26165
rect 18999 26137 19033 26171
rect 18455 26045 18489 26079
rect 18999 26045 19033 26079
rect 18455 25953 18489 25987
rect 18999 25953 19033 25987
rect 18455 25861 18489 25895
rect 18455 25769 18489 25803
rect 18999 25861 19033 25895
rect 18999 25769 19033 25803
rect 18455 25677 18489 25711
rect 18999 25677 19033 25711
rect 18455 25585 18489 25619
rect 18455 25493 18489 25527
rect 18999 25585 19033 25619
rect 18455 25401 18489 25435
rect 18455 25309 18489 25343
rect 18693 25399 18727 25433
rect 18999 25493 19033 25527
rect 18999 25401 19033 25435
rect 18625 25312 18659 25346
rect 18455 25217 18489 25251
rect 18999 25309 19033 25343
rect 18455 25125 18489 25159
rect 18999 25217 19033 25251
rect 18455 25033 18489 25067
rect 18455 24941 18489 24975
rect 18999 25125 19033 25159
rect 18625 25000 18651 25032
rect 18651 25000 18659 25032
rect 18625 24998 18659 25000
rect 18693 24895 18727 24929
rect 18999 25033 19033 25067
rect 18999 24941 19033 24975
rect 18455 24849 18489 24883
rect 18999 24849 19033 24883
rect 18455 24757 18489 24791
rect 18822 24736 18858 24772
rect 18999 24757 19033 24791
rect 18455 24665 18489 24699
rect 18693 24657 18727 24691
rect 18999 24665 19033 24699
rect 18455 24573 18489 24607
rect 18625 24578 18659 24612
rect 18455 24481 18489 24515
rect 18754 24518 18790 24522
rect 18754 24486 18767 24518
rect 18767 24486 18790 24518
rect 18999 24573 19033 24607
rect 18999 24481 19033 24515
rect 7575 23371 7609 23405
rect 7667 23371 7701 23405
rect 7759 23371 7793 23405
rect 7851 23371 7885 23405
rect 7943 23371 7977 23405
rect 8035 23371 8069 23405
rect 8127 23371 8161 23405
rect 8219 23371 8253 23405
rect 8311 23371 8345 23405
rect 8403 23371 8437 23405
rect 8495 23371 8529 23405
rect 8587 23371 8621 23405
rect 8679 23371 8713 23405
rect 8771 23371 8805 23405
rect 8863 23371 8897 23405
rect 8955 23371 8989 23405
rect 9047 23371 9081 23405
rect 9139 23371 9173 23405
rect 9231 23371 9265 23405
rect 9323 23371 9357 23405
rect 9789 23379 9823 23413
rect 9881 23379 9915 23413
rect 9973 23379 10007 23413
rect 10065 23379 10099 23413
rect 10157 23379 10191 23413
rect 10249 23379 10283 23413
rect 10341 23379 10375 23413
rect 10433 23379 10467 23413
rect 10525 23379 10559 23413
rect 10617 23379 10651 23413
rect 10709 23379 10743 23413
rect 10801 23379 10835 23413
rect 10893 23379 10927 23413
rect 10985 23379 11019 23413
rect 11077 23379 11111 23413
rect 11169 23379 11203 23413
rect 11261 23379 11295 23413
rect 11353 23379 11387 23413
rect 11445 23379 11479 23413
rect 11537 23379 11571 23413
rect 7672 23201 7706 23235
rect 7580 23093 7616 23106
rect 7580 23070 7612 23093
rect 7612 23070 7616 23093
rect 7751 23133 7785 23167
rect 7830 23002 7866 23038
rect 8092 23209 8126 23235
rect 8092 23201 8094 23209
rect 8094 23201 8126 23209
rect 7989 23133 8023 23167
rect 8406 23201 8440 23235
rect 8493 23133 8527 23167
rect 9230 23187 9266 23190
rect 9230 23156 9259 23187
rect 9259 23156 9266 23187
rect 9886 23209 9920 23243
rect 9794 23101 9830 23114
rect 9794 23078 9826 23101
rect 9826 23078 9830 23101
rect 9965 23141 9999 23175
rect 10044 23010 10080 23046
rect 10306 23217 10340 23243
rect 10306 23209 10308 23217
rect 10308 23209 10340 23217
rect 10203 23141 10237 23175
rect 10620 23209 10654 23243
rect 10707 23141 10741 23175
rect 11444 23195 11480 23198
rect 11444 23164 11473 23195
rect 11473 23164 11480 23195
rect 11989 23361 12023 23395
rect 12081 23361 12115 23395
rect 12173 23361 12207 23395
rect 12265 23361 12299 23395
rect 12357 23361 12391 23395
rect 12449 23361 12483 23395
rect 12541 23361 12575 23395
rect 12633 23361 12667 23395
rect 12725 23361 12759 23395
rect 12817 23361 12851 23395
rect 12909 23361 12943 23395
rect 13001 23361 13035 23395
rect 13093 23361 13127 23395
rect 13185 23361 13219 23395
rect 13277 23361 13311 23395
rect 13369 23361 13403 23395
rect 13461 23361 13495 23395
rect 13553 23361 13587 23395
rect 13645 23361 13679 23395
rect 13737 23361 13771 23395
rect 14203 23369 14237 23403
rect 14295 23369 14329 23403
rect 14387 23369 14421 23403
rect 14479 23369 14513 23403
rect 14571 23369 14605 23403
rect 14663 23369 14697 23403
rect 14755 23369 14789 23403
rect 14847 23369 14881 23403
rect 14939 23369 14973 23403
rect 15031 23369 15065 23403
rect 15123 23369 15157 23403
rect 15215 23369 15249 23403
rect 15307 23369 15341 23403
rect 15399 23369 15433 23403
rect 15491 23369 15525 23403
rect 15583 23369 15617 23403
rect 15675 23369 15709 23403
rect 15767 23369 15801 23403
rect 15859 23369 15893 23403
rect 15951 23369 15985 23403
rect 16509 23377 16543 23411
rect 16601 23377 16635 23411
rect 16693 23377 16727 23411
rect 16785 23377 16819 23411
rect 16877 23377 16911 23411
rect 16969 23377 17003 23411
rect 17061 23377 17095 23411
rect 17153 23377 17187 23411
rect 17245 23377 17279 23411
rect 17337 23377 17371 23411
rect 17429 23377 17463 23411
rect 17521 23377 17555 23411
rect 17613 23377 17647 23411
rect 17705 23377 17739 23411
rect 17797 23377 17831 23411
rect 17889 23377 17923 23411
rect 17981 23377 18015 23411
rect 18073 23377 18107 23411
rect 18165 23377 18199 23411
rect 18257 23377 18291 23411
rect 12086 23191 12120 23225
rect 11994 23083 12030 23096
rect 11994 23060 12026 23083
rect 12026 23060 12030 23083
rect 12165 23123 12199 23157
rect 12244 22992 12280 23028
rect 12506 23199 12540 23225
rect 12506 23191 12508 23199
rect 12508 23191 12540 23199
rect 12403 23123 12437 23157
rect 7575 22827 7609 22861
rect 7667 22827 7701 22861
rect 7759 22827 7793 22861
rect 7851 22827 7885 22861
rect 7943 22827 7977 22861
rect 8035 22827 8069 22861
rect 8127 22827 8161 22861
rect 8219 22827 8253 22861
rect 8311 22827 8345 22861
rect 8403 22827 8437 22861
rect 8495 22827 8529 22861
rect 8587 22827 8621 22861
rect 8679 22827 8713 22861
rect 8771 22827 8805 22861
rect 8863 22827 8897 22861
rect 8955 22827 8989 22861
rect 9047 22827 9081 22861
rect 9139 22827 9173 22861
rect 9231 22827 9265 22861
rect 9323 22827 9357 22861
rect 9789 22835 9823 22869
rect 9881 22835 9915 22869
rect 9973 22835 10007 22869
rect 10065 22835 10099 22869
rect 10157 22835 10191 22869
rect 10249 22835 10283 22869
rect 10341 22835 10375 22869
rect 10433 22835 10467 22869
rect 10525 22835 10559 22869
rect 10617 22835 10651 22869
rect 10709 22835 10743 22869
rect 10801 22835 10835 22869
rect 10893 22835 10927 22869
rect 10985 22835 11019 22869
rect 11077 22835 11111 22869
rect 11169 22835 11203 22869
rect 11261 22835 11295 22869
rect 11353 22835 11387 22869
rect 11445 22835 11479 22869
rect 11537 22835 11571 22869
rect 12820 23191 12854 23225
rect 12907 23123 12941 23157
rect 13644 23177 13680 23180
rect 13644 23146 13673 23177
rect 13673 23146 13680 23177
rect 14300 23199 14334 23233
rect 14208 23091 14244 23104
rect 14208 23068 14240 23091
rect 14240 23068 14244 23091
rect 14379 23131 14413 23165
rect 14458 23000 14494 23036
rect 14720 23207 14754 23233
rect 14720 23199 14722 23207
rect 14722 23199 14754 23207
rect 14617 23131 14651 23165
rect 15034 23199 15068 23233
rect 15121 23131 15155 23165
rect 15858 23185 15894 23188
rect 15858 23154 15887 23185
rect 15887 23154 15894 23185
rect 16606 23207 16640 23241
rect 16514 23099 16550 23112
rect 16514 23076 16546 23099
rect 16546 23076 16550 23099
rect 16685 23139 16719 23173
rect 16764 23008 16800 23044
rect 17026 23215 17060 23241
rect 17026 23207 17028 23215
rect 17028 23207 17060 23215
rect 16923 23139 16957 23173
rect 17340 23207 17374 23241
rect 17427 23139 17461 23173
rect 18164 23193 18200 23196
rect 18164 23162 18193 23193
rect 18193 23162 18200 23193
rect 11989 22817 12023 22851
rect 12081 22817 12115 22851
rect 12173 22817 12207 22851
rect 12265 22817 12299 22851
rect 12357 22817 12391 22851
rect 12449 22817 12483 22851
rect 12541 22817 12575 22851
rect 12633 22817 12667 22851
rect 12725 22817 12759 22851
rect 12817 22817 12851 22851
rect 12909 22817 12943 22851
rect 13001 22817 13035 22851
rect 13093 22817 13127 22851
rect 13185 22817 13219 22851
rect 13277 22817 13311 22851
rect 13369 22817 13403 22851
rect 13461 22817 13495 22851
rect 13553 22817 13587 22851
rect 13645 22817 13679 22851
rect 13737 22817 13771 22851
rect 14203 22825 14237 22859
rect 14295 22825 14329 22859
rect 14387 22825 14421 22859
rect 14479 22825 14513 22859
rect 14571 22825 14605 22859
rect 14663 22825 14697 22859
rect 14755 22825 14789 22859
rect 14847 22825 14881 22859
rect 14939 22825 14973 22859
rect 15031 22825 15065 22859
rect 15123 22825 15157 22859
rect 15215 22825 15249 22859
rect 15307 22825 15341 22859
rect 15399 22825 15433 22859
rect 15491 22825 15525 22859
rect 15583 22825 15617 22859
rect 15675 22825 15709 22859
rect 15767 22825 15801 22859
rect 15859 22825 15893 22859
rect 15951 22825 15985 22859
rect 16509 22833 16543 22867
rect 16601 22833 16635 22867
rect 16693 22833 16727 22867
rect 16785 22833 16819 22867
rect 16877 22833 16911 22867
rect 16969 22833 17003 22867
rect 17061 22833 17095 22867
rect 17153 22833 17187 22867
rect 17245 22833 17279 22867
rect 17337 22833 17371 22867
rect 17429 22833 17463 22867
rect 17521 22833 17555 22867
rect 17613 22833 17647 22867
rect 17705 22833 17739 22867
rect 17797 22833 17831 22867
rect 17889 22833 17923 22867
rect 17981 22833 18015 22867
rect 18073 22833 18107 22867
rect 18165 22833 18199 22867
rect 18257 22833 18291 22867
rect 16296 17667 16330 17701
rect 16374 17667 16408 17701
rect 16466 17667 16500 17701
rect 16558 17667 16592 17701
rect 17162 17669 17196 17703
rect 17248 17669 17282 17703
rect 17340 17669 17374 17703
rect 17432 17669 17466 17703
rect 15510 17629 15544 17663
rect 15596 17629 15630 17663
rect 15688 17629 15722 17663
rect 15780 17629 15814 17663
rect 9496 17532 9532 17568
rect 9596 17536 9632 17572
rect 17940 17659 17974 17693
rect 18016 17659 18050 17693
rect 18108 17659 18142 17693
rect 18200 17659 18234 17693
rect 19056 17661 19090 17695
rect 19138 17661 19172 17695
rect 19230 17661 19264 17695
rect 19322 17661 19356 17695
rect 19922 17663 19956 17697
rect 20012 17663 20046 17697
rect 20104 17663 20138 17697
rect 20196 17663 20230 17697
rect 15635 17402 15669 17436
rect 16413 17434 16449 17468
rect 15725 17397 15729 17428
rect 15729 17397 15763 17428
rect 15725 17394 15763 17397
rect 16517 17435 16541 17464
rect 16541 17435 16551 17464
rect 16517 17430 16551 17435
rect 17287 17442 17321 17476
rect 17377 17437 17381 17468
rect 17381 17437 17415 17468
rect 17377 17434 17415 17437
rect 18059 17438 18097 17472
rect 20692 17653 20726 17687
rect 20780 17653 20814 17687
rect 20872 17653 20906 17687
rect 20964 17653 20998 17687
rect 16296 17123 16330 17157
rect 16374 17123 16408 17157
rect 16466 17123 16500 17157
rect 16558 17123 16592 17157
rect 17162 17125 17196 17159
rect 17248 17125 17282 17159
rect 17340 17125 17374 17159
rect 17432 17125 17466 17159
rect 18147 17427 18149 17460
rect 18149 17427 18183 17460
rect 18147 17426 18183 17427
rect 19177 17428 19213 17462
rect 19281 17429 19305 17458
rect 19305 17429 19315 17458
rect 19281 17424 19315 17429
rect 20051 17436 20085 17470
rect 21394 17651 21428 17685
rect 21486 17651 21520 17685
rect 21578 17651 21612 17685
rect 21670 17651 21704 17685
rect 22178 17653 22212 17687
rect 22268 17653 22302 17687
rect 22360 17653 22394 17687
rect 22452 17653 22486 17687
rect 20141 17431 20145 17462
rect 20145 17431 20179 17462
rect 20141 17428 20179 17431
rect 20823 17432 20861 17466
rect 15510 17085 15544 17119
rect 15596 17085 15630 17119
rect 15688 17085 15722 17119
rect 15780 17085 15814 17119
rect 17940 17115 17974 17149
rect 18016 17115 18050 17149
rect 18108 17115 18142 17149
rect 18200 17115 18234 17149
rect 19056 17117 19090 17151
rect 19138 17117 19172 17151
rect 19230 17117 19264 17151
rect 19322 17117 19356 17151
rect 19922 17119 19956 17153
rect 20012 17119 20046 17153
rect 20104 17119 20138 17153
rect 20196 17119 20230 17153
rect 20911 17421 20913 17454
rect 20913 17421 20947 17454
rect 20911 17420 20947 17421
rect 23036 17643 23070 17677
rect 23128 17643 23162 17677
rect 23220 17643 23254 17677
rect 23310 17643 23344 17677
rect 21433 17418 21469 17452
rect 21537 17419 21561 17448
rect 21561 17419 21571 17448
rect 21537 17414 21571 17419
rect 22307 17426 22341 17460
rect 20692 17109 20726 17143
rect 20780 17109 20814 17143
rect 20872 17109 20906 17143
rect 20964 17109 20998 17143
rect 22397 17421 22401 17452
rect 22401 17421 22435 17452
rect 22397 17418 22435 17421
rect 23079 17422 23117 17456
rect 23167 17411 23169 17444
rect 23169 17411 23203 17444
rect 23167 17410 23203 17411
rect 21394 17107 21428 17141
rect 21486 17107 21520 17141
rect 21578 17107 21612 17141
rect 21670 17107 21704 17141
rect 22178 17109 22212 17143
rect 22268 17109 22302 17143
rect 22360 17109 22394 17143
rect 22452 17109 22486 17143
rect 23036 17099 23070 17133
rect 23128 17099 23162 17133
rect 23220 17099 23254 17133
rect 23310 17099 23344 17133
rect 9363 16573 9397 16607
rect 9455 16573 9489 16607
rect 9547 16573 9581 16607
rect 9639 16573 9673 16607
rect 9731 16573 9765 16607
rect 9823 16573 9857 16607
rect 9915 16573 9949 16607
rect 9910 16387 9944 16394
rect 9910 16356 9935 16387
rect 9935 16356 9944 16387
rect 16416 16366 16452 16400
rect 16502 16354 16540 16388
rect 17184 16358 17222 16392
rect 9420 16295 9454 16296
rect 9420 16262 9453 16295
rect 9453 16262 9454 16295
rect 9540 16295 9574 16298
rect 9540 16264 9570 16295
rect 9570 16264 9574 16295
rect 17278 16350 17312 16384
rect 18048 16362 18082 16396
rect 18150 16358 18186 16392
rect 18672 16356 18708 16390
rect 18758 16344 18796 16378
rect 19440 16348 19478 16382
rect 19534 16340 19568 16374
rect 20304 16352 20338 16386
rect 20406 16348 20442 16382
rect 21436 16350 21472 16384
rect 21522 16338 21560 16372
rect 22204 16342 22242 16376
rect 22298 16334 22332 16368
rect 23068 16346 23102 16380
rect 23170 16342 23206 16376
rect 9363 16029 9397 16063
rect 9455 16029 9489 16063
rect 9547 16029 9581 16063
rect 9639 16029 9673 16063
rect 9731 16029 9765 16063
rect 9823 16029 9857 16063
rect 9915 16029 9949 16063
rect 9461 15829 9495 15863
rect 9553 15829 9587 15863
rect 9645 15829 9679 15863
rect 9737 15829 9771 15863
rect 9829 15829 9863 15863
rect 11503 15719 11537 15753
rect 11595 15719 11629 15753
rect 11687 15719 11721 15753
rect 11779 15719 11813 15753
rect 11871 15719 11905 15753
rect 11963 15719 11997 15753
rect 12055 15719 12089 15753
rect 9454 15534 9496 15574
rect 9644 15551 9686 15564
rect 9644 15524 9647 15551
rect 9647 15524 9681 15551
rect 9681 15524 9686 15551
rect 9836 15460 9872 15494
rect 11498 15368 11534 15404
rect 9461 15285 9495 15319
rect 9553 15285 9587 15319
rect 9645 15285 9679 15319
rect 9737 15285 9771 15319
rect 9829 15285 9863 15319
rect 11670 15407 11685 15438
rect 11685 15407 11704 15438
rect 11670 15402 11704 15407
rect 11768 15280 11802 15314
rect 11864 15348 11898 15384
rect 12056 15402 12090 15436
rect 10645 15219 10679 15253
rect 10737 15219 10771 15253
rect 10829 15219 10863 15253
rect 10921 15219 10955 15253
rect 11013 15219 11047 15253
rect 9373 15009 9407 15043
rect 9465 15009 9499 15043
rect 9557 15009 9591 15043
rect 9649 15009 9683 15043
rect 9741 15009 9775 15043
rect 9833 15009 9867 15043
rect 9925 15009 9959 15043
rect 11503 15175 11537 15209
rect 11595 15175 11629 15209
rect 11687 15175 11721 15209
rect 11779 15175 11813 15209
rect 11871 15175 11905 15209
rect 11963 15175 11997 15209
rect 12055 15175 12089 15209
rect 11010 15143 11017 15152
rect 11017 15143 11050 15152
rect 11010 15116 11050 15143
rect 9922 14925 9945 14934
rect 9945 14925 9956 14934
rect 9922 14900 9956 14925
rect 10690 14941 10724 14942
rect 10690 14908 10724 14941
rect 10830 14941 10866 14942
rect 10830 14908 10831 14941
rect 10831 14908 10865 14941
rect 10865 14908 10866 14941
rect 9430 14731 9464 14732
rect 9430 14698 9463 14731
rect 9463 14698 9464 14731
rect 9550 14731 9584 14734
rect 9550 14700 9580 14731
rect 9580 14700 9584 14731
rect 10645 14675 10679 14709
rect 10737 14675 10771 14709
rect 10829 14675 10863 14709
rect 10921 14675 10955 14709
rect 11013 14675 11047 14709
rect 24150 14616 24186 14650
rect 23530 14546 23568 14580
rect 23672 14528 23708 14562
rect 24556 14554 24592 14588
rect 24456 14518 24492 14552
rect 24712 14528 24746 14562
rect 25356 14560 25390 14594
rect 9373 14465 9407 14499
rect 9465 14465 9499 14499
rect 9557 14465 9591 14499
rect 9649 14465 9683 14499
rect 9741 14465 9775 14499
rect 9833 14465 9867 14499
rect 9925 14465 9959 14499
rect 9471 14265 9505 14299
rect 9563 14265 9597 14299
rect 9655 14265 9689 14299
rect 9747 14265 9781 14299
rect 9839 14265 9873 14299
rect 10719 14253 10753 14287
rect 10811 14253 10845 14287
rect 10903 14253 10937 14287
rect 10995 14253 11029 14287
rect 11087 14253 11121 14287
rect 11179 14253 11213 14287
rect 11271 14253 11305 14287
rect 8212 14036 8254 14076
rect 9464 13970 9506 14010
rect 9654 13987 9696 14000
rect 9654 13960 9657 13987
rect 9657 13960 9691 13987
rect 9691 13960 9696 13987
rect 7752 13904 7792 13938
rect 9844 13854 9880 13888
rect 12617 14237 12651 14271
rect 12709 14237 12743 14271
rect 12801 14237 12835 14271
rect 12893 14237 12927 14271
rect 12985 14237 13019 14271
rect 13077 14237 13111 14271
rect 12762 14136 12798 14170
rect 10716 13975 10750 13980
rect 10716 13946 10721 13975
rect 10721 13946 10750 13975
rect 10886 13850 10920 13884
rect 10984 13890 11018 13924
rect 11078 13941 11103 13974
rect 11103 13941 11114 13974
rect 11078 13936 11114 13941
rect 13078 14062 13103 14080
rect 13103 14062 13120 14080
rect 11260 13853 11265 13856
rect 11265 13853 11298 13856
rect 11689 13879 11723 13913
rect 11781 13879 11815 13913
rect 11873 13879 11907 13913
rect 11965 13879 11999 13913
rect 12057 13879 12091 13913
rect 12618 13925 12623 13942
rect 12623 13925 12657 13942
rect 12657 13925 12658 13942
rect 12618 13908 12658 13925
rect 13078 14040 13120 14062
rect 12746 13959 12796 13964
rect 12746 13925 12749 13959
rect 12749 13925 12783 13959
rect 12783 13925 12796 13959
rect 12746 13922 12796 13925
rect 12918 13959 12956 13960
rect 12918 13925 12925 13959
rect 12925 13925 12956 13959
rect 12918 13924 12956 13925
rect 11260 13819 11298 13853
rect 11260 13818 11265 13819
rect 11265 13818 11298 13819
rect 9471 13721 9505 13755
rect 9563 13721 9597 13755
rect 9655 13721 9689 13755
rect 9747 13721 9781 13755
rect 9839 13721 9873 13755
rect 10719 13709 10753 13743
rect 10811 13709 10845 13743
rect 10903 13709 10937 13743
rect 10995 13709 11029 13743
rect 11087 13709 11121 13743
rect 11179 13709 11213 13743
rect 11271 13709 11305 13743
rect 12028 13735 12039 13768
rect 12039 13735 12062 13768
rect 12028 13734 12062 13735
rect 11700 13524 11734 13558
rect 11878 13601 11912 13608
rect 11878 13574 11896 13601
rect 11896 13574 11912 13601
rect 12617 13693 12651 13727
rect 12709 13693 12743 13727
rect 12801 13693 12835 13727
rect 12893 13693 12927 13727
rect 12985 13693 13019 13727
rect 13077 13693 13111 13727
rect 10843 13411 10877 13445
rect 10935 13411 10969 13445
rect 11027 13411 11061 13445
rect 11119 13411 11153 13445
rect 11211 13411 11245 13445
rect 9365 13341 9399 13375
rect 9457 13341 9491 13375
rect 9549 13341 9583 13375
rect 9641 13341 9675 13375
rect 9733 13341 9767 13375
rect 9825 13341 9859 13375
rect 9917 13341 9951 13375
rect 11012 13326 11021 13338
rect 11021 13326 11048 13338
rect 11012 13302 11048 13326
rect 11689 13335 11723 13369
rect 11781 13335 11815 13369
rect 11873 13335 11907 13369
rect 11965 13335 11999 13369
rect 12057 13335 12091 13369
rect 9914 13223 9948 13224
rect 9914 13190 9937 13223
rect 9937 13190 9948 13223
rect 11208 13253 11239 13282
rect 11239 13253 11246 13282
rect 11208 13244 11246 13253
rect 9422 13063 9456 13064
rect 9422 13030 9455 13063
rect 9455 13030 9456 13063
rect 9542 13063 9576 13066
rect 9542 13032 9572 13063
rect 9572 13032 9576 13063
rect 10860 13053 10883 13064
rect 10883 13053 10894 13064
rect 10860 13030 10894 13053
rect 11062 13036 11098 13070
rect 10843 12867 10877 12901
rect 10935 12867 10969 12901
rect 11027 12867 11061 12901
rect 11119 12867 11153 12901
rect 11211 12867 11245 12901
rect 9365 12797 9399 12831
rect 9457 12797 9491 12831
rect 9549 12797 9583 12831
rect 9641 12797 9675 12831
rect 9733 12797 9767 12831
rect 9825 12797 9859 12831
rect 9917 12797 9951 12831
rect 9463 12597 9497 12631
rect 9555 12597 9589 12631
rect 9647 12597 9681 12631
rect 9739 12597 9773 12631
rect 9831 12597 9865 12631
rect 9456 12302 9498 12342
rect 10839 12391 10873 12425
rect 10931 12391 10965 12425
rect 11023 12391 11057 12425
rect 11115 12391 11149 12425
rect 11207 12391 11241 12425
rect 9836 12340 9872 12374
rect 9646 12319 9688 12332
rect 9646 12292 9649 12319
rect 9649 12292 9683 12319
rect 9683 12292 9688 12319
rect 11212 12166 11246 12200
rect 9463 12053 9497 12087
rect 9555 12053 9589 12087
rect 9647 12053 9681 12087
rect 9739 12053 9773 12087
rect 9831 12053 9865 12087
rect 10884 12113 10920 12116
rect 10884 12082 10918 12113
rect 10918 12082 10920 12113
rect 11024 12113 11060 12114
rect 11024 12080 11025 12113
rect 11025 12080 11059 12113
rect 11059 12080 11060 12113
rect 10839 11847 10873 11881
rect 10931 11847 10965 11881
rect 11023 11847 11057 11881
rect 11115 11847 11149 11881
rect 11207 11847 11241 11881
rect 9375 11777 9409 11811
rect 9467 11777 9501 11811
rect 9559 11777 9593 11811
rect 9651 11777 9685 11811
rect 9743 11777 9777 11811
rect 9835 11777 9869 11811
rect 9927 11777 9961 11811
rect 9914 11659 9950 11660
rect 9914 11626 9947 11659
rect 9947 11626 9950 11659
rect 9432 11499 9466 11500
rect 9432 11466 9465 11499
rect 9465 11466 9466 11499
rect 9552 11499 9586 11502
rect 9552 11468 9582 11499
rect 9582 11468 9586 11499
rect 9375 11233 9409 11267
rect 9467 11233 9501 11267
rect 9559 11233 9593 11267
rect 9651 11233 9685 11267
rect 9743 11233 9777 11267
rect 9835 11233 9869 11267
rect 9927 11233 9961 11267
rect 9473 11033 9507 11067
rect 9565 11033 9599 11067
rect 9657 11033 9691 11067
rect 9749 11033 9783 11067
rect 9841 11033 9875 11067
rect 9466 10738 9508 10778
rect 4982 10694 5016 10730
rect 9656 10755 9698 10768
rect 9656 10728 9659 10755
rect 9659 10728 9693 10755
rect 9693 10728 9698 10755
rect 9848 10698 9882 10734
rect 9473 10489 9507 10523
rect 9565 10489 9599 10523
rect 9657 10489 9691 10523
rect 9749 10489 9783 10523
rect 9841 10489 9875 10523
rect 6141 6583 6175 6617
rect 6233 6583 6267 6617
rect 6325 6583 6359 6617
rect 6178 6348 6212 6382
rect 6274 6351 6308 6384
rect 6274 6350 6308 6351
rect 6141 6039 6175 6073
rect 6233 6039 6267 6073
rect 6325 6039 6359 6073
rect 10047 5951 10081 5985
rect 10139 5951 10173 5985
rect 10231 5951 10265 5985
rect 10323 5951 10357 5985
rect 10415 5951 10449 5985
rect 10507 5951 10541 5985
rect 10599 5951 10633 5985
rect 10691 5951 10725 5985
rect 10783 5951 10817 5985
rect 10875 5951 10909 5985
rect 10967 5951 11001 5985
rect 11059 5951 11093 5985
rect 11151 5951 11185 5985
rect 11243 5951 11277 5985
rect 11335 5951 11369 5985
rect 11427 5951 11461 5985
rect 10410 5781 10444 5815
rect 12109 5939 12143 5973
rect 12201 5939 12235 5973
rect 12293 5939 12327 5973
rect 12385 5939 12419 5973
rect 12477 5939 12511 5973
rect 12569 5939 12603 5973
rect 12661 5939 12695 5973
rect 12753 5939 12787 5973
rect 12845 5939 12879 5973
rect 12937 5939 12971 5973
rect 13029 5939 13063 5973
rect 13121 5939 13155 5973
rect 13213 5939 13247 5973
rect 13305 5939 13339 5973
rect 13397 5939 13431 5973
rect 13489 5939 13523 5973
rect 14067 5947 14101 5981
rect 14159 5947 14193 5981
rect 14251 5947 14285 5981
rect 14343 5947 14377 5981
rect 14435 5947 14469 5981
rect 14527 5947 14561 5981
rect 14619 5947 14653 5981
rect 14711 5947 14745 5981
rect 14803 5947 14837 5981
rect 14895 5947 14929 5981
rect 14987 5947 15021 5981
rect 15079 5947 15113 5981
rect 15171 5947 15205 5981
rect 15263 5947 15297 5981
rect 15355 5947 15389 5981
rect 15447 5947 15481 5981
rect 16061 5953 16095 5987
rect 16153 5953 16187 5987
rect 16245 5953 16279 5987
rect 16337 5953 16371 5987
rect 16429 5953 16463 5987
rect 16521 5953 16555 5987
rect 16613 5953 16647 5987
rect 16705 5953 16739 5987
rect 16797 5953 16831 5987
rect 16889 5953 16923 5987
rect 16981 5953 17015 5987
rect 17073 5953 17107 5987
rect 17165 5953 17199 5987
rect 17257 5953 17291 5987
rect 17349 5953 17383 5987
rect 17441 5953 17475 5987
rect 11150 5781 11184 5815
rect 10226 5727 10241 5747
rect 10241 5727 10260 5747
rect 10594 5743 10615 5747
rect 10615 5743 10628 5747
rect 10226 5713 10260 5727
rect 10594 5713 10628 5743
rect 1865 5531 1899 5565
rect 1957 5531 1991 5565
rect 2049 5531 2083 5565
rect 2141 5531 2175 5565
rect 2233 5531 2267 5565
rect 2325 5531 2359 5565
rect 2417 5531 2451 5565
rect 2509 5531 2543 5565
rect 2601 5531 2635 5565
rect 2693 5531 2727 5565
rect 2785 5531 2819 5565
rect 2877 5531 2911 5565
rect 2969 5531 3003 5565
rect 3061 5531 3095 5565
rect 3153 5531 3187 5565
rect 3245 5531 3279 5565
rect 2228 5361 2262 5395
rect 3999 5523 4033 5557
rect 4091 5523 4125 5557
rect 4183 5523 4217 5557
rect 4275 5523 4309 5557
rect 4367 5523 4401 5557
rect 4459 5523 4493 5557
rect 4551 5523 4585 5557
rect 4643 5523 4677 5557
rect 4735 5523 4769 5557
rect 4827 5523 4861 5557
rect 4919 5523 4953 5557
rect 5011 5523 5045 5557
rect 5103 5523 5137 5557
rect 5195 5523 5229 5557
rect 5287 5523 5321 5557
rect 5379 5523 5413 5557
rect 5951 5523 5985 5557
rect 6043 5523 6077 5557
rect 6135 5523 6169 5557
rect 6227 5523 6261 5557
rect 6319 5523 6353 5557
rect 6411 5523 6445 5557
rect 6503 5523 6537 5557
rect 6595 5523 6629 5557
rect 6687 5523 6721 5557
rect 6779 5523 6813 5557
rect 6871 5523 6905 5557
rect 6963 5523 6997 5557
rect 7055 5523 7089 5557
rect 7147 5523 7181 5557
rect 7239 5523 7273 5557
rect 7331 5523 7365 5557
rect 7953 5529 7987 5563
rect 8045 5529 8079 5563
rect 8137 5529 8171 5563
rect 8229 5529 8263 5563
rect 8321 5529 8355 5563
rect 8413 5529 8447 5563
rect 8505 5529 8539 5563
rect 8597 5529 8631 5563
rect 8689 5529 8723 5563
rect 8781 5529 8815 5563
rect 8873 5529 8907 5563
rect 8965 5529 8999 5563
rect 9057 5529 9091 5563
rect 9149 5529 9183 5563
rect 9241 5529 9275 5563
rect 9333 5529 9367 5563
rect 10318 5649 10352 5679
rect 10318 5645 10347 5649
rect 10347 5645 10352 5649
rect 10778 5665 10812 5679
rect 10778 5645 10783 5665
rect 10783 5645 10812 5665
rect 10966 5713 11000 5747
rect 11242 5719 11274 5747
rect 11274 5719 11276 5747
rect 11242 5713 11276 5719
rect 11150 5645 11184 5679
rect 10418 5580 10452 5614
rect 2968 5361 3002 5395
rect 2044 5307 2059 5327
rect 2059 5307 2078 5327
rect 2412 5323 2433 5327
rect 2433 5323 2446 5327
rect 2044 5293 2078 5307
rect 2412 5293 2446 5323
rect 2136 5229 2170 5259
rect 2136 5225 2165 5229
rect 2165 5225 2170 5229
rect 2596 5245 2630 5259
rect 2596 5225 2601 5245
rect 2601 5225 2630 5245
rect 2784 5293 2818 5327
rect 3060 5299 3092 5327
rect 3092 5299 3094 5327
rect 3060 5293 3094 5299
rect 2968 5225 3002 5259
rect 2236 5160 2270 5194
rect 3244 5176 3273 5186
rect 3273 5176 3284 5186
rect 3244 5150 3284 5176
rect 4362 5353 4396 5387
rect 5102 5353 5136 5387
rect 4178 5299 4193 5319
rect 4193 5299 4212 5319
rect 4546 5315 4567 5319
rect 4567 5315 4580 5319
rect 4178 5285 4212 5299
rect 4546 5285 4580 5315
rect 4270 5221 4304 5251
rect 4270 5217 4299 5221
rect 4299 5217 4304 5221
rect 4730 5237 4764 5251
rect 4730 5217 4735 5237
rect 4735 5217 4764 5237
rect 4918 5285 4952 5319
rect 5194 5291 5226 5319
rect 5226 5291 5228 5319
rect 5194 5285 5228 5291
rect 5102 5217 5136 5251
rect 4368 5150 4402 5184
rect 1865 4987 1899 5021
rect 1957 4987 1991 5021
rect 2049 4987 2083 5021
rect 2141 4987 2175 5021
rect 2233 4987 2267 5021
rect 2325 4987 2359 5021
rect 2417 4987 2451 5021
rect 2509 4987 2543 5021
rect 2601 4987 2635 5021
rect 2693 4987 2727 5021
rect 2785 4987 2819 5021
rect 2877 4987 2911 5021
rect 2969 4987 3003 5021
rect 3061 4987 3095 5021
rect 3153 4987 3187 5021
rect 3245 4987 3279 5021
rect 5384 5168 5407 5178
rect 5407 5168 5418 5178
rect 5384 5142 5418 5168
rect 6314 5353 6348 5387
rect 7054 5353 7088 5387
rect 6130 5299 6145 5319
rect 6145 5299 6164 5319
rect 6498 5315 6519 5319
rect 6519 5315 6532 5319
rect 6130 5285 6164 5299
rect 6498 5285 6532 5315
rect 6222 5221 6256 5251
rect 6222 5217 6251 5221
rect 6251 5217 6256 5221
rect 6682 5237 6716 5251
rect 6682 5217 6687 5237
rect 6687 5217 6716 5237
rect 6870 5285 6904 5319
rect 7146 5291 7178 5319
rect 7178 5291 7180 5319
rect 7146 5285 7180 5291
rect 7054 5217 7088 5251
rect 6320 5150 6354 5184
rect 7336 5168 7359 5178
rect 7359 5168 7370 5178
rect 7336 5142 7370 5168
rect 8316 5359 8350 5393
rect 9056 5359 9090 5393
rect 8132 5305 8147 5325
rect 8147 5305 8166 5325
rect 8500 5321 8521 5325
rect 8521 5321 8534 5325
rect 8132 5291 8166 5305
rect 8500 5291 8534 5321
rect 11426 5596 11455 5606
rect 11455 5596 11466 5606
rect 11426 5570 11466 5596
rect 12472 5769 12506 5803
rect 13212 5769 13246 5803
rect 12288 5715 12303 5735
rect 12303 5715 12322 5735
rect 12656 5731 12677 5735
rect 12677 5731 12690 5735
rect 12288 5701 12322 5715
rect 12656 5701 12690 5731
rect 12380 5637 12414 5667
rect 12380 5633 12409 5637
rect 12409 5633 12414 5637
rect 12840 5653 12874 5667
rect 12840 5633 12845 5653
rect 12845 5633 12874 5653
rect 13028 5701 13062 5735
rect 13304 5707 13336 5735
rect 13336 5707 13338 5735
rect 13304 5701 13338 5707
rect 13212 5633 13246 5667
rect 12478 5566 12512 5600
rect 10047 5407 10081 5441
rect 10139 5407 10173 5441
rect 10231 5407 10265 5441
rect 10323 5407 10357 5441
rect 10415 5407 10449 5441
rect 10507 5407 10541 5441
rect 10599 5407 10633 5441
rect 10691 5407 10725 5441
rect 10783 5407 10817 5441
rect 10875 5407 10909 5441
rect 10967 5407 11001 5441
rect 11059 5407 11093 5441
rect 11151 5407 11185 5441
rect 11243 5407 11277 5441
rect 11335 5407 11369 5441
rect 11427 5407 11461 5441
rect 13494 5584 13517 5594
rect 13517 5584 13528 5594
rect 13494 5558 13528 5584
rect 14430 5777 14464 5811
rect 15170 5777 15204 5811
rect 14246 5723 14261 5743
rect 14261 5723 14280 5743
rect 14614 5739 14635 5743
rect 14635 5739 14648 5743
rect 14246 5709 14280 5723
rect 14614 5709 14648 5739
rect 14338 5645 14372 5675
rect 14338 5641 14367 5645
rect 14367 5641 14372 5645
rect 14798 5661 14832 5675
rect 14798 5641 14803 5661
rect 14803 5641 14832 5661
rect 14986 5709 15020 5743
rect 15262 5715 15294 5743
rect 15294 5715 15296 5743
rect 15262 5709 15296 5715
rect 15170 5641 15204 5675
rect 14436 5574 14470 5608
rect 15452 5592 15475 5602
rect 15475 5592 15486 5602
rect 15452 5566 15486 5592
rect 16424 5783 16458 5817
rect 17164 5783 17198 5817
rect 16240 5729 16255 5749
rect 16255 5729 16274 5749
rect 16608 5745 16629 5749
rect 16629 5745 16642 5749
rect 16240 5715 16274 5729
rect 16608 5715 16642 5745
rect 16332 5651 16366 5681
rect 16332 5647 16361 5651
rect 16361 5647 16366 5651
rect 16792 5667 16826 5681
rect 16792 5647 16797 5667
rect 16797 5647 16826 5667
rect 16980 5715 17014 5749
rect 17256 5721 17288 5749
rect 17288 5721 17290 5749
rect 17256 5715 17290 5721
rect 17164 5647 17198 5681
rect 16430 5580 16464 5614
rect 17446 5598 17469 5608
rect 17469 5598 17480 5608
rect 17446 5572 17480 5598
rect 12109 5395 12143 5429
rect 12201 5395 12235 5429
rect 12293 5395 12327 5429
rect 12385 5395 12419 5429
rect 12477 5395 12511 5429
rect 12569 5395 12603 5429
rect 12661 5395 12695 5429
rect 12753 5395 12787 5429
rect 12845 5395 12879 5429
rect 12937 5395 12971 5429
rect 13029 5395 13063 5429
rect 13121 5395 13155 5429
rect 13213 5395 13247 5429
rect 13305 5395 13339 5429
rect 13397 5395 13431 5429
rect 13489 5395 13523 5429
rect 14067 5403 14101 5437
rect 14159 5403 14193 5437
rect 14251 5403 14285 5437
rect 14343 5403 14377 5437
rect 14435 5403 14469 5437
rect 14527 5403 14561 5437
rect 14619 5403 14653 5437
rect 14711 5403 14745 5437
rect 14803 5403 14837 5437
rect 14895 5403 14929 5437
rect 14987 5403 15021 5437
rect 15079 5403 15113 5437
rect 15171 5403 15205 5437
rect 15263 5403 15297 5437
rect 15355 5403 15389 5437
rect 15447 5403 15481 5437
rect 16061 5409 16095 5443
rect 16153 5409 16187 5443
rect 16245 5409 16279 5443
rect 16337 5409 16371 5443
rect 16429 5409 16463 5443
rect 16521 5409 16555 5443
rect 16613 5409 16647 5443
rect 16705 5409 16739 5443
rect 16797 5409 16831 5443
rect 16889 5409 16923 5443
rect 16981 5409 17015 5443
rect 17073 5409 17107 5443
rect 17165 5409 17199 5443
rect 17257 5409 17291 5443
rect 17349 5409 17383 5443
rect 17441 5409 17475 5443
rect 8224 5227 8258 5257
rect 8224 5223 8253 5227
rect 8253 5223 8258 5227
rect 8684 5243 8718 5257
rect 8684 5223 8689 5243
rect 8689 5223 8718 5243
rect 8872 5291 8906 5325
rect 9148 5297 9180 5325
rect 9180 5297 9182 5325
rect 9148 5291 9182 5297
rect 9056 5223 9090 5257
rect 8322 5156 8356 5190
rect 18608 5188 18642 5222
rect 9338 5174 9361 5184
rect 9361 5174 9372 5184
rect 9338 5148 9372 5174
rect 18690 5160 18724 5194
rect 10075 5077 10109 5111
rect 10167 5077 10201 5111
rect 10259 5077 10293 5111
rect 10351 5077 10385 5111
rect 10443 5077 10477 5111
rect 10535 5077 10569 5111
rect 10627 5077 10661 5111
rect 10719 5077 10753 5111
rect 10811 5077 10845 5111
rect 10903 5077 10937 5111
rect 10995 5077 11029 5111
rect 11087 5077 11121 5111
rect 11179 5077 11213 5111
rect 11271 5077 11305 5111
rect 11363 5077 11397 5111
rect 11455 5077 11489 5111
rect 3999 4979 4033 5013
rect 4091 4979 4125 5013
rect 4183 4979 4217 5013
rect 4275 4979 4309 5013
rect 4367 4979 4401 5013
rect 4459 4979 4493 5013
rect 4551 4979 4585 5013
rect 4643 4979 4677 5013
rect 4735 4979 4769 5013
rect 4827 4979 4861 5013
rect 4919 4979 4953 5013
rect 5011 4979 5045 5013
rect 5103 4979 5137 5013
rect 5195 4979 5229 5013
rect 5287 4979 5321 5013
rect 5379 4979 5413 5013
rect 5951 4979 5985 5013
rect 6043 4979 6077 5013
rect 6135 4979 6169 5013
rect 6227 4979 6261 5013
rect 6319 4979 6353 5013
rect 6411 4979 6445 5013
rect 6503 4979 6537 5013
rect 6595 4979 6629 5013
rect 6687 4979 6721 5013
rect 6779 4979 6813 5013
rect 6871 4979 6905 5013
rect 6963 4979 6997 5013
rect 7055 4979 7089 5013
rect 7147 4979 7181 5013
rect 7239 4979 7273 5013
rect 7331 4979 7365 5013
rect 7953 4985 7987 5019
rect 8045 4985 8079 5019
rect 8137 4985 8171 5019
rect 8229 4985 8263 5019
rect 8321 4985 8355 5019
rect 8413 4985 8447 5019
rect 8505 4985 8539 5019
rect 8597 4985 8631 5019
rect 8689 4985 8723 5019
rect 8781 4985 8815 5019
rect 8873 4985 8907 5019
rect 8965 4985 8999 5019
rect 9057 4985 9091 5019
rect 9149 4985 9183 5019
rect 9241 4985 9275 5019
rect 9333 4985 9367 5019
rect 10438 4907 10472 4941
rect 18432 5070 18470 5108
rect 12345 5033 12379 5067
rect 12437 5033 12471 5067
rect 12529 5033 12563 5067
rect 12621 5033 12655 5067
rect 12713 5033 12747 5067
rect 12805 5033 12839 5067
rect 12897 5033 12931 5067
rect 12989 5033 13023 5067
rect 13081 5033 13115 5067
rect 13173 5033 13207 5067
rect 13265 5033 13299 5067
rect 13357 5033 13391 5067
rect 13449 5033 13483 5067
rect 13541 5033 13575 5067
rect 13633 5033 13667 5067
rect 13725 5033 13759 5067
rect 11178 4907 11212 4941
rect 10254 4853 10269 4873
rect 10269 4853 10288 4873
rect 10622 4869 10643 4873
rect 10643 4869 10656 4873
rect 10254 4839 10288 4853
rect 10622 4839 10656 4869
rect 10346 4775 10380 4805
rect 10346 4771 10375 4775
rect 10375 4771 10380 4775
rect 10806 4791 10840 4805
rect 10806 4771 10811 4791
rect 10811 4771 10840 4791
rect 10994 4839 11028 4873
rect 11270 4845 11302 4873
rect 11302 4845 11304 4873
rect 11270 4839 11304 4845
rect 11178 4771 11212 4805
rect 10446 4706 10480 4740
rect 11454 4722 11483 4732
rect 11483 4722 11494 4732
rect 11454 4696 11494 4722
rect 12708 4863 12742 4897
rect 14347 5027 14381 5061
rect 14439 5027 14473 5061
rect 14531 5027 14565 5061
rect 14623 5027 14657 5061
rect 14715 5027 14749 5061
rect 14807 5027 14841 5061
rect 14899 5027 14933 5061
rect 14991 5027 15025 5061
rect 15083 5027 15117 5061
rect 15175 5027 15209 5061
rect 15267 5027 15301 5061
rect 15359 5027 15393 5061
rect 15451 5027 15485 5061
rect 15543 5027 15577 5061
rect 15635 5027 15669 5061
rect 15727 5027 15761 5061
rect 13448 4863 13482 4897
rect 12524 4809 12539 4829
rect 12539 4809 12558 4829
rect 12892 4825 12913 4829
rect 12913 4825 12926 4829
rect 12524 4795 12558 4809
rect 12892 4795 12926 4825
rect 12616 4731 12650 4761
rect 12616 4727 12645 4731
rect 12645 4727 12650 4731
rect 13076 4747 13110 4761
rect 13076 4727 13081 4747
rect 13081 4727 13110 4747
rect 13264 4795 13298 4829
rect 13540 4801 13572 4829
rect 13572 4801 13574 4829
rect 13540 4795 13574 4801
rect 13448 4727 13482 4761
rect 12714 4660 12748 4694
rect 10075 4533 10109 4567
rect 10167 4533 10201 4567
rect 10259 4533 10293 4567
rect 10351 4533 10385 4567
rect 10443 4533 10477 4567
rect 10535 4533 10569 4567
rect 10627 4533 10661 4567
rect 10719 4533 10753 4567
rect 10811 4533 10845 4567
rect 10903 4533 10937 4567
rect 10995 4533 11029 4567
rect 11087 4533 11121 4567
rect 11179 4533 11213 4567
rect 11271 4533 11305 4567
rect 11363 4533 11397 4567
rect 11455 4533 11489 4567
rect 13730 4678 13753 4688
rect 13753 4678 13764 4688
rect 13730 4652 13764 4678
rect 14710 4857 14744 4891
rect 16369 5009 16403 5043
rect 16461 5009 16495 5043
rect 16553 5009 16587 5043
rect 16645 5009 16679 5043
rect 16737 5009 16771 5043
rect 16829 5009 16863 5043
rect 16921 5009 16955 5043
rect 17013 5009 17047 5043
rect 17105 5009 17139 5043
rect 17197 5009 17231 5043
rect 17289 5009 17323 5043
rect 17381 5009 17415 5043
rect 17473 5009 17507 5043
rect 17565 5009 17599 5043
rect 17657 5009 17691 5043
rect 17749 5009 17783 5043
rect 15450 4857 15484 4891
rect 14526 4803 14541 4823
rect 14541 4803 14560 4823
rect 14894 4819 14915 4823
rect 14915 4819 14928 4823
rect 14526 4789 14560 4803
rect 14894 4789 14928 4819
rect 14618 4725 14652 4755
rect 14618 4721 14647 4725
rect 14647 4721 14652 4725
rect 15078 4741 15112 4755
rect 15078 4721 15083 4741
rect 15083 4721 15112 4741
rect 15266 4789 15300 4823
rect 15542 4795 15574 4823
rect 15574 4795 15576 4823
rect 15542 4789 15576 4795
rect 15450 4721 15484 4755
rect 14716 4654 14750 4688
rect 12345 4489 12379 4523
rect 12437 4489 12471 4523
rect 12529 4489 12563 4523
rect 12621 4489 12655 4523
rect 12713 4489 12747 4523
rect 12805 4489 12839 4523
rect 12897 4489 12931 4523
rect 12989 4489 13023 4523
rect 13081 4489 13115 4523
rect 13173 4489 13207 4523
rect 13265 4489 13299 4523
rect 13357 4489 13391 4523
rect 13449 4489 13483 4523
rect 13541 4489 13575 4523
rect 13633 4489 13667 4523
rect 13725 4489 13759 4523
rect 15732 4672 15755 4682
rect 15755 4672 15766 4682
rect 15732 4646 15766 4672
rect 16732 4839 16766 4873
rect 19064 5004 19102 5042
rect 17472 4839 17506 4873
rect 16548 4785 16563 4805
rect 16563 4785 16582 4805
rect 16916 4801 16937 4805
rect 16937 4801 16950 4805
rect 16548 4771 16582 4785
rect 16916 4771 16950 4801
rect 16640 4707 16674 4737
rect 16640 4703 16669 4707
rect 16669 4703 16674 4707
rect 17100 4723 17134 4737
rect 17100 4703 17105 4723
rect 17105 4703 17134 4723
rect 17288 4771 17322 4805
rect 17564 4777 17596 4805
rect 17596 4777 17598 4805
rect 17564 4771 17598 4777
rect 17472 4703 17506 4737
rect 16738 4636 16772 4670
rect 14347 4483 14381 4517
rect 14439 4483 14473 4517
rect 14531 4483 14565 4517
rect 14623 4483 14657 4517
rect 14715 4483 14749 4517
rect 14807 4483 14841 4517
rect 14899 4483 14933 4517
rect 14991 4483 15025 4517
rect 15083 4483 15117 4517
rect 15175 4483 15209 4517
rect 15267 4483 15301 4517
rect 15359 4483 15393 4517
rect 15451 4483 15485 4517
rect 15543 4483 15577 4517
rect 15635 4483 15669 4517
rect 15727 4483 15761 4517
rect 17754 4654 17777 4664
rect 17777 4654 17788 4664
rect 17754 4628 17788 4654
rect 16369 4465 16403 4499
rect 16461 4465 16495 4499
rect 16553 4465 16587 4499
rect 16645 4465 16679 4499
rect 16737 4465 16771 4499
rect 16829 4465 16863 4499
rect 16921 4465 16955 4499
rect 17013 4465 17047 4499
rect 17105 4465 17139 4499
rect 17197 4465 17231 4499
rect 17289 4465 17323 4499
rect 17381 4465 17415 4499
rect 17473 4465 17507 4499
rect 17565 4465 17599 4499
rect 17657 4465 17691 4499
rect 17749 4465 17783 4499
rect 6148 3088 6182 3122
rect 6244 3090 6278 3124
rect 1835 2271 1869 2305
rect 1927 2271 1961 2305
rect 2019 2271 2053 2305
rect 2111 2271 2145 2305
rect 2203 2271 2237 2305
rect 2295 2271 2329 2305
rect 2387 2271 2421 2305
rect 2479 2271 2513 2305
rect 2571 2271 2605 2305
rect 2663 2271 2697 2305
rect 2755 2271 2789 2305
rect 2847 2271 2881 2305
rect 2939 2271 2973 2305
rect 3031 2271 3065 2305
rect 3123 2271 3157 2305
rect 3215 2271 3249 2305
rect 2198 2101 2232 2135
rect 3905 2267 3939 2301
rect 3997 2267 4031 2301
rect 4089 2267 4123 2301
rect 4181 2267 4215 2301
rect 4273 2267 4307 2301
rect 4365 2267 4399 2301
rect 4457 2267 4491 2301
rect 4549 2267 4583 2301
rect 4641 2267 4675 2301
rect 4733 2267 4767 2301
rect 4825 2267 4859 2301
rect 4917 2267 4951 2301
rect 5009 2267 5043 2301
rect 5101 2267 5135 2301
rect 5193 2267 5227 2301
rect 5285 2267 5319 2301
rect 5857 2267 5891 2301
rect 5949 2267 5983 2301
rect 6041 2267 6075 2301
rect 6133 2267 6167 2301
rect 6225 2267 6259 2301
rect 6317 2267 6351 2301
rect 6409 2267 6443 2301
rect 6501 2267 6535 2301
rect 6593 2267 6627 2301
rect 6685 2267 6719 2301
rect 6777 2267 6811 2301
rect 6869 2267 6903 2301
rect 6961 2267 6995 2301
rect 7053 2267 7087 2301
rect 7145 2267 7179 2301
rect 7237 2267 7271 2301
rect 7859 2273 7893 2307
rect 7951 2273 7985 2307
rect 8043 2273 8077 2307
rect 8135 2273 8169 2307
rect 8227 2273 8261 2307
rect 8319 2273 8353 2307
rect 8411 2273 8445 2307
rect 8503 2273 8537 2307
rect 8595 2273 8629 2307
rect 8687 2273 8721 2307
rect 8779 2273 8813 2307
rect 8871 2273 8905 2307
rect 8963 2273 8997 2307
rect 9055 2273 9089 2307
rect 9147 2273 9181 2307
rect 9239 2273 9273 2307
rect 9811 2273 9845 2307
rect 9903 2273 9937 2307
rect 9995 2273 10029 2307
rect 10087 2273 10121 2307
rect 10179 2273 10213 2307
rect 10271 2273 10305 2307
rect 10363 2273 10397 2307
rect 10455 2273 10489 2307
rect 10547 2273 10581 2307
rect 10639 2273 10673 2307
rect 10731 2273 10765 2307
rect 10823 2273 10857 2307
rect 10915 2273 10949 2307
rect 11007 2273 11041 2307
rect 11099 2273 11133 2307
rect 11191 2273 11225 2307
rect 11803 2273 11837 2307
rect 11895 2273 11929 2307
rect 11987 2273 12021 2307
rect 12079 2273 12113 2307
rect 12171 2273 12205 2307
rect 12263 2273 12297 2307
rect 12355 2273 12389 2307
rect 12447 2273 12481 2307
rect 12539 2273 12573 2307
rect 12631 2273 12665 2307
rect 12723 2273 12757 2307
rect 12815 2273 12849 2307
rect 12907 2273 12941 2307
rect 12999 2273 13033 2307
rect 13091 2273 13125 2307
rect 13183 2273 13217 2307
rect 13755 2273 13789 2307
rect 13847 2273 13881 2307
rect 13939 2273 13973 2307
rect 14031 2273 14065 2307
rect 14123 2273 14157 2307
rect 14215 2273 14249 2307
rect 14307 2273 14341 2307
rect 14399 2273 14433 2307
rect 14491 2273 14525 2307
rect 14583 2273 14617 2307
rect 14675 2273 14709 2307
rect 14767 2273 14801 2307
rect 14859 2273 14893 2307
rect 14951 2273 14985 2307
rect 15043 2273 15077 2307
rect 15135 2273 15169 2307
rect 15819 2273 15853 2307
rect 15911 2273 15945 2307
rect 16003 2273 16037 2307
rect 16095 2273 16129 2307
rect 16187 2273 16221 2307
rect 16279 2273 16313 2307
rect 16371 2273 16405 2307
rect 16463 2273 16497 2307
rect 16555 2273 16589 2307
rect 16647 2273 16681 2307
rect 16739 2273 16773 2307
rect 16831 2273 16865 2307
rect 16923 2273 16957 2307
rect 17015 2273 17049 2307
rect 17107 2273 17141 2307
rect 17199 2273 17233 2307
rect 2938 2101 2972 2135
rect 2014 2047 2029 2067
rect 2029 2047 2048 2067
rect 2382 2063 2403 2067
rect 2403 2063 2416 2067
rect 2014 2033 2048 2047
rect 2382 2033 2416 2063
rect 2106 1969 2140 1999
rect 2106 1965 2135 1969
rect 2135 1965 2140 1969
rect 2566 1985 2600 1999
rect 2566 1965 2571 1985
rect 2571 1965 2600 1985
rect 2754 2033 2788 2067
rect 3030 2039 3062 2067
rect 3062 2039 3064 2067
rect 3030 2033 3064 2039
rect 2938 1965 2972 1999
rect 2206 1900 2240 1934
rect 3214 1916 3243 1926
rect 3243 1916 3254 1926
rect 3214 1890 3254 1916
rect 4268 2097 4302 2131
rect 5008 2097 5042 2131
rect 4084 2043 4099 2063
rect 4099 2043 4118 2063
rect 4452 2059 4473 2063
rect 4473 2059 4486 2063
rect 4084 2029 4118 2043
rect 4452 2029 4486 2059
rect 4176 1965 4210 1995
rect 4176 1961 4205 1965
rect 4205 1961 4210 1965
rect 4636 1981 4670 1995
rect 4636 1961 4641 1981
rect 4641 1961 4670 1981
rect 4824 2029 4858 2063
rect 5100 2035 5132 2063
rect 5132 2035 5134 2063
rect 5100 2029 5134 2035
rect 5008 1961 5042 1995
rect 4274 1894 4308 1928
rect 1835 1727 1869 1761
rect 1927 1727 1961 1761
rect 2019 1727 2053 1761
rect 2111 1727 2145 1761
rect 2203 1727 2237 1761
rect 2295 1727 2329 1761
rect 2387 1727 2421 1761
rect 2479 1727 2513 1761
rect 2571 1727 2605 1761
rect 2663 1727 2697 1761
rect 2755 1727 2789 1761
rect 2847 1727 2881 1761
rect 2939 1727 2973 1761
rect 3031 1727 3065 1761
rect 3123 1727 3157 1761
rect 3215 1727 3249 1761
rect 5290 1912 5313 1922
rect 5313 1912 5324 1922
rect 5290 1886 5324 1912
rect 6220 2097 6254 2131
rect 6960 2097 6994 2131
rect 6036 2043 6051 2063
rect 6051 2043 6070 2063
rect 6404 2059 6425 2063
rect 6425 2059 6438 2063
rect 6036 2029 6070 2043
rect 6404 2029 6438 2059
rect 6128 1965 6162 1995
rect 6128 1961 6157 1965
rect 6157 1961 6162 1965
rect 6588 1981 6622 1995
rect 6588 1961 6593 1981
rect 6593 1961 6622 1981
rect 6776 2029 6810 2063
rect 7052 2035 7084 2063
rect 7084 2035 7086 2063
rect 7052 2029 7086 2035
rect 6960 1961 6994 1995
rect 6226 1894 6260 1928
rect 7242 1912 7265 1922
rect 7265 1912 7276 1922
rect 7242 1886 7276 1912
rect 8222 2103 8256 2137
rect 8962 2103 8996 2137
rect 8038 2049 8053 2069
rect 8053 2049 8072 2069
rect 8406 2065 8427 2069
rect 8427 2065 8440 2069
rect 8038 2035 8072 2049
rect 8406 2035 8440 2065
rect 8130 1971 8164 2001
rect 8130 1967 8159 1971
rect 8159 1967 8164 1971
rect 8590 1987 8624 2001
rect 8590 1967 8595 1987
rect 8595 1967 8624 1987
rect 8778 2035 8812 2069
rect 9054 2041 9086 2069
rect 9086 2041 9088 2069
rect 9054 2035 9088 2041
rect 8962 1967 8996 2001
rect 8228 1900 8262 1934
rect 9244 1918 9267 1928
rect 9267 1918 9278 1928
rect 9244 1892 9278 1918
rect 10174 2103 10208 2137
rect 10914 2103 10948 2137
rect 9990 2049 10005 2069
rect 10005 2049 10024 2069
rect 10358 2065 10379 2069
rect 10379 2065 10392 2069
rect 9990 2035 10024 2049
rect 10358 2035 10392 2065
rect 10082 1971 10116 2001
rect 10082 1967 10111 1971
rect 10111 1967 10116 1971
rect 10542 1987 10576 2001
rect 10542 1967 10547 1987
rect 10547 1967 10576 1987
rect 10730 2035 10764 2069
rect 11006 2041 11038 2069
rect 11038 2041 11040 2069
rect 11006 2035 11040 2041
rect 10914 1967 10948 2001
rect 10180 1900 10214 1934
rect 11196 1918 11219 1928
rect 11219 1918 11230 1928
rect 11196 1892 11230 1918
rect 12166 2103 12200 2137
rect 12906 2103 12940 2137
rect 11982 2049 11997 2069
rect 11997 2049 12016 2069
rect 12350 2065 12371 2069
rect 12371 2065 12384 2069
rect 11982 2035 12016 2049
rect 12350 2035 12384 2065
rect 12074 1971 12108 2001
rect 12074 1967 12103 1971
rect 12103 1967 12108 1971
rect 12534 1987 12568 2001
rect 12534 1967 12539 1987
rect 12539 1967 12568 1987
rect 12722 2035 12756 2069
rect 12998 2041 13030 2069
rect 13030 2041 13032 2069
rect 12998 2035 13032 2041
rect 12906 1967 12940 2001
rect 12172 1900 12206 1934
rect 13188 1918 13211 1928
rect 13211 1918 13222 1928
rect 13188 1892 13222 1918
rect 14118 2103 14152 2137
rect 14858 2103 14892 2137
rect 13934 2049 13949 2069
rect 13949 2049 13968 2069
rect 14302 2065 14323 2069
rect 14323 2065 14336 2069
rect 13934 2035 13968 2049
rect 14302 2035 14336 2065
rect 14026 1971 14060 2001
rect 14026 1967 14055 1971
rect 14055 1967 14060 1971
rect 14486 1987 14520 2001
rect 14486 1967 14491 1987
rect 14491 1967 14520 1987
rect 14674 2035 14708 2069
rect 14950 2041 14982 2069
rect 14982 2041 14984 2069
rect 14950 2035 14984 2041
rect 14858 1967 14892 2001
rect 14124 1900 14158 1934
rect 15140 1918 15163 1928
rect 15163 1918 15174 1928
rect 15140 1892 15174 1918
rect 16182 2103 16216 2137
rect 16922 2103 16956 2137
rect 15998 2049 16013 2069
rect 16013 2049 16032 2069
rect 16366 2065 16387 2069
rect 16387 2065 16400 2069
rect 15998 2035 16032 2049
rect 16366 2035 16400 2065
rect 16090 1971 16124 2001
rect 16090 1967 16119 1971
rect 16119 1967 16124 1971
rect 16550 1987 16584 2001
rect 16550 1967 16555 1987
rect 16555 1967 16584 1987
rect 16738 2035 16772 2069
rect 17014 2041 17046 2069
rect 17046 2041 17048 2069
rect 17014 2035 17048 2041
rect 16922 1967 16956 2001
rect 16188 1900 16222 1934
rect 17204 1918 17227 1928
rect 17227 1918 17238 1928
rect 17204 1892 17238 1918
rect 3905 1723 3939 1757
rect 3997 1723 4031 1757
rect 4089 1723 4123 1757
rect 4181 1723 4215 1757
rect 4273 1723 4307 1757
rect 4365 1723 4399 1757
rect 4457 1723 4491 1757
rect 4549 1723 4583 1757
rect 4641 1723 4675 1757
rect 4733 1723 4767 1757
rect 4825 1723 4859 1757
rect 4917 1723 4951 1757
rect 5009 1723 5043 1757
rect 5101 1723 5135 1757
rect 5193 1723 5227 1757
rect 5285 1723 5319 1757
rect 5857 1723 5891 1757
rect 5949 1723 5983 1757
rect 6041 1723 6075 1757
rect 6133 1723 6167 1757
rect 6225 1723 6259 1757
rect 6317 1723 6351 1757
rect 6409 1723 6443 1757
rect 6501 1723 6535 1757
rect 6593 1723 6627 1757
rect 6685 1723 6719 1757
rect 6777 1723 6811 1757
rect 6869 1723 6903 1757
rect 6961 1723 6995 1757
rect 7053 1723 7087 1757
rect 7145 1723 7179 1757
rect 7237 1723 7271 1757
rect 7859 1729 7893 1763
rect 7951 1729 7985 1763
rect 8043 1729 8077 1763
rect 8135 1729 8169 1763
rect 8227 1729 8261 1763
rect 8319 1729 8353 1763
rect 8411 1729 8445 1763
rect 8503 1729 8537 1763
rect 8595 1729 8629 1763
rect 8687 1729 8721 1763
rect 8779 1729 8813 1763
rect 8871 1729 8905 1763
rect 8963 1729 8997 1763
rect 9055 1729 9089 1763
rect 9147 1729 9181 1763
rect 9239 1729 9273 1763
rect 9811 1729 9845 1763
rect 9903 1729 9937 1763
rect 9995 1729 10029 1763
rect 10087 1729 10121 1763
rect 10179 1729 10213 1763
rect 10271 1729 10305 1763
rect 10363 1729 10397 1763
rect 10455 1729 10489 1763
rect 10547 1729 10581 1763
rect 10639 1729 10673 1763
rect 10731 1729 10765 1763
rect 10823 1729 10857 1763
rect 10915 1729 10949 1763
rect 11007 1729 11041 1763
rect 11099 1729 11133 1763
rect 11191 1729 11225 1763
rect 11803 1729 11837 1763
rect 11895 1729 11929 1763
rect 11987 1729 12021 1763
rect 12079 1729 12113 1763
rect 12171 1729 12205 1763
rect 12263 1729 12297 1763
rect 12355 1729 12389 1763
rect 12447 1729 12481 1763
rect 12539 1729 12573 1763
rect 12631 1729 12665 1763
rect 12723 1729 12757 1763
rect 12815 1729 12849 1763
rect 12907 1729 12941 1763
rect 12999 1729 13033 1763
rect 13091 1729 13125 1763
rect 13183 1729 13217 1763
rect 13755 1729 13789 1763
rect 13847 1729 13881 1763
rect 13939 1729 13973 1763
rect 14031 1729 14065 1763
rect 14123 1729 14157 1763
rect 14215 1729 14249 1763
rect 14307 1729 14341 1763
rect 14399 1729 14433 1763
rect 14491 1729 14525 1763
rect 14583 1729 14617 1763
rect 14675 1729 14709 1763
rect 14767 1729 14801 1763
rect 14859 1729 14893 1763
rect 14951 1729 14985 1763
rect 15043 1729 15077 1763
rect 15135 1729 15169 1763
rect 15819 1729 15853 1763
rect 15911 1729 15945 1763
rect 16003 1729 16037 1763
rect 16095 1729 16129 1763
rect 16187 1729 16221 1763
rect 16279 1729 16313 1763
rect 16371 1729 16405 1763
rect 16463 1729 16497 1763
rect 16555 1729 16589 1763
rect 16647 1729 16681 1763
rect 16739 1729 16773 1763
rect 16831 1729 16865 1763
rect 16923 1729 16957 1763
rect 17015 1729 17049 1763
rect 17107 1729 17141 1763
rect 17199 1729 17233 1763
<< metal1 >>
rect 18590 44096 19128 44168
rect 18590 43898 18768 44096
rect 18962 43898 19128 44096
rect 18590 43828 19128 43898
rect 18866 43294 18936 43828
rect 18866 43258 18882 43294
rect 18916 43258 18936 43294
rect 18866 43244 18936 43258
rect 18856 42024 18938 42050
rect 18856 41990 18886 42024
rect 18920 41990 18938 42024
rect 18856 41398 18938 41990
rect 18856 41364 18868 41398
rect 18902 41364 18938 41398
rect 18856 41346 18938 41364
rect 18846 40468 18914 40510
rect 18846 40434 18870 40468
rect 18904 40434 18914 40468
rect 18846 39606 18914 40434
rect 18846 39570 18862 39606
rect 18896 39570 18914 39606
rect 18846 39554 18914 39570
rect 18864 39090 18946 39114
rect 18864 39056 18876 39090
rect 18910 39056 18946 39090
rect 18864 38340 18946 39056
rect 18864 38306 18886 38340
rect 18920 38306 18946 38340
rect 18864 38284 18946 38306
rect 18872 37794 18934 37954
rect 18872 37760 18888 37794
rect 18922 37760 18934 37794
rect 18872 37198 18934 37760
rect 18870 37192 18952 37198
rect 18870 37158 18892 37192
rect 18926 37158 18952 37192
rect 18870 37144 18952 37158
rect 18886 36920 18950 36928
rect 18886 36884 18900 36920
rect 18934 36884 18950 36920
rect 18886 36868 18950 36884
rect 18898 36236 18944 36868
rect 18890 36226 18954 36236
rect 18890 36190 18904 36226
rect 18940 36190 18954 36226
rect 18890 36176 18954 36190
rect 18896 36130 18958 36146
rect 18896 36094 18904 36130
rect 18948 36094 18958 36130
rect 18896 36080 18958 36094
rect 18911 35879 18953 36080
rect 18870 35837 18953 35879
rect 18418 35197 18514 35226
rect 18418 35163 18449 35197
rect 18483 35163 18514 35197
rect 18418 35105 18514 35163
rect 18418 35071 18449 35105
rect 18483 35071 18514 35105
rect 18418 35013 18514 35071
rect 18632 35106 18736 35126
rect 18632 35070 18664 35106
rect 18698 35102 18736 35106
rect 18698 35070 18754 35102
rect 18632 35052 18754 35070
rect 18632 35050 18736 35052
rect 18418 34979 18449 35013
rect 18483 34979 18514 35013
rect 18418 34921 18514 34979
rect 18418 34887 18449 34921
rect 18483 34887 18514 34921
rect 18418 34829 18514 34887
rect 18418 34795 18449 34829
rect 18483 34795 18514 34829
rect 18418 34737 18514 34795
rect 18418 34703 18449 34737
rect 18483 34703 18514 34737
rect 18418 34645 18514 34703
rect 18418 34611 18449 34645
rect 18483 34611 18514 34645
rect 18418 34553 18514 34611
rect 18418 34519 18449 34553
rect 18483 34519 18514 34553
rect 18661 34604 18732 35050
rect 18870 34834 18912 35837
rect 18962 35197 19058 35226
rect 18962 35163 18993 35197
rect 19027 35163 19058 35197
rect 18962 35105 19058 35163
rect 18962 35071 18993 35105
rect 19027 35071 19058 35105
rect 18962 35013 19058 35071
rect 18962 34979 18993 35013
rect 19027 34979 19058 35013
rect 18962 34921 19058 34979
rect 18962 34887 18993 34921
rect 19027 34887 19058 34921
rect 18846 34820 18934 34834
rect 18846 34782 18868 34820
rect 18906 34782 18934 34820
rect 18846 34774 18934 34782
rect 18962 34829 19058 34887
rect 18962 34795 18993 34829
rect 19027 34795 19058 34829
rect 18962 34737 19058 34795
rect 18962 34703 18993 34737
rect 19027 34703 19058 34737
rect 18962 34645 19058 34703
rect 18962 34611 18993 34645
rect 19027 34611 19058 34645
rect 18661 34533 18867 34604
rect 18418 34461 18514 34519
rect 18418 34454 18449 34461
rect 18483 34454 18514 34461
rect 18418 34372 18424 34454
rect 18504 34372 18514 34454
rect 18418 34369 18514 34372
rect 18418 34335 18449 34369
rect 18483 34335 18514 34369
rect 18418 34277 18514 34335
rect 18681 34367 18727 34379
rect 18681 34333 18687 34367
rect 18721 34333 18727 34367
rect 18681 34321 18727 34333
rect 18418 34243 18449 34277
rect 18483 34243 18514 34277
rect 18418 34185 18514 34243
rect 18613 34280 18659 34292
rect 18613 34246 18619 34280
rect 18653 34246 18659 34280
rect 18613 34234 18659 34246
rect 18418 34151 18449 34185
rect 18483 34151 18514 34185
rect 18418 34093 18514 34151
rect 18418 34059 18449 34093
rect 18483 34059 18514 34093
rect 18418 34001 18514 34059
rect 18418 33967 18449 34001
rect 18483 33967 18514 34001
rect 18622 33978 18650 34234
rect 18418 33909 18514 33967
rect 18613 33966 18659 33978
rect 18613 33932 18619 33966
rect 18653 33932 18659 33966
rect 18613 33920 18659 33932
rect 18418 33875 18449 33909
rect 18483 33875 18514 33909
rect 18418 33817 18514 33875
rect 18418 33783 18449 33817
rect 18483 33783 18514 33817
rect 18418 33725 18514 33783
rect 18418 33691 18449 33725
rect 18483 33691 18514 33725
rect 18418 33633 18514 33691
rect 18418 33599 18449 33633
rect 18483 33599 18514 33633
rect 18418 33541 18514 33599
rect 18622 33558 18650 33920
rect 18690 33875 18718 34321
rect 18681 33863 18727 33875
rect 18681 33829 18687 33863
rect 18721 33829 18727 33863
rect 18681 33817 18727 33829
rect 18690 33637 18718 33817
rect 18796 33706 18867 34533
rect 18796 33670 18816 33706
rect 18852 33670 18867 33706
rect 18796 33660 18867 33670
rect 18962 34553 19058 34611
rect 18962 34519 18993 34553
rect 19027 34519 19058 34553
rect 18962 34461 19058 34519
rect 18962 34458 18993 34461
rect 19027 34458 19058 34461
rect 18962 34376 18972 34458
rect 19052 34376 19058 34458
rect 18962 34369 19058 34376
rect 18962 34335 18993 34369
rect 19027 34335 19058 34369
rect 18962 34277 19058 34335
rect 18962 34243 18993 34277
rect 19027 34243 19058 34277
rect 18962 34185 19058 34243
rect 18962 34151 18993 34185
rect 19027 34151 19058 34185
rect 18962 34093 19058 34151
rect 18962 34059 18993 34093
rect 19027 34059 19058 34093
rect 18962 34001 19058 34059
rect 18962 33967 18993 34001
rect 19027 33967 19058 34001
rect 18962 33909 19058 33967
rect 18962 33875 18993 33909
rect 19027 33875 19058 33909
rect 18962 33817 19058 33875
rect 18962 33783 18993 33817
rect 19027 33783 19058 33817
rect 18962 33725 19058 33783
rect 18962 33691 18993 33725
rect 19027 33691 19058 33725
rect 18681 33625 18727 33637
rect 18681 33591 18687 33625
rect 18721 33591 18727 33625
rect 18681 33579 18727 33591
rect 18962 33633 19058 33691
rect 18962 33599 18993 33633
rect 19027 33599 19058 33633
rect 18418 33507 18449 33541
rect 18483 33507 18514 33541
rect 18418 33449 18514 33507
rect 18613 33546 18659 33558
rect 18613 33512 18619 33546
rect 18653 33512 18659 33546
rect 18613 33500 18659 33512
rect 18962 33541 19058 33599
rect 18962 33507 18993 33541
rect 19027 33507 19058 33541
rect 18418 33415 18449 33449
rect 18483 33415 18514 33449
rect 18418 33386 18514 33415
rect 18715 33456 18861 33477
rect 18715 33420 18748 33456
rect 18784 33420 18861 33456
rect 18715 33278 18861 33420
rect 18962 33449 19058 33507
rect 18962 33415 18993 33449
rect 19027 33415 19058 33449
rect 18962 33386 19058 33415
rect 18714 33216 18861 33278
rect 18426 32891 18522 32920
rect 18426 32857 18457 32891
rect 18491 32857 18522 32891
rect 18426 32799 18522 32857
rect 18714 32820 18784 33216
rect 18426 32765 18457 32799
rect 18491 32765 18522 32799
rect 18426 32707 18522 32765
rect 18640 32800 18784 32820
rect 18970 32891 19066 32920
rect 18970 32857 19001 32891
rect 19035 32857 19066 32891
rect 18640 32764 18672 32800
rect 18706 32764 18875 32800
rect 18640 32746 18875 32764
rect 18640 32744 18744 32746
rect 18426 32673 18457 32707
rect 18491 32673 18522 32707
rect 18426 32615 18522 32673
rect 18426 32581 18457 32615
rect 18491 32581 18522 32615
rect 18426 32523 18522 32581
rect 18426 32489 18457 32523
rect 18491 32489 18522 32523
rect 18426 32431 18522 32489
rect 18426 32397 18457 32431
rect 18491 32397 18522 32431
rect 18426 32339 18522 32397
rect 18426 32305 18457 32339
rect 18491 32305 18522 32339
rect 18426 32247 18522 32305
rect 18426 32213 18457 32247
rect 18491 32213 18522 32247
rect 18426 32155 18522 32213
rect 18426 32148 18457 32155
rect 18491 32148 18522 32155
rect 18426 32066 18432 32148
rect 18512 32066 18522 32148
rect 18426 32063 18522 32066
rect 18426 32029 18457 32063
rect 18491 32029 18522 32063
rect 18426 31971 18522 32029
rect 18689 32061 18735 32073
rect 18689 32027 18695 32061
rect 18729 32027 18735 32061
rect 18689 32015 18735 32027
rect 18426 31937 18457 31971
rect 18491 31937 18522 31971
rect 18426 31879 18522 31937
rect 18621 31974 18667 31986
rect 18621 31940 18627 31974
rect 18661 31940 18667 31974
rect 18621 31928 18667 31940
rect 18426 31845 18457 31879
rect 18491 31845 18522 31879
rect 18426 31787 18522 31845
rect 18426 31753 18457 31787
rect 18491 31753 18522 31787
rect 18426 31695 18522 31753
rect 18426 31661 18457 31695
rect 18491 31661 18522 31695
rect 18630 31672 18658 31928
rect 18426 31603 18522 31661
rect 18621 31660 18667 31672
rect 18621 31626 18627 31660
rect 18661 31626 18667 31660
rect 18621 31614 18667 31626
rect 18426 31569 18457 31603
rect 18491 31569 18522 31603
rect 18426 31511 18522 31569
rect 18426 31477 18457 31511
rect 18491 31477 18522 31511
rect 18426 31419 18522 31477
rect 18426 31385 18457 31419
rect 18491 31385 18522 31419
rect 18426 31327 18522 31385
rect 18426 31293 18457 31327
rect 18491 31293 18522 31327
rect 18426 31235 18522 31293
rect 18630 31252 18658 31614
rect 18698 31569 18726 32015
rect 18689 31557 18735 31569
rect 18689 31523 18695 31557
rect 18729 31523 18735 31557
rect 18689 31511 18735 31523
rect 18698 31331 18726 31511
rect 18804 31400 18875 32746
rect 18804 31364 18824 31400
rect 18860 31364 18875 31400
rect 18804 31354 18875 31364
rect 18970 32799 19066 32857
rect 18970 32765 19001 32799
rect 19035 32765 19066 32799
rect 18970 32707 19066 32765
rect 18970 32673 19001 32707
rect 19035 32673 19066 32707
rect 18970 32615 19066 32673
rect 18970 32581 19001 32615
rect 19035 32581 19066 32615
rect 18970 32523 19066 32581
rect 18970 32489 19001 32523
rect 19035 32489 19066 32523
rect 18970 32431 19066 32489
rect 18970 32397 19001 32431
rect 19035 32397 19066 32431
rect 18970 32339 19066 32397
rect 18970 32305 19001 32339
rect 19035 32305 19066 32339
rect 18970 32247 19066 32305
rect 18970 32213 19001 32247
rect 19035 32213 19066 32247
rect 18970 32155 19066 32213
rect 18970 32152 19001 32155
rect 19035 32152 19066 32155
rect 18970 32070 18980 32152
rect 19060 32070 19066 32152
rect 18970 32063 19066 32070
rect 18970 32029 19001 32063
rect 19035 32029 19066 32063
rect 18970 31971 19066 32029
rect 18970 31937 19001 31971
rect 19035 31937 19066 31971
rect 18970 31879 19066 31937
rect 18970 31845 19001 31879
rect 19035 31845 19066 31879
rect 18970 31787 19066 31845
rect 18970 31753 19001 31787
rect 19035 31753 19066 31787
rect 18970 31695 19066 31753
rect 18970 31661 19001 31695
rect 19035 31661 19066 31695
rect 18970 31603 19066 31661
rect 18970 31569 19001 31603
rect 19035 31569 19066 31603
rect 18970 31511 19066 31569
rect 18970 31477 19001 31511
rect 19035 31477 19066 31511
rect 18970 31419 19066 31477
rect 18970 31385 19001 31419
rect 19035 31385 19066 31419
rect 18689 31319 18735 31331
rect 18689 31285 18695 31319
rect 18729 31285 18735 31319
rect 18689 31273 18735 31285
rect 18970 31327 19066 31385
rect 18970 31293 19001 31327
rect 19035 31293 19066 31327
rect 18426 31201 18457 31235
rect 18491 31201 18522 31235
rect 18426 31143 18522 31201
rect 18621 31240 18667 31252
rect 18621 31206 18627 31240
rect 18661 31206 18667 31240
rect 18621 31194 18667 31206
rect 18970 31235 19066 31293
rect 18970 31201 19001 31235
rect 19035 31201 19066 31235
rect 18426 31109 18457 31143
rect 18491 31109 18522 31143
rect 18426 31080 18522 31109
rect 18723 31150 18869 31171
rect 18723 31114 18756 31150
rect 18792 31114 18869 31150
rect 18723 30882 18869 31114
rect 18970 31143 19066 31201
rect 18970 31109 19001 31143
rect 19035 31109 19066 31143
rect 18970 31080 19066 31109
rect 18720 30778 18869 30882
rect 18434 30677 18530 30706
rect 18434 30643 18465 30677
rect 18499 30643 18530 30677
rect 18434 30585 18530 30643
rect 18720 30606 18754 30778
rect 18434 30551 18465 30585
rect 18499 30551 18530 30585
rect 18434 30493 18530 30551
rect 18648 30586 18754 30606
rect 18978 30677 19074 30706
rect 18978 30643 19009 30677
rect 19043 30643 19074 30677
rect 18648 30550 18680 30586
rect 18714 30582 18754 30586
rect 18812 30582 18883 30586
rect 18714 30550 18883 30582
rect 18648 30532 18883 30550
rect 18648 30530 18752 30532
rect 18434 30459 18465 30493
rect 18499 30459 18530 30493
rect 18434 30401 18530 30459
rect 18434 30367 18465 30401
rect 18499 30367 18530 30401
rect 18434 30309 18530 30367
rect 18434 30275 18465 30309
rect 18499 30275 18530 30309
rect 18434 30217 18530 30275
rect 18434 30183 18465 30217
rect 18499 30183 18530 30217
rect 18434 30125 18530 30183
rect 18434 30091 18465 30125
rect 18499 30091 18530 30125
rect 18434 30033 18530 30091
rect 18434 29999 18465 30033
rect 18499 29999 18530 30033
rect 18434 29941 18530 29999
rect 18434 29934 18465 29941
rect 18499 29934 18530 29941
rect 18434 29852 18440 29934
rect 18520 29852 18530 29934
rect 18434 29849 18530 29852
rect 18434 29815 18465 29849
rect 18499 29815 18530 29849
rect 18434 29757 18530 29815
rect 18697 29847 18743 29859
rect 18697 29813 18703 29847
rect 18737 29813 18743 29847
rect 18697 29801 18743 29813
rect 18434 29723 18465 29757
rect 18499 29723 18530 29757
rect 18434 29665 18530 29723
rect 18629 29760 18675 29772
rect 18629 29726 18635 29760
rect 18669 29726 18675 29760
rect 18629 29714 18675 29726
rect 18434 29631 18465 29665
rect 18499 29631 18530 29665
rect 18434 29573 18530 29631
rect 18434 29539 18465 29573
rect 18499 29539 18530 29573
rect 18434 29481 18530 29539
rect 18434 29447 18465 29481
rect 18499 29447 18530 29481
rect 18638 29458 18666 29714
rect 18434 29389 18530 29447
rect 18629 29446 18675 29458
rect 18629 29412 18635 29446
rect 18669 29412 18675 29446
rect 18629 29400 18675 29412
rect 18434 29355 18465 29389
rect 18499 29355 18530 29389
rect 18434 29297 18530 29355
rect 18434 29263 18465 29297
rect 18499 29263 18530 29297
rect 18434 29205 18530 29263
rect 18434 29171 18465 29205
rect 18499 29171 18530 29205
rect 18434 29113 18530 29171
rect 18434 29079 18465 29113
rect 18499 29079 18530 29113
rect 18434 29021 18530 29079
rect 18638 29038 18666 29400
rect 18706 29355 18734 29801
rect 18697 29343 18743 29355
rect 18697 29309 18703 29343
rect 18737 29309 18743 29343
rect 18697 29297 18743 29309
rect 18706 29117 18734 29297
rect 18812 29186 18883 30532
rect 18812 29150 18832 29186
rect 18868 29150 18883 29186
rect 18812 29140 18883 29150
rect 18978 30585 19074 30643
rect 18978 30551 19009 30585
rect 19043 30551 19074 30585
rect 18978 30493 19074 30551
rect 18978 30459 19009 30493
rect 19043 30459 19074 30493
rect 18978 30401 19074 30459
rect 18978 30367 19009 30401
rect 19043 30367 19074 30401
rect 18978 30309 19074 30367
rect 18978 30275 19009 30309
rect 19043 30275 19074 30309
rect 18978 30217 19074 30275
rect 18978 30183 19009 30217
rect 19043 30183 19074 30217
rect 18978 30125 19074 30183
rect 18978 30091 19009 30125
rect 19043 30091 19074 30125
rect 18978 30033 19074 30091
rect 18978 29999 19009 30033
rect 19043 29999 19074 30033
rect 18978 29941 19074 29999
rect 18978 29938 19009 29941
rect 19043 29938 19074 29941
rect 18978 29856 18988 29938
rect 19068 29856 19074 29938
rect 18978 29849 19074 29856
rect 18978 29815 19009 29849
rect 19043 29815 19074 29849
rect 18978 29757 19074 29815
rect 18978 29723 19009 29757
rect 19043 29723 19074 29757
rect 18978 29665 19074 29723
rect 18978 29631 19009 29665
rect 19043 29631 19074 29665
rect 18978 29573 19074 29631
rect 18978 29539 19009 29573
rect 19043 29539 19074 29573
rect 18978 29481 19074 29539
rect 18978 29447 19009 29481
rect 19043 29447 19074 29481
rect 18978 29389 19074 29447
rect 18978 29355 19009 29389
rect 19043 29355 19074 29389
rect 18978 29297 19074 29355
rect 18978 29263 19009 29297
rect 19043 29263 19074 29297
rect 18978 29205 19074 29263
rect 18978 29171 19009 29205
rect 19043 29171 19074 29205
rect 18697 29105 18743 29117
rect 18697 29071 18703 29105
rect 18737 29071 18743 29105
rect 18697 29059 18743 29071
rect 18978 29113 19074 29171
rect 18978 29079 19009 29113
rect 19043 29079 19074 29113
rect 18434 28987 18465 29021
rect 18499 28987 18530 29021
rect 18434 28929 18530 28987
rect 18629 29026 18675 29038
rect 18629 28992 18635 29026
rect 18669 28992 18675 29026
rect 18629 28980 18675 28992
rect 18978 29021 19074 29079
rect 18978 28987 19009 29021
rect 19043 28987 19074 29021
rect 18434 28895 18465 28929
rect 18499 28895 18530 28929
rect 18434 28866 18530 28895
rect 18731 28936 18877 28957
rect 18731 28900 18764 28936
rect 18800 28900 18877 28936
rect 18731 28742 18877 28900
rect 18978 28929 19074 28987
rect 18978 28895 19009 28929
rect 19043 28895 19074 28929
rect 18978 28866 19074 28895
rect 18730 28608 18877 28742
rect 18416 28477 18512 28506
rect 18416 28443 18447 28477
rect 18481 28443 18512 28477
rect 18416 28385 18512 28443
rect 18730 28406 18766 28608
rect 18416 28351 18447 28385
rect 18481 28351 18512 28385
rect 18416 28293 18512 28351
rect 18630 28386 18766 28406
rect 18960 28477 19056 28506
rect 18960 28443 18991 28477
rect 19025 28443 19056 28477
rect 18630 28350 18662 28386
rect 18696 28382 18766 28386
rect 18794 28382 18865 28386
rect 18696 28350 18865 28382
rect 18630 28332 18865 28350
rect 18630 28330 18734 28332
rect 18416 28259 18447 28293
rect 18481 28259 18512 28293
rect 18416 28201 18512 28259
rect 18416 28167 18447 28201
rect 18481 28167 18512 28201
rect 18416 28109 18512 28167
rect 18416 28075 18447 28109
rect 18481 28075 18512 28109
rect 18416 28017 18512 28075
rect 18416 27983 18447 28017
rect 18481 27983 18512 28017
rect 18416 27925 18512 27983
rect 18416 27891 18447 27925
rect 18481 27891 18512 27925
rect 18416 27833 18512 27891
rect 18416 27799 18447 27833
rect 18481 27799 18512 27833
rect 18416 27741 18512 27799
rect 18416 27734 18447 27741
rect 18481 27734 18512 27741
rect 18416 27652 18422 27734
rect 18502 27652 18512 27734
rect 18416 27649 18512 27652
rect 18416 27615 18447 27649
rect 18481 27615 18512 27649
rect 18416 27557 18512 27615
rect 18679 27647 18725 27659
rect 18679 27613 18685 27647
rect 18719 27613 18725 27647
rect 18679 27601 18725 27613
rect 18416 27523 18447 27557
rect 18481 27523 18512 27557
rect 18416 27465 18512 27523
rect 18611 27560 18657 27572
rect 18611 27526 18617 27560
rect 18651 27526 18657 27560
rect 18611 27514 18657 27526
rect 18416 27431 18447 27465
rect 18481 27431 18512 27465
rect 18416 27373 18512 27431
rect 18416 27339 18447 27373
rect 18481 27339 18512 27373
rect 18416 27281 18512 27339
rect 18416 27247 18447 27281
rect 18481 27247 18512 27281
rect 18620 27258 18648 27514
rect 18416 27189 18512 27247
rect 18611 27246 18657 27258
rect 18611 27212 18617 27246
rect 18651 27212 18657 27246
rect 18611 27200 18657 27212
rect 18416 27155 18447 27189
rect 18481 27155 18512 27189
rect 18416 27097 18512 27155
rect 18416 27063 18447 27097
rect 18481 27063 18512 27097
rect 18416 27005 18512 27063
rect 18416 26971 18447 27005
rect 18481 26971 18512 27005
rect 18416 26913 18512 26971
rect 18416 26879 18447 26913
rect 18481 26879 18512 26913
rect 18416 26821 18512 26879
rect 18620 26838 18648 27200
rect 18688 27155 18716 27601
rect 18679 27143 18725 27155
rect 18679 27109 18685 27143
rect 18719 27109 18725 27143
rect 18679 27097 18725 27109
rect 18688 26917 18716 27097
rect 18794 26986 18865 28332
rect 18794 26950 18814 26986
rect 18850 26950 18865 26986
rect 18794 26940 18865 26950
rect 18960 28385 19056 28443
rect 18960 28351 18991 28385
rect 19025 28351 19056 28385
rect 18960 28293 19056 28351
rect 18960 28259 18991 28293
rect 19025 28259 19056 28293
rect 18960 28201 19056 28259
rect 18960 28167 18991 28201
rect 19025 28167 19056 28201
rect 18960 28109 19056 28167
rect 18960 28075 18991 28109
rect 19025 28075 19056 28109
rect 18960 28017 19056 28075
rect 18960 27983 18991 28017
rect 19025 27983 19056 28017
rect 18960 27925 19056 27983
rect 18960 27891 18991 27925
rect 19025 27891 19056 27925
rect 18960 27833 19056 27891
rect 18960 27799 18991 27833
rect 19025 27799 19056 27833
rect 18960 27741 19056 27799
rect 18960 27738 18991 27741
rect 19025 27738 19056 27741
rect 18960 27656 18970 27738
rect 19050 27656 19056 27738
rect 18960 27649 19056 27656
rect 18960 27615 18991 27649
rect 19025 27615 19056 27649
rect 18960 27557 19056 27615
rect 18960 27523 18991 27557
rect 19025 27523 19056 27557
rect 18960 27465 19056 27523
rect 18960 27431 18991 27465
rect 19025 27431 19056 27465
rect 18960 27373 19056 27431
rect 18960 27339 18991 27373
rect 19025 27339 19056 27373
rect 18960 27281 19056 27339
rect 18960 27247 18991 27281
rect 19025 27247 19056 27281
rect 18960 27189 19056 27247
rect 18960 27155 18991 27189
rect 19025 27155 19056 27189
rect 18960 27097 19056 27155
rect 18960 27063 18991 27097
rect 19025 27063 19056 27097
rect 18960 27005 19056 27063
rect 18960 26971 18991 27005
rect 19025 26971 19056 27005
rect 18679 26905 18725 26917
rect 18679 26871 18685 26905
rect 18719 26871 18725 26905
rect 18679 26859 18725 26871
rect 18960 26913 19056 26971
rect 18960 26879 18991 26913
rect 19025 26879 19056 26913
rect 18416 26787 18447 26821
rect 18481 26787 18512 26821
rect 18416 26729 18512 26787
rect 18611 26826 18657 26838
rect 18611 26792 18617 26826
rect 18651 26792 18657 26826
rect 18611 26780 18657 26792
rect 18960 26821 19056 26879
rect 18960 26787 18991 26821
rect 19025 26787 19056 26821
rect 18416 26695 18447 26729
rect 18481 26695 18512 26729
rect 18416 26666 18512 26695
rect 18713 26736 18859 26757
rect 18713 26700 18746 26736
rect 18782 26700 18859 26736
rect 18713 26468 18859 26700
rect 18960 26729 19056 26787
rect 18960 26695 18991 26729
rect 19025 26695 19056 26729
rect 18960 26666 19056 26695
rect 18710 26364 18859 26468
rect 18424 26263 18520 26292
rect 18424 26229 18455 26263
rect 18489 26229 18520 26263
rect 18424 26171 18520 26229
rect 18710 26192 18744 26364
rect 18424 26137 18455 26171
rect 18489 26137 18520 26171
rect 18424 26079 18520 26137
rect 18638 26172 18744 26192
rect 18968 26263 19064 26292
rect 18968 26229 18999 26263
rect 19033 26229 19064 26263
rect 18638 26136 18670 26172
rect 18704 26168 18744 26172
rect 18802 26168 18873 26172
rect 18704 26136 18873 26168
rect 18638 26118 18873 26136
rect 18638 26116 18742 26118
rect 18424 26045 18455 26079
rect 18489 26045 18520 26079
rect 18424 25987 18520 26045
rect 18424 25953 18455 25987
rect 18489 25953 18520 25987
rect 18424 25895 18520 25953
rect 18424 25861 18455 25895
rect 18489 25861 18520 25895
rect 18424 25803 18520 25861
rect 18424 25769 18455 25803
rect 18489 25769 18520 25803
rect 18424 25711 18520 25769
rect 18424 25677 18455 25711
rect 18489 25677 18520 25711
rect 18424 25619 18520 25677
rect 18424 25585 18455 25619
rect 18489 25585 18520 25619
rect 18424 25527 18520 25585
rect 18424 25520 18455 25527
rect 18489 25520 18520 25527
rect 18424 25438 18430 25520
rect 18510 25438 18520 25520
rect 18424 25435 18520 25438
rect 18424 25401 18455 25435
rect 18489 25401 18520 25435
rect 18424 25343 18520 25401
rect 18687 25433 18733 25445
rect 18687 25399 18693 25433
rect 18727 25399 18733 25433
rect 18687 25387 18733 25399
rect 18424 25309 18455 25343
rect 18489 25309 18520 25343
rect 18424 25251 18520 25309
rect 18619 25346 18665 25358
rect 18619 25312 18625 25346
rect 18659 25312 18665 25346
rect 18619 25300 18665 25312
rect 18424 25217 18455 25251
rect 18489 25217 18520 25251
rect 18424 25159 18520 25217
rect 18424 25125 18455 25159
rect 18489 25125 18520 25159
rect 18424 25067 18520 25125
rect 18424 25033 18455 25067
rect 18489 25033 18520 25067
rect 18628 25044 18656 25300
rect 18424 24975 18520 25033
rect 18619 25032 18665 25044
rect 18619 24998 18625 25032
rect 18659 24998 18665 25032
rect 18619 24986 18665 24998
rect 18424 24941 18455 24975
rect 18489 24941 18520 24975
rect 18424 24883 18520 24941
rect 18424 24849 18455 24883
rect 18489 24849 18520 24883
rect 18424 24791 18520 24849
rect 18424 24757 18455 24791
rect 18489 24757 18520 24791
rect 18424 24699 18520 24757
rect 18424 24665 18455 24699
rect 18489 24665 18520 24699
rect 18424 24607 18520 24665
rect 18628 24624 18656 24986
rect 18696 24941 18724 25387
rect 18687 24929 18733 24941
rect 18687 24895 18693 24929
rect 18727 24895 18733 24929
rect 18687 24883 18733 24895
rect 18696 24703 18724 24883
rect 18802 24772 18873 26118
rect 18802 24736 18822 24772
rect 18858 24736 18873 24772
rect 18802 24726 18873 24736
rect 18968 26171 19064 26229
rect 18968 26137 18999 26171
rect 19033 26137 19064 26171
rect 18968 26079 19064 26137
rect 18968 26045 18999 26079
rect 19033 26045 19064 26079
rect 18968 25987 19064 26045
rect 18968 25953 18999 25987
rect 19033 25953 19064 25987
rect 18968 25895 19064 25953
rect 18968 25861 18999 25895
rect 19033 25861 19064 25895
rect 18968 25803 19064 25861
rect 18968 25769 18999 25803
rect 19033 25769 19064 25803
rect 18968 25711 19064 25769
rect 18968 25677 18999 25711
rect 19033 25677 19064 25711
rect 18968 25619 19064 25677
rect 18968 25585 18999 25619
rect 19033 25585 19064 25619
rect 18968 25527 19064 25585
rect 18968 25524 18999 25527
rect 19033 25524 19064 25527
rect 18968 25442 18978 25524
rect 19058 25442 19064 25524
rect 18968 25435 19064 25442
rect 18968 25401 18999 25435
rect 19033 25401 19064 25435
rect 18968 25343 19064 25401
rect 18968 25309 18999 25343
rect 19033 25309 19064 25343
rect 18968 25251 19064 25309
rect 18968 25217 18999 25251
rect 19033 25217 19064 25251
rect 18968 25159 19064 25217
rect 18968 25125 18999 25159
rect 19033 25125 19064 25159
rect 18968 25067 19064 25125
rect 18968 25033 18999 25067
rect 19033 25033 19064 25067
rect 18968 24975 19064 25033
rect 18968 24941 18999 24975
rect 19033 24941 19064 24975
rect 18968 24883 19064 24941
rect 18968 24849 18999 24883
rect 19033 24849 19064 24883
rect 18968 24791 19064 24849
rect 18968 24757 18999 24791
rect 19033 24757 19064 24791
rect 18687 24691 18733 24703
rect 18687 24657 18693 24691
rect 18727 24657 18733 24691
rect 18687 24645 18733 24657
rect 18968 24699 19064 24757
rect 18968 24665 18999 24699
rect 19033 24665 19064 24699
rect 18424 24573 18455 24607
rect 18489 24573 18520 24607
rect 18424 24515 18520 24573
rect 18619 24612 18665 24624
rect 18619 24578 18625 24612
rect 18659 24578 18665 24612
rect 18619 24566 18665 24578
rect 18968 24607 19064 24665
rect 18968 24573 18999 24607
rect 19033 24573 19064 24607
rect 18424 24481 18455 24515
rect 18489 24481 18520 24515
rect 18424 24452 18520 24481
rect 18721 24522 18867 24543
rect 18721 24486 18754 24522
rect 18790 24486 18867 24522
rect 18721 24342 18867 24486
rect 18968 24515 19064 24573
rect 18968 24481 18999 24515
rect 19033 24481 19064 24515
rect 18968 24452 19064 24481
rect 9760 23438 11600 23444
rect 7546 23430 9386 23436
rect 7546 23405 8532 23430
rect 8614 23405 9386 23430
rect 7546 23371 7575 23405
rect 7609 23371 7667 23405
rect 7701 23371 7759 23405
rect 7793 23371 7851 23405
rect 7885 23371 7943 23405
rect 7977 23371 8035 23405
rect 8069 23371 8127 23405
rect 8161 23371 8219 23405
rect 8253 23371 8311 23405
rect 8345 23371 8403 23405
rect 8437 23371 8495 23405
rect 8529 23371 8532 23405
rect 8621 23371 8679 23405
rect 8713 23371 8771 23405
rect 8805 23371 8863 23405
rect 8897 23371 8955 23405
rect 8989 23371 9047 23405
rect 9081 23371 9139 23405
rect 9173 23371 9231 23405
rect 9265 23371 9323 23405
rect 9357 23371 9386 23405
rect 7546 23350 8532 23371
rect 8614 23350 9386 23371
rect 7546 23340 9386 23350
rect 9760 23413 10746 23438
rect 10828 23413 11600 23438
rect 16480 23436 18320 23442
rect 14174 23428 16014 23434
rect 9760 23379 9789 23413
rect 9823 23379 9881 23413
rect 9915 23379 9973 23413
rect 10007 23379 10065 23413
rect 10099 23379 10157 23413
rect 10191 23379 10249 23413
rect 10283 23379 10341 23413
rect 10375 23379 10433 23413
rect 10467 23379 10525 23413
rect 10559 23379 10617 23413
rect 10651 23379 10709 23413
rect 10743 23379 10746 23413
rect 10835 23379 10893 23413
rect 10927 23379 10985 23413
rect 11019 23379 11077 23413
rect 11111 23379 11169 23413
rect 11203 23379 11261 23413
rect 11295 23379 11353 23413
rect 11387 23379 11445 23413
rect 11479 23379 11537 23413
rect 11571 23379 11600 23413
rect 9760 23358 10746 23379
rect 10828 23358 11600 23379
rect 9760 23348 11600 23358
rect 11960 23420 13800 23426
rect 11960 23395 12946 23420
rect 13028 23395 13800 23420
rect 11960 23361 11989 23395
rect 12023 23361 12081 23395
rect 12115 23361 12173 23395
rect 12207 23361 12265 23395
rect 12299 23361 12357 23395
rect 12391 23361 12449 23395
rect 12483 23361 12541 23395
rect 12575 23361 12633 23395
rect 12667 23361 12725 23395
rect 12759 23361 12817 23395
rect 12851 23361 12909 23395
rect 12943 23361 12946 23395
rect 13035 23361 13093 23395
rect 13127 23361 13185 23395
rect 13219 23361 13277 23395
rect 13311 23361 13369 23395
rect 13403 23361 13461 23395
rect 13495 23361 13553 23395
rect 13587 23361 13645 23395
rect 13679 23361 13737 23395
rect 13771 23361 13800 23395
rect 11960 23340 12946 23361
rect 13028 23340 13800 23361
rect 11960 23330 13800 23340
rect 14174 23403 15160 23428
rect 15242 23403 16014 23428
rect 14174 23369 14203 23403
rect 14237 23369 14295 23403
rect 14329 23369 14387 23403
rect 14421 23369 14479 23403
rect 14513 23369 14571 23403
rect 14605 23369 14663 23403
rect 14697 23369 14755 23403
rect 14789 23369 14847 23403
rect 14881 23369 14939 23403
rect 14973 23369 15031 23403
rect 15065 23369 15123 23403
rect 15157 23369 15160 23403
rect 15249 23369 15307 23403
rect 15341 23369 15399 23403
rect 15433 23369 15491 23403
rect 15525 23369 15583 23403
rect 15617 23369 15675 23403
rect 15709 23369 15767 23403
rect 15801 23369 15859 23403
rect 15893 23369 15951 23403
rect 15985 23369 16014 23403
rect 14174 23348 15160 23369
rect 15242 23348 16014 23369
rect 14174 23338 16014 23348
rect 16480 23411 17466 23436
rect 17548 23411 18320 23436
rect 16480 23377 16509 23411
rect 16543 23377 16601 23411
rect 16635 23377 16693 23411
rect 16727 23377 16785 23411
rect 16819 23377 16877 23411
rect 16911 23377 16969 23411
rect 17003 23377 17061 23411
rect 17095 23377 17153 23411
rect 17187 23377 17245 23411
rect 17279 23377 17337 23411
rect 17371 23377 17429 23411
rect 17463 23377 17466 23411
rect 17555 23377 17613 23411
rect 17647 23377 17705 23411
rect 17739 23377 17797 23411
rect 17831 23377 17889 23411
rect 17923 23377 17981 23411
rect 18015 23377 18073 23411
rect 18107 23377 18165 23411
rect 18199 23377 18257 23411
rect 18291 23377 18320 23411
rect 16480 23356 17466 23377
rect 17548 23356 18320 23377
rect 16480 23346 18320 23356
rect 9874 23243 9932 23249
rect 7660 23235 7718 23241
rect 7660 23201 7672 23235
rect 7706 23232 7718 23235
rect 8080 23235 8138 23241
rect 8080 23232 8092 23235
rect 7706 23204 8092 23232
rect 7706 23201 7718 23204
rect 7660 23195 7718 23201
rect 8080 23201 8092 23204
rect 8126 23232 8138 23235
rect 8394 23235 8452 23241
rect 8394 23232 8406 23235
rect 8126 23204 8406 23232
rect 8126 23201 8138 23204
rect 8080 23195 8138 23201
rect 8394 23201 8406 23204
rect 8440 23201 8452 23235
rect 8394 23195 8452 23201
rect 9210 23190 9286 23222
rect 9874 23209 9886 23243
rect 9920 23240 9932 23243
rect 10294 23243 10352 23249
rect 10294 23240 10306 23243
rect 9920 23212 10306 23240
rect 9920 23209 9932 23212
rect 9874 23203 9932 23209
rect 10294 23209 10306 23212
rect 10340 23240 10352 23243
rect 10608 23243 10666 23249
rect 10608 23240 10620 23243
rect 10340 23212 10620 23240
rect 10340 23209 10352 23212
rect 10294 23203 10352 23209
rect 10608 23209 10620 23212
rect 10654 23209 10666 23243
rect 16594 23241 16652 23247
rect 14288 23233 14346 23239
rect 10608 23203 10666 23209
rect 7739 23167 7797 23173
rect 6269 23106 7637 23139
rect 7739 23133 7751 23167
rect 7785 23164 7797 23167
rect 7977 23167 8035 23173
rect 7977 23164 7989 23167
rect 7785 23136 7989 23164
rect 7785 23133 7797 23136
rect 7739 23127 7797 23133
rect 7977 23133 7989 23136
rect 8023 23164 8035 23167
rect 8481 23167 8539 23173
rect 8481 23164 8493 23167
rect 8023 23136 8493 23164
rect 8023 23133 8035 23136
rect 7977 23127 8035 23133
rect 8481 23133 8493 23136
rect 8527 23133 8539 23167
rect 8481 23127 8539 23133
rect 9210 23156 9230 23190
rect 9266 23156 9286 23190
rect 11424 23198 11500 23230
rect 9210 23150 9286 23156
rect 9953 23175 10011 23181
rect 9210 23147 9562 23150
rect 9210 23118 9851 23147
rect 9953 23141 9965 23175
rect 9999 23172 10011 23175
rect 10191 23175 10249 23181
rect 10191 23172 10203 23175
rect 9999 23144 10203 23172
rect 9999 23141 10011 23144
rect 9953 23135 10011 23141
rect 10191 23141 10203 23144
rect 10237 23172 10249 23175
rect 10695 23175 10753 23181
rect 10695 23172 10707 23175
rect 10237 23144 10707 23172
rect 10237 23141 10249 23144
rect 10191 23135 10249 23141
rect 10695 23141 10707 23144
rect 10741 23141 10753 23175
rect 10695 23135 10753 23141
rect 11424 23164 11444 23198
rect 11480 23164 11500 23198
rect 12074 23225 12132 23231
rect 12074 23191 12086 23225
rect 12120 23222 12132 23225
rect 12494 23225 12552 23231
rect 12494 23222 12506 23225
rect 12120 23194 12506 23222
rect 12120 23191 12132 23194
rect 12074 23185 12132 23191
rect 12494 23191 12506 23194
rect 12540 23222 12552 23225
rect 12808 23225 12866 23231
rect 12808 23222 12820 23225
rect 12540 23194 12820 23222
rect 12540 23191 12552 23194
rect 12494 23185 12552 23191
rect 12808 23191 12820 23194
rect 12854 23191 12866 23225
rect 12808 23185 12866 23191
rect 11424 23130 11500 23164
rect 13624 23180 13700 23212
rect 14288 23199 14300 23233
rect 14334 23230 14346 23233
rect 14708 23233 14766 23239
rect 14708 23230 14720 23233
rect 14334 23202 14720 23230
rect 14334 23199 14346 23202
rect 14288 23193 14346 23199
rect 14708 23199 14720 23202
rect 14754 23230 14766 23233
rect 15022 23233 15080 23239
rect 15022 23230 15034 23233
rect 14754 23202 15034 23230
rect 14754 23199 14766 23202
rect 14708 23193 14766 23199
rect 15022 23199 15034 23202
rect 15068 23199 15080 23233
rect 15022 23193 15080 23199
rect 12153 23157 12211 23163
rect 11424 23129 11836 23130
rect 11424 23126 12051 23129
rect 6269 23070 7580 23106
rect 7616 23070 7637 23106
rect 6269 22993 7637 23070
rect 9212 23116 9851 23118
rect 9212 23058 9262 23116
rect 9458 23114 9851 23116
rect 9458 23078 9794 23114
rect 9830 23078 9851 23114
rect 7820 23038 9266 23058
rect 7820 23002 7830 23038
rect 7866 23002 9266 23038
rect 6269 18485 6415 22993
rect 7820 22987 9266 23002
rect 9458 23001 9851 23078
rect 11426 23096 12051 23126
rect 12153 23123 12165 23157
rect 12199 23154 12211 23157
rect 12391 23157 12449 23163
rect 12391 23154 12403 23157
rect 12199 23126 12403 23154
rect 12199 23123 12211 23126
rect 12153 23117 12211 23123
rect 12391 23123 12403 23126
rect 12437 23154 12449 23157
rect 12895 23157 12953 23163
rect 12895 23154 12907 23157
rect 12437 23126 12907 23154
rect 12437 23123 12449 23126
rect 12391 23117 12449 23123
rect 12895 23123 12907 23126
rect 12941 23123 12953 23157
rect 12895 23117 12953 23123
rect 13624 23146 13644 23180
rect 13680 23146 13700 23180
rect 15838 23188 15914 23220
rect 16594 23207 16606 23241
rect 16640 23238 16652 23241
rect 17014 23241 17072 23247
rect 17014 23238 17026 23241
rect 16640 23210 17026 23238
rect 16640 23207 16652 23210
rect 16594 23201 16652 23207
rect 17014 23207 17026 23210
rect 17060 23238 17072 23241
rect 17328 23241 17386 23247
rect 17328 23238 17340 23241
rect 17060 23210 17340 23238
rect 17060 23207 17072 23210
rect 17014 23201 17072 23207
rect 17328 23207 17340 23210
rect 17374 23207 17386 23241
rect 17328 23201 17386 23207
rect 13624 23140 13700 23146
rect 14367 23165 14425 23171
rect 13624 23137 13976 23140
rect 13624 23108 14265 23137
rect 14367 23131 14379 23165
rect 14413 23162 14425 23165
rect 14605 23165 14663 23171
rect 14605 23162 14617 23165
rect 14413 23134 14617 23162
rect 14413 23131 14425 23134
rect 14367 23125 14425 23131
rect 14605 23131 14617 23134
rect 14651 23162 14663 23165
rect 15109 23165 15167 23171
rect 15109 23162 15121 23165
rect 14651 23134 15121 23162
rect 14651 23131 14663 23134
rect 14605 23125 14663 23131
rect 15109 23131 15121 23134
rect 15155 23131 15167 23165
rect 15109 23125 15167 23131
rect 15838 23154 15858 23188
rect 15894 23154 15914 23188
rect 18144 23196 18220 23228
rect 15838 23146 15914 23154
rect 16673 23173 16731 23179
rect 15838 23145 16372 23146
rect 15838 23116 16571 23145
rect 16673 23139 16685 23173
rect 16719 23170 16731 23173
rect 16911 23173 16969 23179
rect 16911 23170 16923 23173
rect 16719 23142 16923 23170
rect 16719 23139 16731 23142
rect 16673 23133 16731 23139
rect 16911 23139 16923 23142
rect 16957 23170 16969 23173
rect 17415 23173 17473 23179
rect 18144 23174 18164 23196
rect 17415 23170 17427 23173
rect 16957 23142 17427 23170
rect 16957 23139 16969 23142
rect 16911 23133 16969 23139
rect 17415 23139 17427 23142
rect 17461 23139 17473 23173
rect 17415 23133 17473 23139
rect 18140 23162 18164 23174
rect 18200 23174 18220 23196
rect 18723 23174 18867 24342
rect 18200 23162 18867 23174
rect 11426 23094 11994 23096
rect 11426 23066 11476 23094
rect 10034 23046 11480 23066
rect 10034 23010 10044 23046
rect 10080 23010 11480 23046
rect 10034 22995 11480 23010
rect 11702 23060 11994 23094
rect 12030 23060 12051 23096
rect 11702 22983 12051 23060
rect 13626 23106 14265 23108
rect 13626 23048 13676 23106
rect 13872 23104 14265 23106
rect 13872 23068 14208 23104
rect 14244 23068 14265 23104
rect 12234 23028 13680 23048
rect 12234 22992 12244 23028
rect 12280 22992 13680 23028
rect 12234 22977 13680 22992
rect 13872 22991 14265 23068
rect 15840 23112 16571 23116
rect 15840 23076 16514 23112
rect 16550 23076 16571 23112
rect 15840 23056 15894 23076
rect 14448 23036 15894 23056
rect 14448 23000 14458 23036
rect 14494 23000 15894 23036
rect 14448 22985 15894 23000
rect 16310 22999 16571 23076
rect 18140 23064 18867 23162
rect 16754 23044 18867 23064
rect 16754 23008 16764 23044
rect 16800 23030 18867 23044
rect 16800 23008 18200 23030
rect 16754 22993 18200 23008
rect 7546 22882 9386 22892
rect 7546 22861 8536 22882
rect 8618 22861 9386 22882
rect 7546 22827 7575 22861
rect 7609 22827 7667 22861
rect 7701 22827 7759 22861
rect 7793 22827 7851 22861
rect 7885 22827 7943 22861
rect 7977 22827 8035 22861
rect 8069 22827 8127 22861
rect 8161 22827 8219 22861
rect 8253 22827 8311 22861
rect 8345 22827 8403 22861
rect 8437 22827 8495 22861
rect 8529 22827 8536 22861
rect 8621 22827 8679 22861
rect 8713 22827 8771 22861
rect 8805 22827 8863 22861
rect 8897 22827 8955 22861
rect 8989 22827 9047 22861
rect 9081 22827 9139 22861
rect 9173 22827 9231 22861
rect 9265 22827 9323 22861
rect 9357 22827 9386 22861
rect 7546 22802 8536 22827
rect 8618 22802 9386 22827
rect 9760 22890 11600 22900
rect 9760 22869 10750 22890
rect 10832 22869 11600 22890
rect 9760 22835 9789 22869
rect 9823 22835 9881 22869
rect 9915 22835 9973 22869
rect 10007 22835 10065 22869
rect 10099 22835 10157 22869
rect 10191 22835 10249 22869
rect 10283 22835 10341 22869
rect 10375 22835 10433 22869
rect 10467 22835 10525 22869
rect 10559 22835 10617 22869
rect 10651 22835 10709 22869
rect 10743 22835 10750 22869
rect 10835 22835 10893 22869
rect 10927 22835 10985 22869
rect 11019 22835 11077 22869
rect 11111 22835 11169 22869
rect 11203 22835 11261 22869
rect 11295 22835 11353 22869
rect 11387 22835 11445 22869
rect 11479 22835 11537 22869
rect 11571 22835 11600 22869
rect 9760 22810 10750 22835
rect 10832 22810 11600 22835
rect 9760 22804 11600 22810
rect 11960 22872 13800 22882
rect 11960 22851 12950 22872
rect 13032 22851 13800 22872
rect 11960 22817 11989 22851
rect 12023 22817 12081 22851
rect 12115 22817 12173 22851
rect 12207 22817 12265 22851
rect 12299 22817 12357 22851
rect 12391 22817 12449 22851
rect 12483 22817 12541 22851
rect 12575 22817 12633 22851
rect 12667 22817 12725 22851
rect 12759 22817 12817 22851
rect 12851 22817 12909 22851
rect 12943 22817 12950 22851
rect 13035 22817 13093 22851
rect 13127 22817 13185 22851
rect 13219 22817 13277 22851
rect 13311 22817 13369 22851
rect 13403 22817 13461 22851
rect 13495 22817 13553 22851
rect 13587 22817 13645 22851
rect 13679 22817 13737 22851
rect 13771 22817 13800 22851
rect 7546 22796 9386 22802
rect 11960 22792 12950 22817
rect 13032 22792 13800 22817
rect 14174 22880 16014 22890
rect 14174 22859 15164 22880
rect 15246 22859 16014 22880
rect 14174 22825 14203 22859
rect 14237 22825 14295 22859
rect 14329 22825 14387 22859
rect 14421 22825 14479 22859
rect 14513 22825 14571 22859
rect 14605 22825 14663 22859
rect 14697 22825 14755 22859
rect 14789 22825 14847 22859
rect 14881 22825 14939 22859
rect 14973 22825 15031 22859
rect 15065 22825 15123 22859
rect 15157 22825 15164 22859
rect 15249 22825 15307 22859
rect 15341 22825 15399 22859
rect 15433 22825 15491 22859
rect 15525 22825 15583 22859
rect 15617 22825 15675 22859
rect 15709 22825 15767 22859
rect 15801 22825 15859 22859
rect 15893 22825 15951 22859
rect 15985 22825 16014 22859
rect 14174 22800 15164 22825
rect 15246 22800 16014 22825
rect 16480 22888 18320 22898
rect 16480 22867 17470 22888
rect 17552 22867 18320 22888
rect 16480 22833 16509 22867
rect 16543 22833 16601 22867
rect 16635 22833 16693 22867
rect 16727 22833 16785 22867
rect 16819 22833 16877 22867
rect 16911 22833 16969 22867
rect 17003 22833 17061 22867
rect 17095 22833 17153 22867
rect 17187 22833 17245 22867
rect 17279 22833 17337 22867
rect 17371 22833 17429 22867
rect 17463 22833 17470 22867
rect 17555 22833 17613 22867
rect 17647 22833 17705 22867
rect 17739 22833 17797 22867
rect 17831 22833 17889 22867
rect 17923 22833 17981 22867
rect 18015 22833 18073 22867
rect 18107 22833 18165 22867
rect 18199 22833 18257 22867
rect 18291 22833 18320 22867
rect 16480 22808 17470 22833
rect 17552 22808 18320 22833
rect 16480 22802 18320 22808
rect 14174 22794 16014 22800
rect 11960 22786 13800 22792
rect 6269 18339 26063 18485
rect 9658 17762 9778 17828
rect 16267 17714 16621 17732
rect 16267 17701 16455 17714
rect 16523 17701 16621 17714
rect 15481 17674 15843 17694
rect 15481 17663 15683 17674
rect 15751 17663 15843 17674
rect 15481 17629 15510 17663
rect 15544 17629 15596 17663
rect 15630 17629 15683 17663
rect 15751 17629 15780 17663
rect 15814 17629 15843 17663
rect 16267 17667 16296 17701
rect 16330 17667 16374 17701
rect 16408 17667 16455 17701
rect 16523 17667 16558 17701
rect 16592 17667 16621 17701
rect 16267 17652 16455 17667
rect 16523 17652 16621 17667
rect 16267 17636 16621 17652
rect 17133 17714 17495 17734
rect 17133 17703 17335 17714
rect 17403 17703 17495 17714
rect 17133 17669 17162 17703
rect 17196 17669 17248 17703
rect 17282 17669 17335 17703
rect 17403 17669 17432 17703
rect 17466 17669 17495 17703
rect 17911 17704 18263 17724
rect 19027 17708 19385 17726
rect 19027 17706 19219 17708
rect 17911 17698 18121 17704
rect 17133 17652 17335 17669
rect 17403 17652 17495 17669
rect 17133 17638 17495 17652
rect 17909 17693 18121 17698
rect 18189 17693 18263 17704
rect 17909 17659 17940 17693
rect 17974 17659 18016 17693
rect 18050 17659 18108 17693
rect 18189 17659 18200 17693
rect 18234 17659 18263 17693
rect 17909 17642 18121 17659
rect 18189 17642 18263 17659
rect 17909 17632 18263 17642
rect 19025 17695 19219 17706
rect 19287 17695 19385 17708
rect 19025 17661 19056 17695
rect 19090 17661 19138 17695
rect 19172 17661 19219 17695
rect 19287 17661 19322 17695
rect 19356 17661 19385 17695
rect 19025 17646 19219 17661
rect 19287 17646 19385 17661
rect 19025 17640 19385 17646
rect 15481 17612 15683 17629
rect 15751 17612 15843 17629
rect 17911 17628 18263 17632
rect 19027 17630 19385 17640
rect 19893 17708 20259 17728
rect 19893 17697 20099 17708
rect 20167 17697 20259 17708
rect 19893 17663 19922 17697
rect 19956 17663 20012 17697
rect 20046 17663 20099 17697
rect 20167 17663 20196 17697
rect 20230 17663 20259 17697
rect 19893 17646 20099 17663
rect 20167 17646 20259 17663
rect 19893 17632 20259 17646
rect 20663 17698 21027 17718
rect 20663 17687 20885 17698
rect 20953 17687 21027 17698
rect 20663 17653 20692 17687
rect 20726 17653 20780 17687
rect 20814 17653 20872 17687
rect 20953 17653 20964 17687
rect 20998 17653 21027 17687
rect 20663 17636 20885 17653
rect 20953 17636 21027 17653
rect 20663 17622 21027 17636
rect 21365 17698 21733 17716
rect 21365 17685 21475 17698
rect 21543 17685 21733 17698
rect 21365 17651 21394 17685
rect 21428 17651 21475 17685
rect 21543 17651 21578 17685
rect 21612 17651 21670 17685
rect 21704 17651 21733 17685
rect 21365 17636 21475 17651
rect 21543 17636 21733 17651
rect 21365 17620 21733 17636
rect 22149 17698 22515 17718
rect 22149 17687 22355 17698
rect 22423 17687 22515 17698
rect 22149 17653 22178 17687
rect 22212 17653 22268 17687
rect 22302 17653 22355 17687
rect 22423 17653 22452 17687
rect 22486 17653 22515 17687
rect 22149 17636 22355 17653
rect 22423 17636 22515 17653
rect 22149 17622 22515 17636
rect 23007 17688 23373 17708
rect 23007 17677 23141 17688
rect 23209 17677 23373 17688
rect 23007 17643 23036 17677
rect 23070 17643 23128 17677
rect 23209 17643 23220 17677
rect 23254 17643 23310 17677
rect 23344 17643 23373 17677
rect 23007 17626 23141 17643
rect 23209 17626 23373 17643
rect 23007 17612 23373 17626
rect 15481 17598 15843 17612
rect 6603 17576 9539 17587
rect 6603 17504 6646 17576
rect 6722 17568 9539 17576
rect 6722 17532 9496 17568
rect 9532 17532 9539 17568
rect 6722 17504 9539 17532
rect 6603 17497 9539 17504
rect 9573 17572 13733 17587
rect 9573 17536 9596 17572
rect 9632 17536 13733 17572
rect 9573 17497 13733 17536
rect 9676 17220 9796 17286
rect 9045 17054 11482 17055
rect 9036 17042 11482 17054
rect 9036 17041 11414 17042
rect 8787 16986 11414 17041
rect 11474 16986 11482 17042
rect 8787 16977 11482 16986
rect 8787 16964 9497 16977
rect 8787 16963 9000 16964
rect 9160 16963 9497 16964
rect 4364 16550 4484 16616
rect 4360 16010 4480 16076
rect 4490 15806 4610 15872
rect 6548 15690 6668 15756
rect 6578 15408 6682 15424
rect 6578 15356 6608 15408
rect 6660 15356 6682 15408
rect 7350 15390 7619 15440
rect 6578 15342 6682 15356
rect 4506 15268 4626 15334
rect 5748 15208 5806 15274
rect 6546 15156 6666 15222
rect 4406 14986 4526 15052
rect 5748 14654 5794 14716
rect 7569 14673 7619 15390
rect 5748 14650 5806 14654
rect 7351 14623 7619 14673
rect 4400 14446 4520 14512
rect 4500 14246 4620 14312
rect 5740 14240 5860 14306
rect 8226 14218 8346 14284
rect 8787 14096 8865 16963
rect 9334 16630 9978 16638
rect 9248 16628 9978 16630
rect 9248 16607 9456 16628
rect 9508 16607 9978 16628
rect 9248 16573 9363 16607
rect 9397 16573 9455 16607
rect 9508 16574 9547 16607
rect 9489 16573 9547 16574
rect 9581 16573 9639 16607
rect 9673 16573 9731 16607
rect 9765 16573 9823 16607
rect 9857 16573 9915 16607
rect 9949 16573 9978 16607
rect 9248 16564 9978 16573
rect 9334 16542 9978 16564
rect 9412 16296 9472 16542
rect 10812 16410 11014 16442
rect 10812 16408 10872 16410
rect 9898 16394 10872 16408
rect 9898 16356 9910 16394
rect 9944 16356 10872 16394
rect 9898 16344 10872 16356
rect 10942 16408 11014 16410
rect 10942 16344 11125 16408
rect 9898 16342 11125 16344
rect 10812 16316 11014 16342
rect 9412 16262 9420 16296
rect 9454 16262 9472 16296
rect 9412 16242 9472 16262
rect 9502 16298 9612 16312
rect 9502 16264 9540 16298
rect 9574 16264 9612 16298
rect 9502 16256 9612 16264
rect 9536 16094 9567 16256
rect 9334 16088 9978 16094
rect 9232 16078 9978 16088
rect 9232 16063 9842 16078
rect 9900 16063 9978 16078
rect 9232 16029 9363 16063
rect 9397 16029 9455 16063
rect 9489 16029 9547 16063
rect 9581 16029 9639 16063
rect 9673 16029 9731 16063
rect 9765 16029 9823 16063
rect 9900 16029 9915 16063
rect 9949 16029 9978 16063
rect 9232 16024 9842 16029
rect 9900 16024 9978 16029
rect 9232 16022 9978 16024
rect 9334 15998 9978 16022
rect 9432 15882 9892 15894
rect 9358 15878 9892 15882
rect 9358 15863 9612 15878
rect 9674 15863 9892 15878
rect 9358 15829 9461 15863
rect 9495 15829 9553 15863
rect 9587 15829 9612 15863
rect 9679 15829 9737 15863
rect 9771 15829 9829 15863
rect 9863 15829 9892 15863
rect 9358 15818 9612 15829
rect 9674 15818 9892 15829
rect 9358 15816 9892 15818
rect 9432 15798 9892 15816
rect 9440 15574 9516 15590
rect 9642 15574 9696 15798
rect 11059 15637 11125 16342
rect 11474 15772 12118 15784
rect 11410 15753 11578 15772
rect 11646 15753 12118 15772
rect 11410 15719 11503 15753
rect 11537 15719 11578 15753
rect 11646 15719 11687 15753
rect 11721 15719 11779 15753
rect 11813 15719 11871 15753
rect 11905 15719 11963 15753
rect 11997 15719 12055 15753
rect 12089 15719 12118 15753
rect 11410 15710 11578 15719
rect 11646 15710 12118 15719
rect 11410 15706 12118 15710
rect 11474 15688 12118 15706
rect 9440 15534 9454 15574
rect 9496 15534 9516 15574
rect 9440 15518 9516 15534
rect 9632 15564 9700 15574
rect 11059 15571 11913 15637
rect 11657 15568 11723 15571
rect 9632 15524 9644 15564
rect 9686 15524 9700 15564
rect 9450 15350 9504 15518
rect 9632 15512 9700 15524
rect 9824 15506 9910 15514
rect 9824 15494 9842 15506
rect 9824 15460 9836 15494
rect 9824 15452 9842 15460
rect 9896 15452 9910 15506
rect 9824 15440 9910 15452
rect 10060 15462 11722 15520
rect 10060 15456 11723 15462
rect 9632 15350 9700 15352
rect 9432 15338 9892 15350
rect 9368 15336 9892 15338
rect 9368 15319 9764 15336
rect 9832 15319 9892 15336
rect 9368 15285 9461 15319
rect 9495 15285 9553 15319
rect 9587 15285 9645 15319
rect 9679 15285 9737 15319
rect 9863 15285 9892 15319
rect 9368 15274 9764 15285
rect 9832 15274 9892 15285
rect 9368 15272 9892 15274
rect 9432 15254 9892 15272
rect 9344 15058 9988 15074
rect 9288 15056 9988 15058
rect 9288 15043 9448 15056
rect 9514 15043 9988 15056
rect 9288 15009 9373 15043
rect 9407 15009 9448 15043
rect 9514 15009 9557 15043
rect 9591 15009 9649 15043
rect 9683 15009 9741 15043
rect 9775 15009 9833 15043
rect 9867 15009 9925 15043
rect 9959 15009 9988 15043
rect 9288 14992 9448 15009
rect 9344 14990 9448 14992
rect 9514 14990 9988 15009
rect 9344 14978 9988 14990
rect 9422 14732 9482 14978
rect 10060 14946 10124 15456
rect 11657 15438 11723 15456
rect 11444 15412 11548 15428
rect 11444 15360 11474 15412
rect 11526 15404 11548 15412
rect 11534 15368 11548 15404
rect 11657 15402 11670 15438
rect 11704 15402 11723 15438
rect 11657 15394 11723 15402
rect 11526 15360 11548 15368
rect 11444 15346 11548 15360
rect 11847 15384 11913 15571
rect 12044 15444 12100 15448
rect 12044 15436 12485 15444
rect 12044 15402 12056 15436
rect 12090 15402 12485 15436
rect 12044 15394 12485 15402
rect 12044 15390 12100 15394
rect 12213 15390 12263 15394
rect 11847 15348 11864 15384
rect 11898 15348 11913 15384
rect 11756 15318 11814 15334
rect 11214 15314 11814 15318
rect 10618 15268 11076 15284
rect 11214 15280 11768 15314
rect 11802 15280 11814 15314
rect 11214 15274 11814 15280
rect 10618 15253 10996 15268
rect 10618 15219 10645 15253
rect 10679 15219 10737 15253
rect 10771 15219 10829 15253
rect 10863 15219 10921 15253
rect 10955 15219 10996 15253
rect 10618 15210 10996 15219
rect 10616 15206 10996 15210
rect 11064 15206 11076 15268
rect 10616 15188 11076 15206
rect 11216 15160 11296 15274
rect 11756 15268 11814 15274
rect 11847 15270 11913 15348
rect 11474 15230 12118 15240
rect 11404 15222 12118 15230
rect 11404 15209 11980 15222
rect 12048 15209 12118 15222
rect 11404 15175 11503 15209
rect 11537 15175 11595 15209
rect 11629 15175 11687 15209
rect 11721 15175 11779 15209
rect 11813 15175 11871 15209
rect 11905 15175 11963 15209
rect 12048 15175 12055 15209
rect 12089 15175 12118 15209
rect 11404 15164 11980 15175
rect 10970 15152 11296 15160
rect 9906 14934 10124 14946
rect 9906 14900 9922 14934
rect 9956 14900 10124 14934
rect 9906 14882 10124 14900
rect 10156 15084 10886 15136
rect 10970 15116 11010 15152
rect 11050 15116 11296 15152
rect 11474 15160 11980 15164
rect 12048 15160 12118 15175
rect 11474 15144 12118 15160
rect 10970 15102 11296 15116
rect 9422 14698 9430 14732
rect 9464 14698 9482 14732
rect 9422 14678 9482 14698
rect 9512 14734 9622 14748
rect 9512 14700 9550 14734
rect 9584 14700 9622 14734
rect 9512 14692 9622 14700
rect 9546 14530 9577 14692
rect 9344 14518 9988 14530
rect 9272 14512 9988 14518
rect 9272 14499 9878 14512
rect 9944 14499 9988 14512
rect 9272 14465 9373 14499
rect 9407 14465 9465 14499
rect 9499 14465 9557 14499
rect 9591 14465 9649 14499
rect 9683 14465 9741 14499
rect 9775 14465 9833 14499
rect 9867 14465 9878 14499
rect 9959 14465 9988 14499
rect 9272 14452 9878 14465
rect 9344 14446 9878 14452
rect 9944 14446 9988 14465
rect 9344 14434 9988 14446
rect 9442 14320 9902 14330
rect 9368 14318 9902 14320
rect 9368 14299 9548 14318
rect 9620 14299 9902 14318
rect 9368 14265 9471 14299
rect 9505 14265 9548 14299
rect 9620 14265 9655 14299
rect 9689 14265 9747 14299
rect 9781 14265 9839 14299
rect 9873 14265 9902 14299
rect 9368 14254 9548 14265
rect 9442 14248 9548 14254
rect 9620 14248 9902 14265
rect 9442 14234 9902 14248
rect 8182 14076 8865 14096
rect 8182 14036 8212 14076
rect 8254 14036 8865 14076
rect 8182 14018 8865 14036
rect 8602 13990 8638 14018
rect 9450 14010 9526 14028
rect 9654 14010 9700 14234
rect 7636 13974 7742 13976
rect 7636 13938 7806 13974
rect 9450 13970 9464 14010
rect 9506 13970 9526 14010
rect 9450 13954 9526 13970
rect 9642 14000 9710 14010
rect 9642 13960 9654 14000
rect 9696 13960 9710 14000
rect 7636 13936 7752 13938
rect 7208 13854 7328 13920
rect 7636 13882 7652 13936
rect 7704 13904 7752 13936
rect 7792 13904 7806 13938
rect 7704 13882 7806 13904
rect 7636 13856 7806 13882
rect 9458 13786 9512 13954
rect 9642 13948 9710 13960
rect 9832 13904 10004 13918
rect 9832 13888 9896 13904
rect 9832 13854 9844 13888
rect 9880 13854 9896 13888
rect 9832 13842 9896 13854
rect 9956 13842 10004 13904
rect 9832 13824 10004 13842
rect 9442 13774 9902 13786
rect 4490 13702 4610 13768
rect 9442 13768 9750 13774
rect 5734 13690 5854 13756
rect 9368 13755 9750 13768
rect 9822 13755 9902 13774
rect 7640 13738 7734 13754
rect 7640 13676 7656 13738
rect 7724 13676 7734 13738
rect 8244 13676 8364 13742
rect 9368 13721 9471 13755
rect 9505 13721 9563 13755
rect 9597 13721 9655 13755
rect 9689 13721 9747 13755
rect 9822 13721 9839 13755
rect 9873 13721 9902 13755
rect 9368 13704 9750 13721
rect 9822 13704 9902 13721
rect 9368 13702 9902 13704
rect 9442 13690 9902 13702
rect 7640 13656 7734 13676
rect 5874 13450 5994 13454
rect 5874 13390 5984 13450
rect 5874 13388 5994 13390
rect 9336 13388 9980 13406
rect 4394 13316 4514 13382
rect 7188 13378 7308 13388
rect 9336 13380 9442 13388
rect 7204 13322 7308 13378
rect 9264 13375 9442 13380
rect 9514 13375 9980 13388
rect 9264 13341 9365 13375
rect 9399 13341 9442 13375
rect 9514 13341 9549 13375
rect 9583 13341 9641 13375
rect 9675 13341 9733 13375
rect 9767 13341 9825 13375
rect 9859 13341 9917 13375
rect 9951 13341 9980 13375
rect 9264 13322 9442 13341
rect 9514 13322 9980 13341
rect 9264 13314 9980 13322
rect 9336 13310 9980 13314
rect 10156 13370 10208 15084
rect 10834 14960 10886 15084
rect 10636 14955 10772 14956
rect 10428 14942 10772 14955
rect 10428 14908 10690 14942
rect 10724 14908 10772 14942
rect 10428 14882 10772 14908
rect 10806 14942 10886 14960
rect 10806 14908 10830 14942
rect 10866 14908 10886 14942
rect 10806 14894 10886 14908
rect 10428 14877 10711 14882
rect 10428 13975 10506 14877
rect 12435 14741 12485 15394
rect 12341 14740 12485 14741
rect 10618 14720 11076 14740
rect 10618 14709 10660 14720
rect 10728 14709 11076 14720
rect 10618 14675 10645 14709
rect 10728 14675 10737 14709
rect 10771 14675 10829 14709
rect 10863 14675 10921 14709
rect 10955 14675 11013 14709
rect 11047 14675 11076 14709
rect 12209 14691 12485 14740
rect 13643 14697 13733 17497
rect 16399 17468 16461 17478
rect 16399 17466 16413 17468
rect 15360 17436 15683 17458
rect 14960 17407 15026 17436
rect 15122 17407 15635 17436
rect 14960 16366 14989 17407
rect 15360 17402 15635 17407
rect 15669 17402 15683 17436
rect 15360 17368 15683 17402
rect 15713 17428 15902 17448
rect 15713 17394 15725 17428
rect 15763 17411 15902 17428
rect 15943 17436 16413 17466
rect 15943 17411 15973 17436
rect 16187 17434 16217 17436
rect 16399 17434 16413 17436
rect 16449 17434 16461 17468
rect 15763 17394 15973 17411
rect 16399 17410 16461 17434
rect 16493 17476 17335 17498
rect 16493 17464 17287 17476
rect 16493 17430 16517 17464
rect 16551 17442 17287 17464
rect 17321 17442 17335 17476
rect 16551 17430 17335 17442
rect 16493 17408 17335 17430
rect 17365 17472 18103 17488
rect 17365 17468 18059 17472
rect 17365 17434 17377 17468
rect 17415 17438 18059 17468
rect 18097 17438 18103 17472
rect 17415 17434 18103 17438
rect 17365 17414 18103 17434
rect 18133 17474 18201 17490
rect 18133 17472 19179 17474
rect 18133 17462 19225 17472
rect 18133 17460 19177 17462
rect 18133 17426 18147 17460
rect 18183 17428 19177 17460
rect 19213 17428 19225 17462
rect 18183 17426 19225 17428
rect 18133 17418 19225 17426
rect 18133 17406 18201 17418
rect 19163 17404 19225 17418
rect 19257 17470 20099 17492
rect 20897 17483 20963 17484
rect 19257 17458 20051 17470
rect 19257 17424 19281 17458
rect 19315 17436 20051 17458
rect 20085 17436 20099 17470
rect 19315 17424 20099 17436
rect 19257 17402 20099 17424
rect 20129 17466 20867 17482
rect 20129 17462 20823 17466
rect 20129 17428 20141 17462
rect 20179 17432 20823 17462
rect 20861 17432 20867 17466
rect 20179 17428 20867 17432
rect 20129 17408 20867 17428
rect 20897 17468 21107 17483
rect 20897 17462 21425 17468
rect 20897 17454 21481 17462
rect 20897 17420 20911 17454
rect 20947 17452 21481 17454
rect 20947 17422 21433 17452
rect 20947 17420 20963 17422
rect 21305 17420 21433 17422
rect 20897 17400 20963 17420
rect 21419 17418 21433 17420
rect 21469 17418 21481 17452
rect 21419 17394 21481 17418
rect 21513 17460 22355 17482
rect 23153 17473 23219 17474
rect 21513 17448 22307 17460
rect 21513 17414 21537 17448
rect 21571 17426 22307 17448
rect 22341 17426 22355 17460
rect 21571 17414 22355 17426
rect 15713 17381 15973 17394
rect 21513 17392 22355 17414
rect 22385 17456 23123 17472
rect 22385 17452 23079 17456
rect 22385 17418 22397 17452
rect 22435 17422 23079 17452
rect 23117 17422 23123 17456
rect 22435 17418 23123 17422
rect 22385 17398 23123 17418
rect 23153 17444 23432 17473
rect 23153 17410 23167 17444
rect 23203 17443 23432 17444
rect 23203 17410 23219 17443
rect 23153 17390 23219 17410
rect 15713 17374 15902 17381
rect 16267 17172 16621 17188
rect 16267 17157 16453 17172
rect 16521 17157 16621 17172
rect 15481 17134 15843 17150
rect 15481 17119 15691 17134
rect 15759 17119 15843 17134
rect 15481 17085 15510 17119
rect 15544 17085 15596 17119
rect 15630 17085 15688 17119
rect 15759 17085 15780 17119
rect 15814 17085 15843 17119
rect 16267 17123 16296 17157
rect 16330 17123 16374 17157
rect 16408 17123 16453 17157
rect 16521 17123 16558 17157
rect 16592 17123 16621 17157
rect 16267 17110 16453 17123
rect 16521 17110 16621 17123
rect 16267 17092 16621 17110
rect 17133 17174 17495 17190
rect 17133 17159 17343 17174
rect 17411 17159 17495 17174
rect 17911 17166 18263 17180
rect 17911 17160 18101 17166
rect 17133 17125 17162 17159
rect 17196 17125 17248 17159
rect 17282 17125 17340 17159
rect 17411 17125 17432 17159
rect 17466 17125 17495 17159
rect 17133 17112 17343 17125
rect 17411 17112 17495 17125
rect 17133 17094 17495 17112
rect 17905 17149 18101 17160
rect 18169 17149 18263 17166
rect 17905 17115 17940 17149
rect 17974 17115 18016 17149
rect 18050 17115 18101 17149
rect 18169 17115 18200 17149
rect 18234 17115 18263 17149
rect 17905 17104 18101 17115
rect 18169 17104 18263 17115
rect 17905 17094 18263 17104
rect 15481 17072 15691 17085
rect 15759 17072 15843 17085
rect 17911 17084 18263 17094
rect 19027 17166 19385 17182
rect 19027 17151 19217 17166
rect 19285 17151 19385 17166
rect 19027 17117 19056 17151
rect 19090 17117 19138 17151
rect 19172 17117 19217 17151
rect 19285 17117 19322 17151
rect 19356 17117 19385 17151
rect 19027 17104 19217 17117
rect 19285 17104 19385 17117
rect 19027 17086 19385 17104
rect 19893 17168 20259 17184
rect 19893 17153 20107 17168
rect 20175 17153 20259 17168
rect 19893 17119 19922 17153
rect 19956 17119 20012 17153
rect 20046 17119 20104 17153
rect 20175 17119 20196 17153
rect 20230 17119 20259 17153
rect 19893 17106 20107 17119
rect 20175 17106 20259 17119
rect 19893 17088 20259 17106
rect 20663 17160 21027 17174
rect 20663 17143 20865 17160
rect 20933 17143 21027 17160
rect 20663 17109 20692 17143
rect 20726 17109 20780 17143
rect 20814 17109 20865 17143
rect 20933 17109 20964 17143
rect 20998 17109 21027 17143
rect 20663 17098 20865 17109
rect 20933 17098 21027 17109
rect 20663 17078 21027 17098
rect 21365 17156 21733 17172
rect 21365 17141 21473 17156
rect 21541 17141 21733 17156
rect 21365 17107 21394 17141
rect 21428 17107 21473 17141
rect 21541 17107 21578 17141
rect 21612 17107 21670 17141
rect 21704 17107 21733 17141
rect 21365 17094 21473 17107
rect 21541 17094 21733 17107
rect 21365 17076 21733 17094
rect 22149 17158 22515 17174
rect 22149 17143 22363 17158
rect 22431 17143 22515 17158
rect 22149 17109 22178 17143
rect 22212 17109 22268 17143
rect 22302 17109 22360 17143
rect 22431 17109 22452 17143
rect 22486 17109 22515 17143
rect 22149 17096 22363 17109
rect 22431 17096 22515 17109
rect 22149 17078 22515 17096
rect 23007 17150 23373 17164
rect 23007 17133 23121 17150
rect 23189 17133 23373 17150
rect 23007 17099 23036 17133
rect 23070 17099 23121 17133
rect 23189 17099 23220 17133
rect 23254 17099 23310 17133
rect 23344 17099 23373 17133
rect 23007 17088 23121 17099
rect 23189 17088 23373 17099
rect 15481 17054 15843 17072
rect 23007 17068 23373 17088
rect 23402 16937 23432 17443
rect 23402 16906 23479 16937
rect 23403 16877 23479 16906
rect 16260 16658 16380 16724
rect 17346 16652 17466 16718
rect 17902 16662 18022 16728
rect 18828 16652 18948 16718
rect 19596 16644 19716 16710
rect 20468 16644 20588 16710
rect 21594 16650 21714 16716
rect 22346 16640 22466 16706
rect 23224 16644 23344 16710
rect 16400 16400 16466 16420
rect 16400 16367 16416 16400
rect 16224 16366 16416 16367
rect 16452 16366 16466 16400
rect 14960 16337 15026 16366
rect 15122 16337 16466 16366
rect 16496 16392 17234 16412
rect 16496 16388 17184 16392
rect 16496 16354 16502 16388
rect 16540 16358 17184 16388
rect 17222 16358 17234 16392
rect 16540 16354 17234 16358
rect 16496 16338 17234 16354
rect 17264 16396 18106 16418
rect 17264 16384 18048 16396
rect 17264 16350 17278 16384
rect 17312 16362 18048 16384
rect 18082 16362 18106 16396
rect 17312 16350 18106 16362
rect 16400 16336 16466 16337
rect 17264 16328 18106 16350
rect 18138 16392 18200 16416
rect 18138 16358 18150 16392
rect 18186 16390 18200 16392
rect 18656 16390 18722 16410
rect 18186 16388 18314 16390
rect 18656 16388 18672 16390
rect 18186 16358 18672 16388
rect 18138 16356 18672 16358
rect 18708 16356 18722 16390
rect 18138 16348 18722 16356
rect 18194 16342 18722 16348
rect 18512 16327 18722 16342
rect 18752 16382 19490 16402
rect 18752 16378 19440 16382
rect 18752 16344 18758 16378
rect 18796 16348 19440 16378
rect 19478 16348 19490 16382
rect 18796 16344 19490 16348
rect 18752 16328 19490 16344
rect 19520 16386 20362 16408
rect 19520 16374 20304 16386
rect 19520 16340 19534 16374
rect 19568 16352 20304 16374
rect 20338 16352 20362 16386
rect 19568 16340 20362 16352
rect 18656 16326 18722 16327
rect 19520 16318 20362 16340
rect 20394 16392 20456 16406
rect 21418 16392 21486 16404
rect 20394 16384 21486 16392
rect 20394 16382 21436 16384
rect 20394 16348 20406 16382
rect 20442 16350 21436 16382
rect 21472 16350 21486 16384
rect 20442 16348 21486 16350
rect 20394 16338 21486 16348
rect 20440 16336 21486 16338
rect 21418 16320 21486 16336
rect 21516 16376 22254 16396
rect 21516 16372 22204 16376
rect 21516 16338 21522 16372
rect 21560 16342 22204 16372
rect 22242 16342 22254 16376
rect 21560 16338 22254 16342
rect 21516 16322 22254 16338
rect 22284 16380 23126 16402
rect 22284 16368 23068 16380
rect 22284 16334 22298 16368
rect 22332 16346 23068 16368
rect 23102 16346 23126 16380
rect 22332 16334 23126 16346
rect 22284 16312 23126 16334
rect 23158 16376 23220 16400
rect 23158 16342 23170 16376
rect 23206 16374 23220 16376
rect 23449 16374 23479 16877
rect 23206 16344 23479 16374
rect 23206 16342 23220 16344
rect 23158 16332 23220 16342
rect 16252 16118 16372 16184
rect 21575 16178 21605 16182
rect 17334 16108 17454 16174
rect 17898 16104 18018 16170
rect 18820 16104 18940 16170
rect 19584 16104 19704 16170
rect 20474 16104 20594 16170
rect 21575 16112 21710 16178
rect 21575 16086 21605 16112
rect 22364 16090 22484 16156
rect 23218 16100 23338 16166
rect 23373 15915 23403 15918
rect 23449 15915 23479 16344
rect 23373 15885 23479 15915
rect 23373 15607 23403 15885
rect 23372 15606 23403 15607
rect 22975 15577 23403 15606
rect 22975 14749 23005 15577
rect 25382 14808 25502 14874
rect 22975 14719 23418 14749
rect 10618 14658 10660 14675
rect 10728 14658 11076 14675
rect 10618 14656 11076 14658
rect 10616 14644 11076 14656
rect 10690 14312 11334 14318
rect 10606 14298 11334 14312
rect 10606 14287 11216 14298
rect 11284 14287 11334 14298
rect 10606 14253 10719 14287
rect 10753 14253 10811 14287
rect 10845 14253 10903 14287
rect 10937 14253 10995 14287
rect 11029 14253 11087 14287
rect 11121 14253 11179 14287
rect 11213 14253 11216 14287
rect 11305 14253 11334 14287
rect 10606 14246 11216 14253
rect 10690 14236 11216 14246
rect 11284 14236 11334 14253
rect 10690 14222 11334 14236
rect 12213 14181 12263 14691
rect 13643 14607 22797 14697
rect 23388 14675 23418 14719
rect 24138 14714 24198 14726
rect 23388 14674 23700 14675
rect 23388 14645 23731 14674
rect 23701 14614 23731 14645
rect 24138 14662 24144 14714
rect 24196 14662 24198 14714
rect 24138 14650 24198 14662
rect 25917 14658 26063 18339
rect 24138 14616 24150 14650
rect 24186 14616 24198 14650
rect 12588 14288 13140 14302
rect 12588 14271 12782 14288
rect 12850 14280 13140 14288
rect 12850 14271 13220 14280
rect 12588 14237 12617 14271
rect 12651 14237 12709 14271
rect 12743 14237 12782 14271
rect 12850 14237 12893 14271
rect 12927 14237 12985 14271
rect 13019 14237 13077 14271
rect 13111 14237 13220 14271
rect 12588 14226 12782 14237
rect 12850 14226 13220 14237
rect 12588 14214 13220 14226
rect 12588 14206 13140 14214
rect 13643 14182 13733 14607
rect 22618 14599 22797 14607
rect 22618 14580 23581 14599
rect 22618 14546 23530 14580
rect 23568 14546 23581 14580
rect 22618 14509 23581 14546
rect 23644 14562 23732 14614
rect 24138 14578 24198 14616
rect 23644 14528 23672 14562
rect 23708 14528 23732 14562
rect 22618 14508 22736 14509
rect 23644 14490 23732 14528
rect 24444 14564 24510 14620
rect 24444 14512 24452 14564
rect 24504 14512 24510 14564
rect 24444 14502 24510 14512
rect 24550 14588 24604 14620
rect 24550 14578 24556 14588
rect 24592 14578 24604 14588
rect 24550 14526 24552 14578
rect 24550 14502 24604 14526
rect 24684 14602 24770 14618
rect 24684 14550 24698 14602
rect 24750 14550 24770 14602
rect 24684 14528 24712 14550
rect 24746 14528 24770 14550
rect 24684 14518 24770 14528
rect 25348 14594 26063 14658
rect 25348 14560 25356 14594
rect 25390 14560 26063 14594
rect 25348 14516 26063 14560
rect 25917 14514 26063 14516
rect 24684 14444 24770 14472
rect 23850 14318 24212 14334
rect 23850 14258 23992 14318
rect 24054 14258 24212 14318
rect 25370 14258 25490 14324
rect 23850 14240 24212 14258
rect 12213 14176 12264 14181
rect 12213 14170 12940 14176
rect 12213 14136 12762 14170
rect 12798 14136 12940 14170
rect 12213 14129 12940 14136
rect 12256 14128 12940 14129
rect 13470 14132 13733 14182
rect 13470 14100 13732 14132
rect 12312 14034 12980 14094
rect 10689 13980 10767 14033
rect 12312 14022 12386 14034
rect 10689 13975 10716 13980
rect 10428 13946 10716 13975
rect 10750 13946 10767 13980
rect 10428 13897 10767 13946
rect 10156 13360 10242 13370
rect 9414 13064 9474 13310
rect 10156 13308 10164 13360
rect 10226 13308 10242 13360
rect 10156 13300 10242 13308
rect 10156 13232 10208 13300
rect 9902 13224 10208 13232
rect 9902 13190 9914 13224
rect 9948 13190 10208 13224
rect 9902 13180 10208 13190
rect 10428 13089 10506 13897
rect 10868 13894 10938 13940
rect 10868 13842 10878 13894
rect 10930 13842 10938 13894
rect 10868 13802 10938 13842
rect 10966 13934 11034 13990
rect 10966 13882 10976 13934
rect 11028 13882 11034 13934
rect 10966 13804 11034 13882
rect 11068 13974 11140 13992
rect 11068 13936 11078 13974
rect 11114 13936 11140 13974
rect 11068 13890 11140 13936
rect 11068 13834 11074 13890
rect 11126 13834 11140 13890
rect 11660 13932 12120 13944
rect 12312 13934 12384 14022
rect 12702 13984 12842 13996
rect 12502 13978 12608 13980
rect 12502 13942 12672 13978
rect 12502 13940 12618 13942
rect 11660 13922 12188 13932
rect 11660 13913 11694 13922
rect 11762 13913 12188 13922
rect 11660 13879 11689 13913
rect 11762 13879 11781 13913
rect 11815 13879 11873 13913
rect 11907 13879 11965 13913
rect 11999 13879 12057 13913
rect 12091 13879 12188 13913
rect 11068 13808 11140 13834
rect 11246 13856 11532 13876
rect 11246 13818 11260 13856
rect 11298 13818 11532 13856
rect 11660 13860 11694 13879
rect 11762 13866 12188 13879
rect 11762 13860 12120 13866
rect 11660 13848 12120 13860
rect 11246 13802 11532 13818
rect 11451 13789 11532 13802
rect 12312 13790 12382 13934
rect 12502 13886 12518 13940
rect 12570 13908 12618 13940
rect 12658 13908 12672 13942
rect 12570 13886 12672 13908
rect 12702 13908 12732 13984
rect 12812 13962 12842 13984
rect 12908 13976 12980 14034
rect 13048 14080 13732 14100
rect 13048 14040 13078 14080
rect 13120 14040 13732 14080
rect 13048 14022 13732 14040
rect 13468 13996 13732 14022
rect 13468 13994 13504 13996
rect 12812 13908 12840 13962
rect 12886 13960 12980 13976
rect 12886 13924 12918 13960
rect 12956 13924 12980 13960
rect 12886 13908 12980 13924
rect 12702 13894 12840 13908
rect 12502 13860 12672 13886
rect 10690 13762 11334 13774
rect 10608 13758 11334 13762
rect 10608 13743 10728 13758
rect 10796 13743 11334 13758
rect 10608 13709 10719 13743
rect 10796 13709 10811 13743
rect 10845 13709 10903 13743
rect 10937 13709 10995 13743
rect 11029 13709 11087 13743
rect 11121 13709 11179 13743
rect 11213 13709 11271 13743
rect 11305 13709 11334 13743
rect 11451 13715 11929 13789
rect 11986 13768 12382 13790
rect 11986 13734 12028 13768
rect 12062 13734 12382 13768
rect 11986 13718 12382 13734
rect 12506 13748 13140 13758
rect 12506 13742 13204 13748
rect 10608 13696 10728 13709
rect 10796 13696 11334 13709
rect 10690 13678 11334 13696
rect 11855 13608 11929 13715
rect 12506 13680 12522 13742
rect 12590 13727 13204 13742
rect 12590 13693 12617 13727
rect 12651 13693 12709 13727
rect 12743 13693 12801 13727
rect 12835 13693 12893 13727
rect 12927 13693 12985 13727
rect 13019 13693 13077 13727
rect 13111 13693 13204 13727
rect 12590 13682 13204 13693
rect 12590 13680 13140 13682
rect 12506 13662 13140 13680
rect 12506 13660 12600 13662
rect 11410 13558 11759 13581
rect 11410 13524 11700 13558
rect 11734 13524 11759 13558
rect 11410 13507 11759 13524
rect 11855 13574 11878 13608
rect 11912 13574 11929 13608
rect 10814 13462 11274 13476
rect 10728 13454 11274 13462
rect 10728 13445 10850 13454
rect 10918 13445 11274 13454
rect 10728 13411 10843 13445
rect 10918 13411 10935 13445
rect 10969 13411 11027 13445
rect 11061 13411 11119 13445
rect 11153 13411 11211 13445
rect 11245 13411 11274 13445
rect 10728 13396 10850 13411
rect 10814 13394 10850 13396
rect 10918 13394 11274 13411
rect 10814 13380 11274 13394
rect 10986 13342 11084 13348
rect 10986 13290 11006 13342
rect 11060 13290 11084 13342
rect 11410 13302 11484 13507
rect 11855 13493 11929 13574
rect 11660 13394 12120 13400
rect 11660 13382 12220 13394
rect 11660 13369 12002 13382
rect 12070 13369 12220 13382
rect 11660 13335 11689 13369
rect 11723 13335 11781 13369
rect 11815 13335 11873 13369
rect 11907 13335 11965 13369
rect 11999 13335 12002 13369
rect 12091 13335 12220 13369
rect 11660 13320 12002 13335
rect 12070 13328 12220 13335
rect 12070 13320 12120 13328
rect 11660 13304 12120 13320
rect 10986 13272 11084 13290
rect 11198 13282 11484 13302
rect 11198 13244 11208 13282
rect 11246 13244 11484 13282
rect 11198 13228 11484 13244
rect 9414 13030 9422 13064
rect 9456 13030 9474 13064
rect 9414 13010 9474 13030
rect 9504 13066 9614 13080
rect 9504 13032 9542 13066
rect 9576 13032 9614 13066
rect 9504 13024 9614 13032
rect 10428 13064 10947 13089
rect 10428 13030 10860 13064
rect 10894 13030 10947 13064
rect 5862 12848 5982 12914
rect 9538 12862 9569 13024
rect 10428 13011 10947 13030
rect 11042 13086 11124 13158
rect 11042 13032 11062 13086
rect 11114 13032 11124 13086
rect 9336 12852 9980 12862
rect 9266 12848 9980 12852
rect 4400 12772 4520 12838
rect 9266 12831 9856 12848
rect 9928 12831 9980 12848
rect 9266 12797 9365 12831
rect 9399 12797 9457 12831
rect 9491 12797 9549 12831
rect 9583 12797 9641 12831
rect 9675 12797 9733 12831
rect 9767 12797 9825 12831
rect 9951 12797 9980 12831
rect 9266 12786 9856 12797
rect 9336 12782 9856 12786
rect 9928 12782 9980 12797
rect 9336 12766 9980 12782
rect 9434 12646 9894 12662
rect 9434 12642 9500 12646
rect 4480 12570 4600 12636
rect 9358 12631 9500 12642
rect 9574 12631 9894 12646
rect 9358 12597 9463 12631
rect 9497 12597 9500 12631
rect 9589 12597 9647 12631
rect 9681 12597 9739 12631
rect 9773 12597 9831 12631
rect 9865 12597 9894 12631
rect 9358 12580 9500 12597
rect 9574 12580 9894 12597
rect 9358 12576 9894 12580
rect 9434 12566 9894 12576
rect 5856 12364 5976 12430
rect 9442 12342 9518 12368
rect 9642 12342 9692 12566
rect 9826 12394 9976 12408
rect 9826 12374 9872 12394
rect 9442 12302 9456 12342
rect 9498 12302 9518 12342
rect 9442 12286 9518 12302
rect 9634 12332 9702 12342
rect 9634 12292 9646 12332
rect 9688 12292 9702 12332
rect 9826 12340 9836 12374
rect 9826 12326 9872 12340
rect 9934 12326 9976 12394
rect 9826 12310 9976 12326
rect 9456 12118 9508 12286
rect 9634 12280 9702 12292
rect 10428 12125 10506 13011
rect 11042 12974 11124 13032
rect 10814 12920 11274 12932
rect 10728 12901 10862 12920
rect 10930 12901 11274 12920
rect 10728 12867 10843 12901
rect 10930 12867 10935 12901
rect 10969 12867 11027 12901
rect 11061 12867 11119 12901
rect 11153 12867 11211 12901
rect 11245 12867 11274 12901
rect 10728 12860 10862 12867
rect 10930 12860 11274 12867
rect 10728 12854 11274 12860
rect 10814 12836 11274 12854
rect 10810 12436 11270 12456
rect 10810 12432 11146 12436
rect 10706 12425 11146 12432
rect 11214 12425 11270 12436
rect 10706 12391 10839 12425
rect 10873 12391 10931 12425
rect 10965 12391 11023 12425
rect 11057 12391 11115 12425
rect 11241 12391 11270 12425
rect 10706 12374 11146 12391
rect 11214 12374 11270 12391
rect 10706 12366 11270 12374
rect 10810 12360 11270 12366
rect 11200 12212 11268 12222
rect 11200 12160 11206 12212
rect 11258 12160 11268 12212
rect 11200 12154 11268 12160
rect 9434 12108 9894 12118
rect 9358 12104 9894 12108
rect 4484 12036 4604 12102
rect 9358 12087 9772 12104
rect 9846 12087 9894 12104
rect 9358 12053 9463 12087
rect 9497 12053 9555 12087
rect 9589 12053 9647 12087
rect 9681 12053 9739 12087
rect 9865 12053 9894 12087
rect 9358 12042 9772 12053
rect 9434 12038 9772 12042
rect 9846 12038 9894 12053
rect 9434 12022 9894 12038
rect 10428 12116 10961 12125
rect 10428 12082 10884 12116
rect 10920 12082 10961 12116
rect 10428 12047 10961 12082
rect 11008 12122 11078 12130
rect 11008 12070 11016 12122
rect 11068 12070 11078 12122
rect 11008 12064 11078 12070
rect 5844 11822 5964 11888
rect 9346 11826 9990 11842
rect 9278 11824 9990 11826
rect 4402 11748 4522 11814
rect 9278 11811 9426 11824
rect 9506 11811 9990 11824
rect 9278 11777 9375 11811
rect 9409 11777 9426 11811
rect 9506 11777 9559 11811
rect 9593 11777 9651 11811
rect 9685 11777 9743 11811
rect 9777 11777 9835 11811
rect 9869 11777 9927 11811
rect 9961 11777 9990 11811
rect 9278 11760 9426 11777
rect 9506 11760 9990 11777
rect 9346 11746 9990 11760
rect 9424 11500 9484 11746
rect 10428 11674 10506 12047
rect 10810 11898 11270 11912
rect 10714 11896 11270 11898
rect 10714 11881 10868 11896
rect 10936 11881 11270 11896
rect 10714 11847 10839 11881
rect 10965 11847 11023 11881
rect 11057 11847 11115 11881
rect 11149 11847 11207 11881
rect 11241 11847 11270 11881
rect 10714 11834 10868 11847
rect 10936 11834 11270 11847
rect 10714 11832 11270 11834
rect 10810 11816 11270 11832
rect 9908 11660 10506 11674
rect 9908 11626 9914 11660
rect 9950 11626 10506 11660
rect 9908 11596 10506 11626
rect 9424 11466 9432 11500
rect 9466 11466 9484 11500
rect 9424 11446 9484 11466
rect 9514 11502 9624 11516
rect 9514 11468 9552 11502
rect 9586 11468 9624 11502
rect 9514 11460 9624 11468
rect 9548 11298 9579 11460
rect 4392 11222 4512 11288
rect 9346 11286 9990 11298
rect 9270 11282 9990 11286
rect 9270 11267 9860 11282
rect 9940 11267 9990 11282
rect 9270 11233 9375 11267
rect 9409 11233 9467 11267
rect 9501 11233 9559 11267
rect 9593 11233 9651 11267
rect 9685 11233 9743 11267
rect 9777 11233 9835 11267
rect 9961 11233 9990 11267
rect 9270 11220 9860 11233
rect 9346 11218 9860 11220
rect 9940 11218 9990 11233
rect 9346 11202 9990 11218
rect 9444 11086 9904 11098
rect 4494 11014 4614 11080
rect 9372 11078 9904 11086
rect 9372 11067 9492 11078
rect 9572 11067 9904 11078
rect 9372 11033 9473 11067
rect 9599 11033 9657 11067
rect 9691 11033 9749 11067
rect 9783 11033 9841 11067
rect 9875 11033 9904 11067
rect 9372 11020 9492 11033
rect 9444 11014 9492 11020
rect 9572 11014 9904 11033
rect 9444 11002 9904 11014
rect 9452 10778 9528 10790
rect 4970 10732 5202 10762
rect 4970 10730 5054 10732
rect 4970 10694 4982 10730
rect 5016 10694 5054 10730
rect 4970 10676 5054 10694
rect 5108 10676 5202 10732
rect 9452 10738 9466 10778
rect 9508 10738 9528 10778
rect 9452 10722 9528 10738
rect 9642 10768 9714 11002
rect 9642 10734 9656 10768
rect 9644 10728 9656 10734
rect 9698 10734 9714 10768
rect 9836 10736 10068 10766
rect 9836 10734 9920 10736
rect 9698 10728 9712 10734
rect 4970 10652 5202 10676
rect 9472 10554 9522 10722
rect 9644 10712 9712 10728
rect 9836 10698 9848 10734
rect 9882 10698 9920 10734
rect 9836 10680 9920 10698
rect 9974 10680 10068 10736
rect 9836 10656 10068 10680
rect 9644 10554 9712 10558
rect 9444 10544 9904 10554
rect 4496 10476 4616 10542
rect 9444 10540 9770 10544
rect 9370 10523 9770 10540
rect 9850 10523 9904 10544
rect 9370 10489 9473 10523
rect 9507 10489 9565 10523
rect 9599 10489 9657 10523
rect 9691 10489 9749 10523
rect 9875 10489 9904 10523
rect 9370 10480 9770 10489
rect 9850 10480 9904 10489
rect 9370 10474 9904 10480
rect 9444 10458 9904 10474
rect 6112 6638 6388 6648
rect 6112 6617 6226 6638
rect 6282 6628 6388 6638
rect 6282 6617 6484 6628
rect 6112 6583 6141 6617
rect 6175 6583 6226 6617
rect 6282 6583 6325 6617
rect 6359 6583 6484 6617
rect 6112 6580 6226 6583
rect 6282 6580 6484 6583
rect 6112 6562 6484 6580
rect 6112 6552 6388 6562
rect 6134 6390 6228 6398
rect 6134 6338 6168 6390
rect 6220 6338 6228 6390
rect 6262 6396 6328 6398
rect 6262 6344 6268 6396
rect 6320 6344 6328 6396
rect 6262 6338 6328 6344
rect 6134 6332 6228 6338
rect 6112 6090 6388 6104
rect 6112 6088 6468 6090
rect 6112 6073 6170 6088
rect 6226 6073 6468 6088
rect 6112 6039 6141 6073
rect 6226 6039 6233 6073
rect 6267 6039 6325 6073
rect 6359 6039 6468 6073
rect 6112 6030 6170 6039
rect 6226 6030 6468 6039
rect 6112 6024 6468 6030
rect 6112 6008 6388 6024
rect 10018 6006 11490 6016
rect 9932 6002 11490 6006
rect 9932 5985 10406 6002
rect 10464 6000 11490 6002
rect 10464 5985 10774 6000
rect 10832 5985 11490 6000
rect 12080 5994 13552 6004
rect 14038 5996 15510 6012
rect 16032 6008 17504 6018
rect 9932 5951 10047 5985
rect 10081 5951 10139 5985
rect 10173 5951 10231 5985
rect 10265 5951 10323 5985
rect 10357 5951 10406 5985
rect 10464 5951 10507 5985
rect 10541 5951 10599 5985
rect 10633 5951 10691 5985
rect 10725 5951 10774 5985
rect 10832 5951 10875 5985
rect 10909 5951 10967 5985
rect 11001 5951 11059 5985
rect 11093 5951 11151 5985
rect 11185 5951 11243 5985
rect 11277 5951 11335 5985
rect 11369 5951 11427 5985
rect 11461 5951 11490 5985
rect 9932 5940 10406 5951
rect 10464 5940 10774 5951
rect 10018 5936 10774 5940
rect 10832 5936 11490 5951
rect 10018 5920 11490 5936
rect 12010 5986 13552 5994
rect 12010 5973 12796 5986
rect 12852 5973 13552 5986
rect 12010 5939 12109 5973
rect 12143 5939 12201 5973
rect 12235 5939 12293 5973
rect 12327 5939 12385 5973
rect 12419 5939 12477 5973
rect 12511 5939 12569 5973
rect 12603 5939 12661 5973
rect 12695 5939 12753 5973
rect 12787 5939 12796 5973
rect 12879 5939 12937 5973
rect 12971 5939 13029 5973
rect 13063 5939 13121 5973
rect 13155 5939 13213 5973
rect 13247 5939 13305 5973
rect 13339 5939 13397 5973
rect 13431 5939 13489 5973
rect 13523 5939 13552 5973
rect 12010 5928 12796 5939
rect 12852 5928 13552 5939
rect 13944 5994 15510 5996
rect 13944 5981 14754 5994
rect 14810 5981 15510 5994
rect 13944 5947 14067 5981
rect 14101 5947 14159 5981
rect 14193 5947 14251 5981
rect 14285 5947 14343 5981
rect 14377 5947 14435 5981
rect 14469 5947 14527 5981
rect 14561 5947 14619 5981
rect 14653 5947 14711 5981
rect 14745 5947 14754 5981
rect 14837 5947 14895 5981
rect 14929 5947 14987 5981
rect 15021 5947 15079 5981
rect 15113 5947 15171 5981
rect 15205 5947 15263 5981
rect 15297 5947 15355 5981
rect 15389 5947 15447 5981
rect 15481 5947 15510 5981
rect 13944 5936 14754 5947
rect 14810 5936 15510 5947
rect 15938 6000 17504 6008
rect 15938 5987 16748 6000
rect 16804 5987 17504 6000
rect 15938 5953 16061 5987
rect 16095 5953 16153 5987
rect 16187 5953 16245 5987
rect 16279 5953 16337 5987
rect 16371 5953 16429 5987
rect 16463 5953 16521 5987
rect 16555 5953 16613 5987
rect 16647 5953 16705 5987
rect 16739 5953 16748 5987
rect 16831 5953 16889 5987
rect 16923 5953 16981 5987
rect 17015 5953 17073 5987
rect 17107 5953 17165 5987
rect 17199 5953 17257 5987
rect 17291 5953 17349 5987
rect 17383 5953 17441 5987
rect 17475 5953 17504 5987
rect 15938 5942 16748 5953
rect 16804 5942 17504 5953
rect 13944 5930 15510 5936
rect 10214 5747 10272 5753
rect 10214 5713 10226 5747
rect 10260 5744 10272 5747
rect 10300 5744 10328 5920
rect 12080 5908 13552 5928
rect 14038 5916 15510 5930
rect 16032 5922 17504 5942
rect 10398 5815 10456 5821
rect 10398 5781 10410 5815
rect 10444 5812 10456 5815
rect 11138 5815 11196 5821
rect 11138 5812 11150 5815
rect 10444 5784 11150 5812
rect 10444 5781 10456 5784
rect 10398 5775 10456 5781
rect 11138 5781 11150 5784
rect 11184 5781 11196 5815
rect 11138 5775 11196 5781
rect 10582 5747 10640 5753
rect 10582 5744 10594 5747
rect 10260 5716 10594 5744
rect 10260 5713 10272 5716
rect 10214 5707 10272 5713
rect 10582 5713 10594 5716
rect 10628 5744 10640 5747
rect 10954 5747 11012 5753
rect 10954 5744 10966 5747
rect 10628 5716 10966 5744
rect 10628 5713 10640 5716
rect 10582 5707 10640 5713
rect 10954 5713 10966 5716
rect 11000 5744 11012 5747
rect 11230 5747 11288 5753
rect 11230 5744 11242 5747
rect 11000 5716 11242 5744
rect 11000 5713 11012 5716
rect 10954 5707 11012 5713
rect 11230 5713 11242 5716
rect 11276 5713 11288 5747
rect 11230 5707 11288 5713
rect 12276 5735 12334 5741
rect 12276 5701 12288 5735
rect 12322 5732 12334 5735
rect 12362 5732 12390 5908
rect 12460 5803 12518 5809
rect 12460 5769 12472 5803
rect 12506 5800 12518 5803
rect 13200 5803 13258 5809
rect 13200 5800 13212 5803
rect 12506 5772 13212 5800
rect 12506 5769 12518 5772
rect 12460 5763 12518 5769
rect 13200 5769 13212 5772
rect 13246 5769 13258 5803
rect 13200 5763 13258 5769
rect 14234 5743 14292 5749
rect 12644 5735 12702 5741
rect 12644 5732 12656 5735
rect 12322 5704 12656 5732
rect 12322 5701 12334 5704
rect 12276 5695 12334 5701
rect 12644 5701 12656 5704
rect 12690 5732 12702 5735
rect 13016 5735 13074 5741
rect 13016 5732 13028 5735
rect 12690 5704 13028 5732
rect 12690 5701 12702 5704
rect 12644 5695 12702 5701
rect 13016 5701 13028 5704
rect 13062 5732 13074 5735
rect 13292 5735 13350 5741
rect 13292 5732 13304 5735
rect 13062 5704 13304 5732
rect 13062 5701 13074 5704
rect 13016 5695 13074 5701
rect 13292 5701 13304 5704
rect 13338 5701 13350 5735
rect 14234 5709 14246 5743
rect 14280 5740 14292 5743
rect 14320 5740 14348 5916
rect 14418 5811 14476 5817
rect 14418 5777 14430 5811
rect 14464 5808 14476 5811
rect 15158 5811 15216 5817
rect 15158 5808 15170 5811
rect 14464 5780 15170 5808
rect 14464 5777 14476 5780
rect 14418 5771 14476 5777
rect 15158 5777 15170 5780
rect 15204 5777 15216 5811
rect 15158 5771 15216 5777
rect 16228 5749 16286 5755
rect 14602 5743 14660 5749
rect 14602 5740 14614 5743
rect 14280 5712 14614 5740
rect 14280 5709 14292 5712
rect 14234 5703 14292 5709
rect 14602 5709 14614 5712
rect 14648 5740 14660 5743
rect 14974 5743 15032 5749
rect 14974 5740 14986 5743
rect 14648 5712 14986 5740
rect 14648 5709 14660 5712
rect 14602 5703 14660 5709
rect 14974 5709 14986 5712
rect 15020 5740 15032 5743
rect 15250 5743 15308 5749
rect 15250 5740 15262 5743
rect 15020 5712 15262 5740
rect 15020 5709 15032 5712
rect 14974 5703 15032 5709
rect 15250 5709 15262 5712
rect 15296 5709 15308 5743
rect 16228 5715 16240 5749
rect 16274 5746 16286 5749
rect 16314 5746 16342 5922
rect 16412 5817 16470 5823
rect 16412 5783 16424 5817
rect 16458 5814 16470 5817
rect 17152 5817 17210 5823
rect 17152 5814 17164 5817
rect 16458 5786 17164 5814
rect 16458 5783 16470 5786
rect 16412 5777 16470 5783
rect 17152 5783 17164 5786
rect 17198 5783 17210 5817
rect 17152 5777 17210 5783
rect 16596 5749 16654 5755
rect 16596 5746 16608 5749
rect 16274 5718 16608 5746
rect 16274 5715 16286 5718
rect 16228 5709 16286 5715
rect 16596 5715 16608 5718
rect 16642 5746 16654 5749
rect 16968 5749 17026 5755
rect 16968 5746 16980 5749
rect 16642 5718 16980 5746
rect 16642 5715 16654 5718
rect 16596 5709 16654 5715
rect 16968 5715 16980 5718
rect 17014 5746 17026 5749
rect 17244 5749 17302 5755
rect 17244 5746 17256 5749
rect 17014 5718 17256 5746
rect 17014 5715 17026 5718
rect 16968 5709 17026 5715
rect 17244 5715 17256 5718
rect 17290 5715 17302 5749
rect 17244 5709 17302 5715
rect 15250 5703 15308 5709
rect 13292 5695 13350 5701
rect 10306 5679 10364 5685
rect 10306 5645 10318 5679
rect 10352 5676 10364 5679
rect 10766 5679 10824 5685
rect 10766 5676 10778 5679
rect 10352 5648 10778 5676
rect 10352 5645 10364 5648
rect 10306 5639 10364 5645
rect 10766 5645 10778 5648
rect 10812 5676 10824 5679
rect 11138 5679 11196 5685
rect 16320 5681 16378 5687
rect 11138 5676 11150 5679
rect 10812 5648 11150 5676
rect 10812 5645 10824 5648
rect 10766 5639 10824 5645
rect 10404 5618 10470 5620
rect 1836 5590 3308 5596
rect 1736 5578 3308 5590
rect 1736 5565 2564 5578
rect 2620 5565 3308 5578
rect 3970 5576 5442 5588
rect 5922 5584 7394 5588
rect 1736 5531 1865 5565
rect 1899 5531 1957 5565
rect 1991 5531 2049 5565
rect 2083 5531 2141 5565
rect 2175 5531 2233 5565
rect 2267 5531 2325 5565
rect 2359 5531 2417 5565
rect 2451 5531 2509 5565
rect 2543 5531 2564 5565
rect 2635 5531 2693 5565
rect 2727 5531 2785 5565
rect 2819 5531 2877 5565
rect 2911 5531 2969 5565
rect 3003 5531 3061 5565
rect 3095 5531 3153 5565
rect 3187 5531 3245 5565
rect 3279 5531 3308 5565
rect 1736 5524 2564 5531
rect 1836 5520 2564 5524
rect 2620 5520 3308 5531
rect 1836 5500 3308 5520
rect 3904 5570 5442 5576
rect 3904 5557 4686 5570
rect 4742 5557 5442 5570
rect 3904 5523 3999 5557
rect 4033 5523 4091 5557
rect 4125 5523 4183 5557
rect 4217 5523 4275 5557
rect 4309 5523 4367 5557
rect 4401 5523 4459 5557
rect 4493 5523 4551 5557
rect 4585 5523 4643 5557
rect 4677 5523 4686 5557
rect 4769 5523 4827 5557
rect 4861 5523 4919 5557
rect 4953 5523 5011 5557
rect 5045 5523 5103 5557
rect 5137 5523 5195 5557
rect 5229 5523 5287 5557
rect 5321 5523 5379 5557
rect 5413 5523 5442 5557
rect 3904 5512 4686 5523
rect 4742 5512 5442 5523
rect 5848 5570 7394 5584
rect 7924 5582 9396 5594
rect 5848 5557 6638 5570
rect 6694 5557 7394 5570
rect 5848 5523 5951 5557
rect 5985 5523 6043 5557
rect 6077 5523 6135 5557
rect 6169 5523 6227 5557
rect 6261 5523 6319 5557
rect 6353 5523 6411 5557
rect 6445 5523 6503 5557
rect 6537 5523 6595 5557
rect 6629 5523 6638 5557
rect 6721 5523 6779 5557
rect 6813 5523 6871 5557
rect 6905 5523 6963 5557
rect 6997 5523 7055 5557
rect 7089 5523 7147 5557
rect 7181 5523 7239 5557
rect 7273 5523 7331 5557
rect 7365 5523 7394 5557
rect 5848 5518 6638 5523
rect 3904 5510 5442 5512
rect 2032 5327 2090 5333
rect 2032 5293 2044 5327
rect 2078 5324 2090 5327
rect 2118 5324 2146 5500
rect 3970 5492 5442 5510
rect 5922 5512 6638 5518
rect 6694 5512 7394 5523
rect 7850 5576 9396 5582
rect 7850 5563 8640 5576
rect 8696 5563 9396 5576
rect 7850 5529 7953 5563
rect 7987 5529 8045 5563
rect 8079 5529 8137 5563
rect 8171 5529 8229 5563
rect 8263 5529 8321 5563
rect 8355 5529 8413 5563
rect 8447 5529 8505 5563
rect 8539 5529 8597 5563
rect 8631 5529 8640 5563
rect 8723 5529 8781 5563
rect 8815 5529 8873 5563
rect 8907 5529 8965 5563
rect 8999 5529 9057 5563
rect 9091 5529 9149 5563
rect 9183 5529 9241 5563
rect 9275 5529 9333 5563
rect 9367 5529 9396 5563
rect 10404 5566 10410 5618
rect 10462 5566 10470 5618
rect 10404 5562 10470 5566
rect 7850 5518 8640 5529
rect 8696 5518 9396 5529
rect 7850 5516 9396 5518
rect 5922 5492 7394 5512
rect 7924 5498 9396 5516
rect 2216 5395 2274 5401
rect 2216 5361 2228 5395
rect 2262 5392 2274 5395
rect 2956 5395 3014 5401
rect 2956 5392 2968 5395
rect 2262 5364 2968 5392
rect 2262 5361 2274 5364
rect 2216 5355 2274 5361
rect 2956 5361 2968 5364
rect 3002 5361 3014 5395
rect 2956 5355 3014 5361
rect 2400 5327 2458 5333
rect 2400 5324 2412 5327
rect 2078 5296 2412 5324
rect 2078 5293 2090 5296
rect 2032 5287 2090 5293
rect 2400 5293 2412 5296
rect 2446 5324 2458 5327
rect 2772 5327 2830 5333
rect 2772 5324 2784 5327
rect 2446 5296 2784 5324
rect 2446 5293 2458 5296
rect 2400 5287 2458 5293
rect 2772 5293 2784 5296
rect 2818 5324 2830 5327
rect 3048 5327 3106 5333
rect 3048 5324 3060 5327
rect 2818 5296 3060 5324
rect 2818 5293 2830 5296
rect 2772 5287 2830 5293
rect 3048 5293 3060 5296
rect 3094 5293 3106 5327
rect 3048 5287 3106 5293
rect 4166 5319 4224 5325
rect 4166 5285 4178 5319
rect 4212 5316 4224 5319
rect 4252 5316 4280 5492
rect 4350 5387 4408 5393
rect 4350 5353 4362 5387
rect 4396 5384 4408 5387
rect 5090 5387 5148 5393
rect 5090 5384 5102 5387
rect 4396 5356 5102 5384
rect 4396 5353 4408 5356
rect 4350 5347 4408 5353
rect 5090 5353 5102 5356
rect 5136 5353 5148 5387
rect 5090 5347 5148 5353
rect 4534 5319 4592 5325
rect 4534 5316 4546 5319
rect 4212 5288 4546 5316
rect 4212 5285 4224 5288
rect 4166 5279 4224 5285
rect 4534 5285 4546 5288
rect 4580 5316 4592 5319
rect 4906 5319 4964 5325
rect 4906 5316 4918 5319
rect 4580 5288 4918 5316
rect 4580 5285 4592 5288
rect 4534 5279 4592 5285
rect 4906 5285 4918 5288
rect 4952 5316 4964 5319
rect 5182 5319 5240 5325
rect 5182 5316 5194 5319
rect 4952 5288 5194 5316
rect 4952 5285 4964 5288
rect 4906 5279 4964 5285
rect 5182 5285 5194 5288
rect 5228 5285 5240 5319
rect 5182 5279 5240 5285
rect 6118 5319 6176 5325
rect 6118 5285 6130 5319
rect 6164 5316 6176 5319
rect 6204 5316 6232 5492
rect 6302 5387 6360 5393
rect 6302 5353 6314 5387
rect 6348 5384 6360 5387
rect 7042 5387 7100 5393
rect 7042 5384 7054 5387
rect 6348 5356 7054 5384
rect 6348 5353 6360 5356
rect 6302 5347 6360 5353
rect 7042 5353 7054 5356
rect 7088 5353 7100 5387
rect 7042 5347 7100 5353
rect 8120 5325 8178 5331
rect 6486 5319 6544 5325
rect 6486 5316 6498 5319
rect 6164 5288 6498 5316
rect 6164 5285 6176 5288
rect 6118 5279 6176 5285
rect 6486 5285 6498 5288
rect 6532 5316 6544 5319
rect 6858 5319 6916 5325
rect 6858 5316 6870 5319
rect 6532 5288 6870 5316
rect 6532 5285 6544 5288
rect 6486 5279 6544 5285
rect 6858 5285 6870 5288
rect 6904 5316 6916 5319
rect 7134 5319 7192 5325
rect 7134 5316 7146 5319
rect 6904 5288 7146 5316
rect 6904 5285 6916 5288
rect 6858 5279 6916 5285
rect 7134 5285 7146 5288
rect 7180 5285 7192 5319
rect 8120 5291 8132 5325
rect 8166 5322 8178 5325
rect 8206 5322 8234 5498
rect 10860 5472 10888 5648
rect 11138 5645 11150 5648
rect 11184 5645 11196 5679
rect 14326 5675 14384 5681
rect 11138 5639 11196 5645
rect 12368 5667 12426 5673
rect 12368 5633 12380 5667
rect 12414 5664 12426 5667
rect 12828 5667 12886 5673
rect 12828 5664 12840 5667
rect 12414 5636 12840 5664
rect 12414 5633 12426 5636
rect 11412 5606 11472 5630
rect 12368 5627 12426 5633
rect 12828 5633 12840 5636
rect 12874 5664 12886 5667
rect 13200 5667 13258 5673
rect 13200 5664 13212 5667
rect 12874 5636 13212 5664
rect 12874 5633 12886 5636
rect 12828 5627 12886 5633
rect 11412 5570 11426 5606
rect 11466 5604 11472 5606
rect 11466 5596 11818 5604
rect 12464 5600 12524 5606
rect 12464 5596 12478 5600
rect 11466 5570 12478 5596
rect 11412 5566 12478 5570
rect 12512 5566 12524 5600
rect 11412 5554 11472 5566
rect 11804 5562 12524 5566
rect 11896 5558 12524 5562
rect 12464 5544 12524 5558
rect 10018 5460 11490 5472
rect 12922 5460 12950 5636
rect 13200 5633 13212 5636
rect 13246 5633 13258 5667
rect 14326 5641 14338 5675
rect 14372 5672 14384 5675
rect 14786 5675 14844 5681
rect 14786 5672 14798 5675
rect 14372 5644 14798 5672
rect 14372 5641 14384 5644
rect 14326 5635 14384 5641
rect 14786 5641 14798 5644
rect 14832 5672 14844 5675
rect 15158 5675 15216 5681
rect 15158 5672 15170 5675
rect 14832 5644 15170 5672
rect 14832 5641 14844 5644
rect 14786 5635 14844 5641
rect 13200 5627 13258 5633
rect 13482 5594 13534 5612
rect 14422 5608 14482 5614
rect 14422 5604 14436 5608
rect 13565 5594 14436 5604
rect 13480 5558 13494 5594
rect 13528 5574 14436 5594
rect 14470 5574 14482 5608
rect 13528 5566 14482 5574
rect 13528 5558 13588 5566
rect 13480 5556 13588 5558
rect 13482 5546 13534 5556
rect 14422 5552 14482 5566
rect 14880 5468 14908 5644
rect 15158 5641 15170 5644
rect 15204 5641 15216 5675
rect 16320 5647 16332 5681
rect 16366 5678 16378 5681
rect 16780 5681 16838 5687
rect 16780 5678 16792 5681
rect 16366 5650 16792 5678
rect 16366 5647 16378 5650
rect 16320 5641 16378 5647
rect 16780 5647 16792 5650
rect 16826 5678 16838 5681
rect 17152 5681 17210 5687
rect 17152 5678 17164 5681
rect 16826 5650 17164 5678
rect 16826 5647 16838 5650
rect 16780 5641 16838 5647
rect 15158 5635 15216 5641
rect 15440 5602 15492 5620
rect 16416 5614 16476 5620
rect 16416 5610 16430 5614
rect 15848 5606 16430 5610
rect 15524 5602 16430 5606
rect 15438 5566 15452 5602
rect 15486 5580 16430 5602
rect 16464 5580 16476 5614
rect 15486 5572 16476 5580
rect 15486 5566 15884 5572
rect 15438 5564 15884 5566
rect 15440 5554 15492 5564
rect 16416 5558 16476 5572
rect 16874 5474 16902 5650
rect 17152 5647 17164 5650
rect 17198 5647 17210 5681
rect 17152 5641 17210 5647
rect 17434 5608 17486 5626
rect 17432 5572 17446 5608
rect 17480 5596 17540 5608
rect 17480 5572 17822 5596
rect 17432 5570 17822 5572
rect 17434 5564 17822 5570
rect 17434 5560 17514 5564
rect 9940 5452 11490 5460
rect 9940 5441 11214 5452
rect 11270 5441 11490 5452
rect 12080 5444 13552 5460
rect 14038 5458 15510 5468
rect 16032 5460 17504 5474
rect 9940 5407 10047 5441
rect 10081 5407 10139 5441
rect 10173 5407 10231 5441
rect 10265 5407 10323 5441
rect 10357 5407 10415 5441
rect 10449 5407 10507 5441
rect 10541 5407 10599 5441
rect 10633 5407 10691 5441
rect 10725 5407 10783 5441
rect 10817 5407 10875 5441
rect 10909 5407 10967 5441
rect 11001 5407 11059 5441
rect 11093 5407 11151 5441
rect 11185 5407 11214 5441
rect 11277 5407 11335 5441
rect 11369 5407 11427 5441
rect 11461 5407 11490 5441
rect 8304 5393 8362 5399
rect 8304 5359 8316 5393
rect 8350 5390 8362 5393
rect 9044 5393 9102 5399
rect 9940 5394 11214 5407
rect 11270 5394 11490 5407
rect 9044 5390 9056 5393
rect 8350 5362 9056 5390
rect 8350 5359 8362 5362
rect 8304 5353 8362 5359
rect 9044 5359 9056 5362
rect 9090 5359 9102 5393
rect 10018 5376 11490 5394
rect 12002 5440 13552 5444
rect 12002 5429 12800 5440
rect 12856 5429 13552 5440
rect 12002 5395 12109 5429
rect 12143 5395 12201 5429
rect 12235 5395 12293 5429
rect 12327 5395 12385 5429
rect 12419 5395 12477 5429
rect 12511 5395 12569 5429
rect 12603 5395 12661 5429
rect 12695 5395 12753 5429
rect 12787 5395 12800 5429
rect 12879 5395 12937 5429
rect 12971 5395 13029 5429
rect 13063 5395 13121 5429
rect 13155 5395 13213 5429
rect 13247 5395 13305 5429
rect 13339 5395 13397 5429
rect 13431 5395 13489 5429
rect 13523 5395 13552 5429
rect 12002 5382 12800 5395
rect 12856 5382 13552 5395
rect 13950 5448 15510 5458
rect 13950 5437 14758 5448
rect 14814 5437 15510 5448
rect 13950 5403 14067 5437
rect 14101 5403 14159 5437
rect 14193 5403 14251 5437
rect 14285 5403 14343 5437
rect 14377 5403 14435 5437
rect 14469 5403 14527 5437
rect 14561 5403 14619 5437
rect 14653 5403 14711 5437
rect 14745 5403 14758 5437
rect 14837 5403 14895 5437
rect 14929 5403 14987 5437
rect 15021 5403 15079 5437
rect 15113 5403 15171 5437
rect 15205 5403 15263 5437
rect 15297 5403 15355 5437
rect 15389 5403 15447 5437
rect 15481 5403 15510 5437
rect 13950 5392 14758 5403
rect 12002 5378 13552 5382
rect 12080 5364 13552 5378
rect 14038 5390 14758 5392
rect 14814 5390 15510 5403
rect 15946 5454 17504 5460
rect 15946 5443 16752 5454
rect 16808 5443 17504 5454
rect 15946 5409 16061 5443
rect 16095 5409 16153 5443
rect 16187 5409 16245 5443
rect 16279 5409 16337 5443
rect 16371 5409 16429 5443
rect 16463 5409 16521 5443
rect 16555 5409 16613 5443
rect 16647 5409 16705 5443
rect 16739 5409 16752 5443
rect 16831 5409 16889 5443
rect 16923 5409 16981 5443
rect 17015 5409 17073 5443
rect 17107 5409 17165 5443
rect 17199 5409 17257 5443
rect 17291 5409 17349 5443
rect 17383 5409 17441 5443
rect 17475 5409 17504 5443
rect 15946 5396 16752 5409
rect 16808 5396 17504 5409
rect 15946 5394 17504 5396
rect 14038 5372 15510 5390
rect 16032 5378 17504 5394
rect 9044 5353 9102 5359
rect 8488 5325 8546 5331
rect 8488 5322 8500 5325
rect 8166 5294 8500 5322
rect 8166 5291 8178 5294
rect 8120 5285 8178 5291
rect 8488 5291 8500 5294
rect 8534 5322 8546 5325
rect 8860 5325 8918 5331
rect 8860 5322 8872 5325
rect 8534 5294 8872 5322
rect 8534 5291 8546 5294
rect 8488 5285 8546 5291
rect 8860 5291 8872 5294
rect 8906 5322 8918 5325
rect 9136 5325 9194 5331
rect 9136 5322 9148 5325
rect 8906 5294 9148 5322
rect 8906 5291 8918 5294
rect 8860 5285 8918 5291
rect 9136 5291 9148 5294
rect 9182 5291 9194 5325
rect 9136 5285 9194 5291
rect 17790 5302 17822 5564
rect 19106 5374 19226 5440
rect 7134 5279 7192 5285
rect 17790 5270 18732 5302
rect 2124 5259 2182 5265
rect 2124 5225 2136 5259
rect 2170 5256 2182 5259
rect 2584 5259 2642 5265
rect 2584 5256 2596 5259
rect 2170 5228 2596 5256
rect 2170 5225 2182 5228
rect 2124 5219 2182 5225
rect 2584 5225 2596 5228
rect 2630 5256 2642 5259
rect 2956 5259 3014 5265
rect 2956 5256 2968 5259
rect 2630 5228 2968 5256
rect 2630 5225 2642 5228
rect 2584 5219 2642 5225
rect 2222 5198 2288 5200
rect 2222 5146 2228 5198
rect 2280 5146 2288 5198
rect 2222 5142 2288 5146
rect 2678 5052 2706 5228
rect 2956 5225 2968 5228
rect 3002 5225 3014 5259
rect 8212 5257 8270 5263
rect 2956 5219 3014 5225
rect 4258 5251 4316 5257
rect 4258 5217 4270 5251
rect 4304 5248 4316 5251
rect 4718 5251 4776 5257
rect 4718 5248 4730 5251
rect 4304 5220 4730 5248
rect 4304 5217 4316 5220
rect 4258 5211 4316 5217
rect 4718 5217 4730 5220
rect 4764 5248 4776 5251
rect 5090 5251 5148 5257
rect 5090 5248 5102 5251
rect 4764 5220 5102 5248
rect 4764 5217 4776 5220
rect 4718 5211 4776 5217
rect 3230 5186 3290 5210
rect 3230 5150 3244 5186
rect 3284 5184 3290 5186
rect 4354 5184 4414 5190
rect 3284 5180 3837 5184
rect 4354 5180 4368 5184
rect 3284 5150 4368 5180
rect 4402 5150 4414 5184
rect 3230 5146 4414 5150
rect 3230 5134 3290 5146
rect 3636 5142 4414 5146
rect 4354 5128 4414 5142
rect 1836 5040 3308 5052
rect 4812 5044 4840 5220
rect 5090 5217 5102 5220
rect 5136 5217 5148 5251
rect 5090 5211 5148 5217
rect 6210 5251 6268 5257
rect 6210 5217 6222 5251
rect 6256 5248 6268 5251
rect 6670 5251 6728 5257
rect 6670 5248 6682 5251
rect 6256 5220 6682 5248
rect 6256 5217 6268 5220
rect 6210 5211 6268 5217
rect 6670 5217 6682 5220
rect 6716 5248 6728 5251
rect 7042 5251 7100 5257
rect 7042 5248 7054 5251
rect 6716 5220 7054 5248
rect 6716 5217 6728 5220
rect 6670 5211 6728 5217
rect 5372 5178 5424 5196
rect 6306 5184 6366 5190
rect 6306 5180 6320 5184
rect 5612 5178 6320 5180
rect 5370 5142 5384 5178
rect 5418 5150 6320 5178
rect 6354 5150 6366 5184
rect 5418 5142 6366 5150
rect 5370 5140 5659 5142
rect 5372 5130 5424 5140
rect 6306 5128 6366 5142
rect 6764 5044 6792 5220
rect 7042 5217 7054 5220
rect 7088 5217 7100 5251
rect 8212 5223 8224 5257
rect 8258 5254 8270 5257
rect 8672 5257 8730 5263
rect 8672 5254 8684 5257
rect 8258 5226 8684 5254
rect 8258 5223 8270 5226
rect 8212 5217 8270 5223
rect 8672 5223 8684 5226
rect 8718 5254 8730 5257
rect 9044 5257 9102 5263
rect 9044 5254 9056 5257
rect 8718 5226 9056 5254
rect 8718 5223 8730 5226
rect 8672 5217 8730 5223
rect 7042 5211 7100 5217
rect 7324 5178 7376 5196
rect 8308 5190 8368 5196
rect 8308 5186 8322 5190
rect 7550 5178 8322 5186
rect 7322 5142 7336 5178
rect 7370 5156 8322 5178
rect 8356 5156 8368 5190
rect 7370 5148 8368 5156
rect 7370 5142 7611 5148
rect 7322 5140 7611 5142
rect 7324 5130 7376 5140
rect 8308 5134 8368 5148
rect 8766 5050 8794 5226
rect 9044 5223 9056 5226
rect 9090 5223 9102 5257
rect 9044 5217 9102 5223
rect 9906 5210 17524 5242
rect 9326 5184 9378 5202
rect 9906 5184 9938 5210
rect 9324 5148 9338 5184
rect 9372 5148 9938 5184
rect 9324 5146 9938 5148
rect 9326 5136 9378 5146
rect 9762 5144 9938 5146
rect 17492 5146 17524 5210
rect 18598 5222 18648 5242
rect 18598 5188 18608 5222
rect 18642 5188 18648 5222
rect 10046 5138 11518 5142
rect 10046 5120 11614 5138
rect 10046 5111 10188 5120
rect 10244 5111 11614 5120
rect 17492 5114 18178 5146
rect 18598 5134 18648 5188
rect 18678 5194 18732 5270
rect 18678 5160 18690 5194
rect 18724 5160 18732 5194
rect 10046 5077 10075 5111
rect 10109 5077 10167 5111
rect 10244 5077 10259 5111
rect 10293 5077 10351 5111
rect 10385 5077 10443 5111
rect 10477 5077 10535 5111
rect 10569 5077 10627 5111
rect 10661 5077 10719 5111
rect 10753 5077 10811 5111
rect 10845 5077 10903 5111
rect 10937 5077 10995 5111
rect 11029 5077 11087 5111
rect 11121 5077 11179 5111
rect 11213 5077 11271 5111
rect 11305 5077 11363 5111
rect 11397 5077 11455 5111
rect 11489 5077 11614 5111
rect 18146 5102 18178 5114
rect 18426 5108 18480 5120
rect 18250 5102 18432 5108
rect 12316 5088 13788 5098
rect 10046 5062 10188 5077
rect 10244 5072 11614 5077
rect 12234 5080 13788 5088
rect 14318 5082 15790 5092
rect 10244 5062 11518 5072
rect 7924 5044 9396 5050
rect 10046 5046 11518 5062
rect 12234 5067 13032 5080
rect 13088 5067 13788 5080
rect 1836 5036 2584 5040
rect 1750 5021 2584 5036
rect 2640 5021 3308 5040
rect 3970 5036 5442 5044
rect 1750 4987 1865 5021
rect 1899 4987 1957 5021
rect 1991 4987 2049 5021
rect 2083 4987 2141 5021
rect 2175 4987 2233 5021
rect 2267 4987 2325 5021
rect 2359 4987 2417 5021
rect 2451 4987 2509 5021
rect 2543 4987 2584 5021
rect 2640 4987 2693 5021
rect 2727 4987 2785 5021
rect 2819 4987 2877 5021
rect 2911 4987 2969 5021
rect 3003 4987 3061 5021
rect 3095 4987 3153 5021
rect 3187 4987 3245 5021
rect 3279 4987 3308 5021
rect 1750 4982 2584 4987
rect 2640 4982 3308 4987
rect 1750 4970 3308 4982
rect 3884 5024 5442 5036
rect 5922 5030 7394 5044
rect 3884 5013 4690 5024
rect 4746 5013 5442 5024
rect 3884 4979 3999 5013
rect 4033 4979 4091 5013
rect 4125 4979 4183 5013
rect 4217 4979 4275 5013
rect 4309 4979 4367 5013
rect 4401 4979 4459 5013
rect 4493 4979 4551 5013
rect 4585 4979 4643 5013
rect 4677 4979 4690 5013
rect 4769 4979 4827 5013
rect 4861 4979 4919 5013
rect 4953 4979 5011 5013
rect 5045 4979 5103 5013
rect 5137 4979 5195 5013
rect 5229 4979 5287 5013
rect 5321 4979 5379 5013
rect 5413 4979 5442 5013
rect 3884 4970 4690 4979
rect 1836 4956 3308 4970
rect 3970 4966 4690 4970
rect 4746 4966 5442 4979
rect 3970 4948 5442 4966
rect 5836 5024 7394 5030
rect 5836 5013 6642 5024
rect 6698 5013 7394 5024
rect 5836 4979 5951 5013
rect 5985 4979 6043 5013
rect 6077 4979 6135 5013
rect 6169 4979 6227 5013
rect 6261 4979 6319 5013
rect 6353 4979 6411 5013
rect 6445 4979 6503 5013
rect 6537 4979 6595 5013
rect 6629 4979 6642 5013
rect 6721 4979 6779 5013
rect 6813 4979 6871 5013
rect 6905 4979 6963 5013
rect 6997 4979 7055 5013
rect 7089 4979 7147 5013
rect 7181 4979 7239 5013
rect 7273 4979 7331 5013
rect 7365 4979 7394 5013
rect 5836 4966 6642 4979
rect 6698 4966 7394 4979
rect 7848 5030 9396 5044
rect 7848 5019 8644 5030
rect 8700 5019 9396 5030
rect 7848 4985 7953 5019
rect 7987 4985 8045 5019
rect 8079 4985 8137 5019
rect 8171 4985 8229 5019
rect 8263 4985 8321 5019
rect 8355 4985 8413 5019
rect 8447 4985 8505 5019
rect 8539 4985 8597 5019
rect 8631 4985 8644 5019
rect 8723 4985 8781 5019
rect 8815 4985 8873 5019
rect 8907 4985 8965 5019
rect 8999 4985 9057 5019
rect 9091 4985 9149 5019
rect 9183 4985 9241 5019
rect 9275 4985 9333 5019
rect 9367 4985 9396 5019
rect 7848 4978 8644 4985
rect 5836 4964 7394 4966
rect 5922 4948 7394 4964
rect 7924 4972 8644 4978
rect 8700 4972 9396 4985
rect 7924 4954 9396 4972
rect 10242 4873 10300 4879
rect 10242 4839 10254 4873
rect 10288 4870 10300 4873
rect 10328 4870 10356 5046
rect 12234 5033 12345 5067
rect 12379 5033 12437 5067
rect 12471 5033 12529 5067
rect 12563 5033 12621 5067
rect 12655 5033 12713 5067
rect 12747 5033 12805 5067
rect 12839 5033 12897 5067
rect 12931 5033 12989 5067
rect 13023 5033 13032 5067
rect 13115 5033 13173 5067
rect 13207 5033 13265 5067
rect 13299 5033 13357 5067
rect 13391 5033 13449 5067
rect 13483 5033 13541 5067
rect 13575 5033 13633 5067
rect 13667 5033 13725 5067
rect 13759 5033 13788 5067
rect 12234 5022 13032 5033
rect 13088 5022 13788 5033
rect 12316 5002 13788 5022
rect 14240 5074 15790 5082
rect 14240 5061 15034 5074
rect 15090 5061 15790 5074
rect 14240 5027 14347 5061
rect 14381 5027 14439 5061
rect 14473 5027 14531 5061
rect 14565 5027 14623 5061
rect 14657 5027 14715 5061
rect 14749 5027 14807 5061
rect 14841 5027 14899 5061
rect 14933 5027 14991 5061
rect 15025 5027 15034 5061
rect 15117 5027 15175 5061
rect 15209 5027 15267 5061
rect 15301 5027 15359 5061
rect 15393 5027 15451 5061
rect 15485 5027 15543 5061
rect 15577 5027 15635 5061
rect 15669 5027 15727 5061
rect 15761 5027 15790 5061
rect 16340 5058 17812 5074
rect 18146 5070 18432 5102
rect 18470 5070 18572 5108
rect 14240 5016 15034 5027
rect 15090 5016 15790 5027
rect 10426 4941 10484 4947
rect 10426 4907 10438 4941
rect 10472 4938 10484 4941
rect 11166 4941 11224 4947
rect 11166 4938 11178 4941
rect 10472 4910 11178 4938
rect 10472 4907 10484 4910
rect 10426 4901 10484 4907
rect 11166 4907 11178 4910
rect 11212 4907 11224 4941
rect 11166 4901 11224 4907
rect 10610 4873 10668 4879
rect 10610 4870 10622 4873
rect 10288 4842 10622 4870
rect 10288 4839 10300 4842
rect 10242 4833 10300 4839
rect 10610 4839 10622 4842
rect 10656 4870 10668 4873
rect 10982 4873 11040 4879
rect 10982 4870 10994 4873
rect 10656 4842 10994 4870
rect 10656 4839 10668 4842
rect 10610 4833 10668 4839
rect 10982 4839 10994 4842
rect 11028 4870 11040 4873
rect 11258 4873 11316 4879
rect 11258 4870 11270 4873
rect 11028 4842 11270 4870
rect 11028 4839 11040 4842
rect 10982 4833 11040 4839
rect 11258 4839 11270 4842
rect 11304 4839 11316 4873
rect 11258 4833 11316 4839
rect 12512 4829 12570 4835
rect 10334 4805 10392 4811
rect 10334 4771 10346 4805
rect 10380 4802 10392 4805
rect 10794 4805 10852 4811
rect 10794 4802 10806 4805
rect 10380 4774 10806 4802
rect 10380 4771 10392 4774
rect 10334 4765 10392 4771
rect 10794 4771 10806 4774
rect 10840 4802 10852 4805
rect 11166 4805 11224 4811
rect 11166 4802 11178 4805
rect 10840 4774 11178 4802
rect 10840 4771 10852 4774
rect 10794 4765 10852 4771
rect 10432 4744 10498 4746
rect 10432 4692 10438 4744
rect 10490 4692 10498 4744
rect 10432 4688 10498 4692
rect 10888 4598 10916 4774
rect 11166 4771 11178 4774
rect 11212 4771 11224 4805
rect 12512 4795 12524 4829
rect 12558 4826 12570 4829
rect 12598 4826 12626 5002
rect 14318 4996 15790 5016
rect 16272 5056 17812 5058
rect 16272 5043 17056 5056
rect 17112 5043 17812 5056
rect 18426 5054 18480 5070
rect 16272 5009 16369 5043
rect 16403 5009 16461 5043
rect 16495 5009 16553 5043
rect 16587 5009 16645 5043
rect 16679 5009 16737 5043
rect 16771 5009 16829 5043
rect 16863 5009 16921 5043
rect 16955 5009 17013 5043
rect 17047 5009 17056 5043
rect 17139 5009 17197 5043
rect 17231 5009 17289 5043
rect 17323 5009 17381 5043
rect 17415 5009 17473 5043
rect 17507 5009 17565 5043
rect 17599 5009 17657 5043
rect 17691 5009 17749 5043
rect 17783 5009 17812 5043
rect 18608 5024 18640 5134
rect 18678 5114 18732 5160
rect 18678 5110 18716 5114
rect 18250 5023 18640 5024
rect 16272 4998 17056 5009
rect 17112 4998 17812 5009
rect 12696 4897 12754 4903
rect 12696 4863 12708 4897
rect 12742 4894 12754 4897
rect 13436 4897 13494 4903
rect 13436 4894 13448 4897
rect 12742 4866 13448 4894
rect 12742 4863 12754 4866
rect 12696 4857 12754 4863
rect 13436 4863 13448 4866
rect 13482 4863 13494 4897
rect 13436 4857 13494 4863
rect 12880 4829 12938 4835
rect 12880 4826 12892 4829
rect 12558 4798 12892 4826
rect 12558 4795 12570 4798
rect 12512 4789 12570 4795
rect 12880 4795 12892 4798
rect 12926 4826 12938 4829
rect 13252 4829 13310 4835
rect 13252 4826 13264 4829
rect 12926 4798 13264 4826
rect 12926 4795 12938 4798
rect 12880 4789 12938 4795
rect 13252 4795 13264 4798
rect 13298 4826 13310 4829
rect 13528 4829 13586 4835
rect 13528 4826 13540 4829
rect 13298 4798 13540 4826
rect 13298 4795 13310 4798
rect 13252 4789 13310 4795
rect 13528 4795 13540 4798
rect 13574 4795 13586 4829
rect 13528 4789 13586 4795
rect 14514 4823 14572 4829
rect 14514 4789 14526 4823
rect 14560 4820 14572 4823
rect 14600 4820 14628 4996
rect 16272 4992 17812 4998
rect 16340 4978 17812 4992
rect 18169 4992 18640 5023
rect 19046 5050 19112 5098
rect 19046 4998 19056 5050
rect 19108 4998 19112 5050
rect 18169 4985 18277 4992
rect 14698 4891 14756 4897
rect 14698 4857 14710 4891
rect 14744 4888 14756 4891
rect 15438 4891 15496 4897
rect 15438 4888 15450 4891
rect 14744 4860 15450 4888
rect 14744 4857 14756 4860
rect 14698 4851 14756 4857
rect 15438 4857 15450 4860
rect 15484 4857 15496 4891
rect 15438 4851 15496 4857
rect 14882 4823 14940 4829
rect 14882 4820 14894 4823
rect 14560 4792 14894 4820
rect 14560 4789 14572 4792
rect 14514 4783 14572 4789
rect 14882 4789 14894 4792
rect 14928 4820 14940 4823
rect 15254 4823 15312 4829
rect 15254 4820 15266 4823
rect 14928 4792 15266 4820
rect 14928 4789 14940 4792
rect 14882 4783 14940 4789
rect 15254 4789 15266 4792
rect 15300 4820 15312 4823
rect 15530 4823 15588 4829
rect 15530 4820 15542 4823
rect 15300 4792 15542 4820
rect 15300 4789 15312 4792
rect 15254 4783 15312 4789
rect 15530 4789 15542 4792
rect 15576 4789 15588 4823
rect 15530 4783 15588 4789
rect 16536 4805 16594 4811
rect 11166 4765 11224 4771
rect 16536 4771 16548 4805
rect 16582 4802 16594 4805
rect 16622 4802 16650 4978
rect 16720 4873 16778 4879
rect 16720 4839 16732 4873
rect 16766 4870 16778 4873
rect 17460 4873 17518 4879
rect 17460 4870 17472 4873
rect 16766 4842 17472 4870
rect 16766 4839 16778 4842
rect 16720 4833 16778 4839
rect 17460 4839 17472 4842
rect 17506 4839 17518 4873
rect 17460 4833 17518 4839
rect 16904 4805 16962 4811
rect 16904 4802 16916 4805
rect 16582 4774 16916 4802
rect 16582 4771 16594 4774
rect 12604 4761 12662 4767
rect 11440 4732 11500 4756
rect 11440 4696 11454 4732
rect 11494 4730 11500 4732
rect 11494 4712 11818 4730
rect 12604 4727 12616 4761
rect 12650 4758 12662 4761
rect 13064 4761 13122 4767
rect 13064 4758 13076 4761
rect 12650 4730 13076 4758
rect 12650 4727 12662 4730
rect 12604 4721 12662 4727
rect 13064 4727 13076 4730
rect 13110 4758 13122 4761
rect 13436 4761 13494 4767
rect 16536 4765 16594 4771
rect 16904 4771 16916 4774
rect 16950 4802 16962 4805
rect 17276 4805 17334 4811
rect 17276 4802 17288 4805
rect 16950 4774 17288 4802
rect 16950 4771 16962 4774
rect 16904 4765 16962 4771
rect 17276 4771 17288 4774
rect 17322 4802 17334 4805
rect 17552 4805 17610 4811
rect 17552 4802 17564 4805
rect 17322 4774 17564 4802
rect 17322 4771 17334 4774
rect 17276 4765 17334 4771
rect 17552 4771 17564 4774
rect 17598 4771 17610 4805
rect 17552 4765 17610 4771
rect 13436 4758 13448 4761
rect 13110 4730 13448 4758
rect 13110 4727 13122 4730
rect 13064 4721 13122 4727
rect 11494 4696 12102 4712
rect 11440 4692 12102 4696
rect 11440 4680 11500 4692
rect 11774 4690 12102 4692
rect 12700 4694 12760 4700
rect 12700 4690 12714 4694
rect 11774 4660 12714 4690
rect 12748 4660 12760 4694
rect 11774 4652 12760 4660
rect 12700 4638 12760 4652
rect 10046 4590 11518 4598
rect 10046 4580 11612 4590
rect 10046 4567 10788 4580
rect 10844 4567 11612 4580
rect 10046 4533 10075 4567
rect 10109 4533 10167 4567
rect 10201 4533 10259 4567
rect 10293 4533 10351 4567
rect 10385 4566 10443 4567
rect 10477 4566 10535 4567
rect 10385 4533 10440 4566
rect 10492 4533 10535 4566
rect 10569 4533 10627 4567
rect 10661 4533 10719 4567
rect 10753 4533 10788 4567
rect 10845 4533 10903 4567
rect 10937 4533 10995 4567
rect 11029 4533 11087 4567
rect 11121 4533 11179 4567
rect 11213 4533 11271 4567
rect 11305 4533 11363 4567
rect 11397 4533 11455 4567
rect 11489 4533 11612 4567
rect 13158 4554 13186 4730
rect 13436 4727 13448 4730
rect 13482 4727 13494 4761
rect 13436 4721 13494 4727
rect 14606 4755 14664 4761
rect 14606 4721 14618 4755
rect 14652 4752 14664 4755
rect 15066 4755 15124 4761
rect 15066 4752 15078 4755
rect 14652 4724 15078 4752
rect 14652 4721 14664 4724
rect 14606 4715 14664 4721
rect 15066 4721 15078 4724
rect 15112 4752 15124 4755
rect 15438 4755 15496 4761
rect 15438 4752 15450 4755
rect 15112 4724 15450 4752
rect 15112 4721 15124 4724
rect 15066 4715 15124 4721
rect 13718 4688 13770 4706
rect 14702 4688 14762 4694
rect 13716 4652 13730 4688
rect 13764 4684 14105 4688
rect 14702 4684 14716 4688
rect 13764 4654 14716 4684
rect 14750 4654 14762 4688
rect 13764 4652 14762 4654
rect 13716 4650 14762 4652
rect 13718 4640 13770 4650
rect 14082 4646 14762 4650
rect 14702 4632 14762 4646
rect 12316 4546 13788 4554
rect 15160 4548 15188 4724
rect 15438 4721 15450 4724
rect 15484 4721 15496 4755
rect 15438 4715 15496 4721
rect 16628 4737 16686 4743
rect 16628 4703 16640 4737
rect 16674 4734 16686 4737
rect 17088 4737 17146 4743
rect 17088 4734 17100 4737
rect 16674 4706 17100 4734
rect 16674 4703 16686 4706
rect 15720 4682 15772 4700
rect 16628 4697 16686 4703
rect 17088 4703 17100 4706
rect 17134 4734 17146 4737
rect 17460 4737 17518 4743
rect 17460 4734 17472 4737
rect 17134 4706 17472 4734
rect 17134 4703 17146 4706
rect 17088 4697 17146 4703
rect 15718 4646 15732 4682
rect 15766 4666 15870 4682
rect 16724 4670 16784 4676
rect 16724 4666 16738 4670
rect 15766 4646 16738 4666
rect 15718 4644 16738 4646
rect 15720 4634 15772 4644
rect 15845 4636 16738 4644
rect 16772 4636 16784 4670
rect 15845 4628 16784 4636
rect 16724 4614 16784 4628
rect 10046 4512 10440 4533
rect 10492 4522 10788 4533
rect 10844 4524 11612 4533
rect 12228 4534 13788 4546
rect 14318 4534 15790 4548
rect 10844 4522 11518 4524
rect 10492 4512 11518 4522
rect 10046 4502 11518 4512
rect 12228 4523 13036 4534
rect 13092 4523 13788 4534
rect 12228 4489 12345 4523
rect 12379 4489 12437 4523
rect 12471 4489 12529 4523
rect 12563 4489 12621 4523
rect 12655 4489 12713 4523
rect 12747 4489 12805 4523
rect 12839 4489 12897 4523
rect 12931 4489 12989 4523
rect 13023 4489 13036 4523
rect 13115 4489 13173 4523
rect 13207 4489 13265 4523
rect 13299 4489 13357 4523
rect 13391 4489 13449 4523
rect 13483 4489 13541 4523
rect 13575 4489 13633 4523
rect 13667 4489 13725 4523
rect 13759 4489 13788 4523
rect 12228 4480 13036 4489
rect 12316 4476 13036 4480
rect 13092 4476 13788 4489
rect 12316 4458 13788 4476
rect 14228 4528 15790 4534
rect 17182 4530 17210 4706
rect 17460 4703 17472 4706
rect 17506 4703 17518 4737
rect 17460 4697 17518 4703
rect 17742 4664 17794 4682
rect 18169 4664 18207 4985
rect 19046 4944 19112 4998
rect 19106 4828 19226 4894
rect 17740 4628 17754 4664
rect 17788 4628 18207 4664
rect 17740 4626 18207 4628
rect 17742 4616 17794 4626
rect 14228 4517 15038 4528
rect 15094 4517 15790 4528
rect 14228 4483 14347 4517
rect 14381 4483 14439 4517
rect 14473 4483 14531 4517
rect 14565 4483 14623 4517
rect 14657 4483 14715 4517
rect 14749 4483 14807 4517
rect 14841 4483 14899 4517
rect 14933 4483 14991 4517
rect 15025 4483 15038 4517
rect 15117 4483 15175 4517
rect 15209 4483 15267 4517
rect 15301 4483 15359 4517
rect 15393 4483 15451 4517
rect 15485 4483 15543 4517
rect 15577 4483 15635 4517
rect 15669 4483 15727 4517
rect 15761 4483 15790 4517
rect 16340 4510 17812 4530
rect 14228 4470 15038 4483
rect 15094 4470 15790 4483
rect 14228 4468 15790 4470
rect 14318 4452 15790 4468
rect 16254 4499 17060 4510
rect 17116 4499 17812 4510
rect 16254 4465 16369 4499
rect 16403 4465 16461 4499
rect 16495 4465 16553 4499
rect 16587 4465 16645 4499
rect 16679 4465 16737 4499
rect 16771 4465 16829 4499
rect 16863 4465 16921 4499
rect 16955 4465 17013 4499
rect 17047 4465 17060 4499
rect 17139 4465 17197 4499
rect 17231 4465 17289 4499
rect 17323 4465 17381 4499
rect 17415 4465 17473 4499
rect 17507 4465 17565 4499
rect 17599 4465 17657 4499
rect 17691 4465 17749 4499
rect 17783 4465 17812 4499
rect 16254 4452 17060 4465
rect 17116 4452 17812 4465
rect 16254 4444 17812 4452
rect 16340 4434 17812 4444
rect 6037 3357 6133 3388
rect 6104 3130 6198 3138
rect 6104 3078 6138 3130
rect 6190 3078 6198 3130
rect 6232 3136 6298 3138
rect 6232 3084 6238 3136
rect 6290 3084 6298 3136
rect 6232 3078 6298 3084
rect 6104 3072 6198 3078
rect 6006 2756 6128 2822
rect 7733 2338 7899 2340
rect 9700 2338 9883 2340
rect 11684 2338 11827 2340
rect 13613 2338 13829 2340
rect 15706 2338 15935 2340
rect 1806 2332 3278 2336
rect 1695 2318 3278 2332
rect 1695 2305 2604 2318
rect 2660 2305 3278 2318
rect 1695 2301 1835 2305
rect 1806 2271 1835 2301
rect 1869 2271 1927 2305
rect 1961 2271 2019 2305
rect 2053 2271 2111 2305
rect 2145 2271 2203 2305
rect 2237 2271 2295 2305
rect 2329 2271 2387 2305
rect 2421 2271 2479 2305
rect 2513 2271 2571 2305
rect 2660 2271 2663 2305
rect 2697 2271 2755 2305
rect 2789 2271 2847 2305
rect 2881 2271 2939 2305
rect 2973 2271 3031 2305
rect 3065 2271 3123 2305
rect 3157 2271 3215 2305
rect 3249 2271 3278 2305
rect 3788 2332 3961 2334
rect 5747 2332 5875 2334
rect 3788 2314 5348 2332
rect 3788 2303 4592 2314
rect 1806 2260 2604 2271
rect 2660 2260 3278 2271
rect 1806 2240 3278 2260
rect 3876 2301 4592 2303
rect 4648 2301 5348 2314
rect 5747 2314 7300 2332
rect 5747 2303 6544 2314
rect 3876 2267 3905 2301
rect 3939 2267 3997 2301
rect 4031 2267 4089 2301
rect 4123 2267 4181 2301
rect 4215 2267 4273 2301
rect 4307 2267 4365 2301
rect 4399 2267 4457 2301
rect 4491 2267 4549 2301
rect 4583 2267 4592 2301
rect 4675 2267 4733 2301
rect 4767 2267 4825 2301
rect 4859 2267 4917 2301
rect 4951 2267 5009 2301
rect 5043 2267 5101 2301
rect 5135 2267 5193 2301
rect 5227 2267 5285 2301
rect 5319 2267 5348 2301
rect 3876 2256 4592 2267
rect 4648 2256 5348 2267
rect 2002 2067 2060 2073
rect 2002 2033 2014 2067
rect 2048 2064 2060 2067
rect 2088 2064 2116 2240
rect 3876 2236 5348 2256
rect 5828 2301 6544 2303
rect 6600 2301 7300 2314
rect 7733 2320 9302 2338
rect 7733 2309 8546 2320
rect 5828 2267 5857 2301
rect 5891 2267 5949 2301
rect 5983 2267 6041 2301
rect 6075 2267 6133 2301
rect 6167 2267 6225 2301
rect 6259 2267 6317 2301
rect 6351 2267 6409 2301
rect 6443 2267 6501 2301
rect 6535 2267 6544 2301
rect 6627 2267 6685 2301
rect 6719 2267 6777 2301
rect 6811 2267 6869 2301
rect 6903 2267 6961 2301
rect 6995 2267 7053 2301
rect 7087 2267 7145 2301
rect 7179 2267 7237 2301
rect 7271 2267 7300 2301
rect 5828 2256 6544 2267
rect 6600 2256 7300 2267
rect 5828 2236 7300 2256
rect 7830 2307 8546 2309
rect 8602 2307 9302 2320
rect 9700 2320 11254 2338
rect 9700 2309 10498 2320
rect 7830 2273 7859 2307
rect 7893 2273 7951 2307
rect 7985 2273 8043 2307
rect 8077 2273 8135 2307
rect 8169 2273 8227 2307
rect 8261 2273 8319 2307
rect 8353 2273 8411 2307
rect 8445 2273 8503 2307
rect 8537 2273 8546 2307
rect 8629 2273 8687 2307
rect 8721 2273 8779 2307
rect 8813 2273 8871 2307
rect 8905 2273 8963 2307
rect 8997 2273 9055 2307
rect 9089 2273 9147 2307
rect 9181 2273 9239 2307
rect 9273 2273 9302 2307
rect 7830 2262 8546 2273
rect 8602 2262 9302 2273
rect 7830 2242 9302 2262
rect 9782 2307 10498 2309
rect 10554 2307 11254 2320
rect 11684 2320 13246 2338
rect 11684 2309 12490 2320
rect 9782 2273 9811 2307
rect 9845 2273 9903 2307
rect 9937 2273 9995 2307
rect 10029 2273 10087 2307
rect 10121 2273 10179 2307
rect 10213 2273 10271 2307
rect 10305 2273 10363 2307
rect 10397 2273 10455 2307
rect 10489 2273 10498 2307
rect 10581 2273 10639 2307
rect 10673 2273 10731 2307
rect 10765 2273 10823 2307
rect 10857 2273 10915 2307
rect 10949 2273 11007 2307
rect 11041 2273 11099 2307
rect 11133 2273 11191 2307
rect 11225 2273 11254 2307
rect 9782 2262 10498 2273
rect 10554 2262 11254 2273
rect 9782 2242 11254 2262
rect 11774 2307 12490 2309
rect 12546 2307 13246 2320
rect 13613 2320 15198 2338
rect 13613 2309 14442 2320
rect 11774 2273 11803 2307
rect 11837 2273 11895 2307
rect 11929 2273 11987 2307
rect 12021 2273 12079 2307
rect 12113 2273 12171 2307
rect 12205 2273 12263 2307
rect 12297 2273 12355 2307
rect 12389 2273 12447 2307
rect 12481 2273 12490 2307
rect 12573 2273 12631 2307
rect 12665 2273 12723 2307
rect 12757 2273 12815 2307
rect 12849 2273 12907 2307
rect 12941 2273 12999 2307
rect 13033 2273 13091 2307
rect 13125 2273 13183 2307
rect 13217 2273 13246 2307
rect 11774 2262 12490 2273
rect 12546 2262 13246 2273
rect 11774 2242 13246 2262
rect 13726 2307 14442 2309
rect 14498 2307 15198 2320
rect 15706 2320 17262 2338
rect 15706 2309 16506 2320
rect 13726 2273 13755 2307
rect 13789 2273 13847 2307
rect 13881 2273 13939 2307
rect 13973 2273 14031 2307
rect 14065 2273 14123 2307
rect 14157 2273 14215 2307
rect 14249 2273 14307 2307
rect 14341 2273 14399 2307
rect 14433 2273 14442 2307
rect 14525 2273 14583 2307
rect 14617 2273 14675 2307
rect 14709 2273 14767 2307
rect 14801 2273 14859 2307
rect 14893 2273 14951 2307
rect 14985 2273 15043 2307
rect 15077 2273 15135 2307
rect 15169 2273 15198 2307
rect 13726 2262 14442 2273
rect 14498 2262 15198 2273
rect 13726 2242 15198 2262
rect 15790 2307 16506 2309
rect 16562 2307 17262 2320
rect 15790 2273 15819 2307
rect 15853 2273 15911 2307
rect 15945 2273 16003 2307
rect 16037 2273 16095 2307
rect 16129 2273 16187 2307
rect 16221 2273 16279 2307
rect 16313 2273 16371 2307
rect 16405 2273 16463 2307
rect 16497 2273 16506 2307
rect 16589 2273 16647 2307
rect 16681 2273 16739 2307
rect 16773 2273 16831 2307
rect 16865 2273 16923 2307
rect 16957 2273 17015 2307
rect 17049 2273 17107 2307
rect 17141 2273 17199 2307
rect 17233 2273 17262 2307
rect 15790 2262 16506 2273
rect 16562 2262 17262 2273
rect 15790 2242 17262 2262
rect 2186 2135 2244 2141
rect 2186 2101 2198 2135
rect 2232 2132 2244 2135
rect 2926 2135 2984 2141
rect 2926 2132 2938 2135
rect 2232 2104 2938 2132
rect 2232 2101 2244 2104
rect 2186 2095 2244 2101
rect 2926 2101 2938 2104
rect 2972 2101 2984 2135
rect 2926 2095 2984 2101
rect 2370 2067 2428 2073
rect 2370 2064 2382 2067
rect 2048 2036 2382 2064
rect 2048 2033 2060 2036
rect 2002 2027 2060 2033
rect 2370 2033 2382 2036
rect 2416 2064 2428 2067
rect 2742 2067 2800 2073
rect 2742 2064 2754 2067
rect 2416 2036 2754 2064
rect 2416 2033 2428 2036
rect 2370 2027 2428 2033
rect 2742 2033 2754 2036
rect 2788 2064 2800 2067
rect 3018 2067 3076 2073
rect 3018 2064 3030 2067
rect 2788 2036 3030 2064
rect 2788 2033 2800 2036
rect 2742 2027 2800 2033
rect 3018 2033 3030 2036
rect 3064 2033 3076 2067
rect 3018 2027 3076 2033
rect 4072 2063 4130 2069
rect 4072 2029 4084 2063
rect 4118 2060 4130 2063
rect 4158 2060 4186 2236
rect 4256 2131 4314 2137
rect 4256 2097 4268 2131
rect 4302 2128 4314 2131
rect 4996 2131 5054 2137
rect 4996 2128 5008 2131
rect 4302 2100 5008 2128
rect 4302 2097 4314 2100
rect 4256 2091 4314 2097
rect 4996 2097 5008 2100
rect 5042 2097 5054 2131
rect 4996 2091 5054 2097
rect 4440 2063 4498 2069
rect 4440 2060 4452 2063
rect 4118 2032 4452 2060
rect 4118 2029 4130 2032
rect 4072 2023 4130 2029
rect 4440 2029 4452 2032
rect 4486 2060 4498 2063
rect 4812 2063 4870 2069
rect 4812 2060 4824 2063
rect 4486 2032 4824 2060
rect 4486 2029 4498 2032
rect 4440 2023 4498 2029
rect 4812 2029 4824 2032
rect 4858 2060 4870 2063
rect 5088 2063 5146 2069
rect 5088 2060 5100 2063
rect 4858 2032 5100 2060
rect 4858 2029 4870 2032
rect 4812 2023 4870 2029
rect 5088 2029 5100 2032
rect 5134 2029 5146 2063
rect 5088 2023 5146 2029
rect 6024 2063 6082 2069
rect 6024 2029 6036 2063
rect 6070 2060 6082 2063
rect 6110 2060 6138 2236
rect 6208 2131 6266 2137
rect 6208 2097 6220 2131
rect 6254 2128 6266 2131
rect 6948 2131 7006 2137
rect 6948 2128 6960 2131
rect 6254 2100 6960 2128
rect 6254 2097 6266 2100
rect 6208 2091 6266 2097
rect 6948 2097 6960 2100
rect 6994 2097 7006 2131
rect 6948 2091 7006 2097
rect 8026 2069 8084 2075
rect 6392 2063 6450 2069
rect 6392 2060 6404 2063
rect 6070 2032 6404 2060
rect 6070 2029 6082 2032
rect 6024 2023 6082 2029
rect 6392 2029 6404 2032
rect 6438 2060 6450 2063
rect 6764 2063 6822 2069
rect 6764 2060 6776 2063
rect 6438 2032 6776 2060
rect 6438 2029 6450 2032
rect 6392 2023 6450 2029
rect 6764 2029 6776 2032
rect 6810 2060 6822 2063
rect 7040 2063 7098 2069
rect 7040 2060 7052 2063
rect 6810 2032 7052 2060
rect 6810 2029 6822 2032
rect 6764 2023 6822 2029
rect 7040 2029 7052 2032
rect 7086 2029 7098 2063
rect 8026 2035 8038 2069
rect 8072 2066 8084 2069
rect 8112 2066 8140 2242
rect 8210 2137 8268 2143
rect 8210 2103 8222 2137
rect 8256 2134 8268 2137
rect 8950 2137 9008 2143
rect 8950 2134 8962 2137
rect 8256 2106 8962 2134
rect 8256 2103 8268 2106
rect 8210 2097 8268 2103
rect 8950 2103 8962 2106
rect 8996 2103 9008 2137
rect 8950 2097 9008 2103
rect 8394 2069 8452 2075
rect 8394 2066 8406 2069
rect 8072 2038 8406 2066
rect 8072 2035 8084 2038
rect 8026 2029 8084 2035
rect 8394 2035 8406 2038
rect 8440 2066 8452 2069
rect 8766 2069 8824 2075
rect 8766 2066 8778 2069
rect 8440 2038 8778 2066
rect 8440 2035 8452 2038
rect 8394 2029 8452 2035
rect 8766 2035 8778 2038
rect 8812 2066 8824 2069
rect 9042 2069 9100 2075
rect 9042 2066 9054 2069
rect 8812 2038 9054 2066
rect 8812 2035 8824 2038
rect 8766 2029 8824 2035
rect 9042 2035 9054 2038
rect 9088 2035 9100 2069
rect 9042 2029 9100 2035
rect 9978 2069 10036 2075
rect 9978 2035 9990 2069
rect 10024 2066 10036 2069
rect 10064 2066 10092 2242
rect 10162 2137 10220 2143
rect 10162 2103 10174 2137
rect 10208 2134 10220 2137
rect 10902 2137 10960 2143
rect 10902 2134 10914 2137
rect 10208 2106 10914 2134
rect 10208 2103 10220 2106
rect 10162 2097 10220 2103
rect 10902 2103 10914 2106
rect 10948 2103 10960 2137
rect 10902 2097 10960 2103
rect 10346 2069 10404 2075
rect 10346 2066 10358 2069
rect 10024 2038 10358 2066
rect 10024 2035 10036 2038
rect 9978 2029 10036 2035
rect 10346 2035 10358 2038
rect 10392 2066 10404 2069
rect 10718 2069 10776 2075
rect 10718 2066 10730 2069
rect 10392 2038 10730 2066
rect 10392 2035 10404 2038
rect 10346 2029 10404 2035
rect 10718 2035 10730 2038
rect 10764 2066 10776 2069
rect 10994 2069 11052 2075
rect 10994 2066 11006 2069
rect 10764 2038 11006 2066
rect 10764 2035 10776 2038
rect 10718 2029 10776 2035
rect 10994 2035 11006 2038
rect 11040 2035 11052 2069
rect 10994 2029 11052 2035
rect 11970 2069 12028 2075
rect 11970 2035 11982 2069
rect 12016 2066 12028 2069
rect 12056 2066 12084 2242
rect 12154 2137 12212 2143
rect 12154 2103 12166 2137
rect 12200 2134 12212 2137
rect 12894 2137 12952 2143
rect 12894 2134 12906 2137
rect 12200 2106 12906 2134
rect 12200 2103 12212 2106
rect 12154 2097 12212 2103
rect 12894 2103 12906 2106
rect 12940 2103 12952 2137
rect 12894 2097 12952 2103
rect 12338 2069 12396 2075
rect 12338 2066 12350 2069
rect 12016 2038 12350 2066
rect 12016 2035 12028 2038
rect 11970 2029 12028 2035
rect 12338 2035 12350 2038
rect 12384 2066 12396 2069
rect 12710 2069 12768 2075
rect 12710 2066 12722 2069
rect 12384 2038 12722 2066
rect 12384 2035 12396 2038
rect 12338 2029 12396 2035
rect 12710 2035 12722 2038
rect 12756 2066 12768 2069
rect 12986 2069 13044 2075
rect 12986 2066 12998 2069
rect 12756 2038 12998 2066
rect 12756 2035 12768 2038
rect 12710 2029 12768 2035
rect 12986 2035 12998 2038
rect 13032 2035 13044 2069
rect 12986 2029 13044 2035
rect 13922 2069 13980 2075
rect 13922 2035 13934 2069
rect 13968 2066 13980 2069
rect 14008 2066 14036 2242
rect 14106 2137 14164 2143
rect 14106 2103 14118 2137
rect 14152 2134 14164 2137
rect 14846 2137 14904 2143
rect 14846 2134 14858 2137
rect 14152 2106 14858 2134
rect 14152 2103 14164 2106
rect 14106 2097 14164 2103
rect 14846 2103 14858 2106
rect 14892 2103 14904 2137
rect 14846 2097 14904 2103
rect 14290 2069 14348 2075
rect 14290 2066 14302 2069
rect 13968 2038 14302 2066
rect 13968 2035 13980 2038
rect 13922 2029 13980 2035
rect 14290 2035 14302 2038
rect 14336 2066 14348 2069
rect 14662 2069 14720 2075
rect 14662 2066 14674 2069
rect 14336 2038 14674 2066
rect 14336 2035 14348 2038
rect 14290 2029 14348 2035
rect 14662 2035 14674 2038
rect 14708 2066 14720 2069
rect 14938 2069 14996 2075
rect 14938 2066 14950 2069
rect 14708 2038 14950 2066
rect 14708 2035 14720 2038
rect 14662 2029 14720 2035
rect 14938 2035 14950 2038
rect 14984 2035 14996 2069
rect 14938 2029 14996 2035
rect 15986 2069 16044 2075
rect 15986 2035 15998 2069
rect 16032 2066 16044 2069
rect 16072 2066 16100 2242
rect 16170 2137 16228 2143
rect 16170 2103 16182 2137
rect 16216 2134 16228 2137
rect 16910 2137 16968 2143
rect 16910 2134 16922 2137
rect 16216 2106 16922 2134
rect 16216 2103 16228 2106
rect 16170 2097 16228 2103
rect 16910 2103 16922 2106
rect 16956 2103 16968 2137
rect 16910 2097 16968 2103
rect 16354 2069 16412 2075
rect 16354 2066 16366 2069
rect 16032 2038 16366 2066
rect 16032 2035 16044 2038
rect 15986 2029 16044 2035
rect 16354 2035 16366 2038
rect 16400 2066 16412 2069
rect 16726 2069 16784 2075
rect 16726 2066 16738 2069
rect 16400 2038 16738 2066
rect 16400 2035 16412 2038
rect 16354 2029 16412 2035
rect 16726 2035 16738 2038
rect 16772 2066 16784 2069
rect 17002 2069 17060 2075
rect 17002 2066 17014 2069
rect 16772 2038 17014 2066
rect 16772 2035 16784 2038
rect 16726 2029 16784 2035
rect 17002 2035 17014 2038
rect 17048 2035 17060 2069
rect 17002 2029 17060 2035
rect 7040 2023 7098 2029
rect 2094 1999 2152 2005
rect 2094 1965 2106 1999
rect 2140 1996 2152 1999
rect 2554 1999 2612 2005
rect 2554 1996 2566 1999
rect 2140 1968 2566 1996
rect 2140 1965 2152 1968
rect 2094 1959 2152 1965
rect 2554 1965 2566 1968
rect 2600 1996 2612 1999
rect 2926 1999 2984 2005
rect 8118 2001 8176 2007
rect 2926 1996 2938 1999
rect 2600 1968 2938 1996
rect 2600 1965 2612 1968
rect 2554 1959 2612 1965
rect 2192 1938 2258 1940
rect 2192 1886 2198 1938
rect 2250 1886 2258 1938
rect 2192 1882 2258 1886
rect 2648 1792 2676 1968
rect 2926 1965 2938 1968
rect 2972 1965 2984 1999
rect 2926 1959 2984 1965
rect 4164 1995 4222 2001
rect 4164 1961 4176 1995
rect 4210 1992 4222 1995
rect 4624 1995 4682 2001
rect 4624 1992 4636 1995
rect 4210 1964 4636 1992
rect 4210 1961 4222 1964
rect 4164 1955 4222 1961
rect 4624 1961 4636 1964
rect 4670 1992 4682 1995
rect 4996 1995 5054 2001
rect 4996 1992 5008 1995
rect 4670 1964 5008 1992
rect 4670 1961 4682 1964
rect 4624 1955 4682 1961
rect 3200 1926 3260 1950
rect 3200 1890 3214 1926
rect 3254 1924 3260 1926
rect 4260 1928 4320 1934
rect 4260 1924 4274 1928
rect 3254 1894 4274 1924
rect 4308 1894 4320 1928
rect 3254 1890 4320 1894
rect 3200 1886 4320 1890
rect 3200 1874 3260 1886
rect 4260 1872 4320 1886
rect 1806 1778 3278 1792
rect 4718 1788 4746 1964
rect 4996 1961 5008 1964
rect 5042 1961 5054 1995
rect 4996 1955 5054 1961
rect 6116 1995 6174 2001
rect 6116 1961 6128 1995
rect 6162 1992 6174 1995
rect 6576 1995 6634 2001
rect 6576 1992 6588 1995
rect 6162 1964 6588 1992
rect 6162 1961 6174 1964
rect 6116 1955 6174 1961
rect 6576 1961 6588 1964
rect 6622 1992 6634 1995
rect 6948 1995 7006 2001
rect 6948 1992 6960 1995
rect 6622 1964 6960 1992
rect 6622 1961 6634 1964
rect 6576 1955 6634 1961
rect 5278 1922 5330 1940
rect 6212 1928 6272 1934
rect 6212 1924 6226 1928
rect 5518 1922 6226 1924
rect 5276 1886 5290 1922
rect 5324 1894 6226 1922
rect 6260 1894 6272 1928
rect 5324 1886 6272 1894
rect 5276 1884 5565 1886
rect 5278 1874 5330 1884
rect 6212 1872 6272 1886
rect 6670 1788 6698 1964
rect 6948 1961 6960 1964
rect 6994 1961 7006 1995
rect 8118 1967 8130 2001
rect 8164 1998 8176 2001
rect 8578 2001 8636 2007
rect 8578 1998 8590 2001
rect 8164 1970 8590 1998
rect 8164 1967 8176 1970
rect 8118 1961 8176 1967
rect 8578 1967 8590 1970
rect 8624 1998 8636 2001
rect 8950 2001 9008 2007
rect 8950 1998 8962 2001
rect 8624 1970 8962 1998
rect 8624 1967 8636 1970
rect 8578 1961 8636 1967
rect 6948 1955 7006 1961
rect 7230 1922 7282 1940
rect 8214 1934 8274 1940
rect 8214 1930 8228 1934
rect 7456 1922 8228 1930
rect 7228 1886 7242 1922
rect 7276 1900 8228 1922
rect 8262 1900 8274 1934
rect 7276 1892 8274 1900
rect 7276 1886 7517 1892
rect 7228 1884 7517 1886
rect 7230 1874 7282 1884
rect 8214 1878 8274 1892
rect 8672 1794 8700 1970
rect 8950 1967 8962 1970
rect 8996 1967 9008 2001
rect 8950 1961 9008 1967
rect 10070 2001 10128 2007
rect 10070 1967 10082 2001
rect 10116 1998 10128 2001
rect 10530 2001 10588 2007
rect 10530 1998 10542 2001
rect 10116 1970 10542 1998
rect 10116 1967 10128 1970
rect 10070 1961 10128 1967
rect 10530 1967 10542 1970
rect 10576 1998 10588 2001
rect 10902 2001 10960 2007
rect 10902 1998 10914 2001
rect 10576 1970 10914 1998
rect 10576 1967 10588 1970
rect 10530 1961 10588 1967
rect 9232 1928 9284 1946
rect 10166 1934 10226 1940
rect 10166 1930 10180 1934
rect 9472 1928 10180 1930
rect 9230 1892 9244 1928
rect 9278 1900 10180 1928
rect 10214 1900 10226 1934
rect 9278 1892 10226 1900
rect 9230 1890 9519 1892
rect 9232 1880 9284 1890
rect 10166 1878 10226 1892
rect 10624 1794 10652 1970
rect 10902 1967 10914 1970
rect 10948 1967 10960 2001
rect 10902 1961 10960 1967
rect 12062 2001 12120 2007
rect 12062 1967 12074 2001
rect 12108 1998 12120 2001
rect 12522 2001 12580 2007
rect 12522 1998 12534 2001
rect 12108 1970 12534 1998
rect 12108 1967 12120 1970
rect 12062 1961 12120 1967
rect 12522 1967 12534 1970
rect 12568 1998 12580 2001
rect 12894 2001 12952 2007
rect 12894 1998 12906 2001
rect 12568 1970 12906 1998
rect 12568 1967 12580 1970
rect 12522 1961 12580 1967
rect 11184 1928 11236 1946
rect 12158 1934 12218 1940
rect 12158 1930 12172 1934
rect 11317 1928 12172 1930
rect 11182 1892 11196 1928
rect 11230 1900 12172 1928
rect 12206 1900 12218 1934
rect 11230 1892 12218 1900
rect 11182 1890 11382 1892
rect 11184 1880 11236 1890
rect 12158 1878 12218 1892
rect 12616 1794 12644 1970
rect 12894 1967 12906 1970
rect 12940 1967 12952 2001
rect 12894 1961 12952 1967
rect 14014 2001 14072 2007
rect 14014 1967 14026 2001
rect 14060 1998 14072 2001
rect 14474 2001 14532 2007
rect 14474 1998 14486 2001
rect 14060 1970 14486 1998
rect 14060 1967 14072 1970
rect 14014 1961 14072 1967
rect 14474 1967 14486 1970
rect 14520 1998 14532 2001
rect 14846 2001 14904 2007
rect 14846 1998 14858 2001
rect 14520 1970 14858 1998
rect 14520 1967 14532 1970
rect 14474 1961 14532 1967
rect 13176 1928 13228 1946
rect 14110 1934 14170 1940
rect 14110 1930 14124 1934
rect 13416 1928 14124 1930
rect 13174 1892 13188 1928
rect 13222 1900 14124 1928
rect 14158 1900 14170 1934
rect 13222 1892 14170 1900
rect 13174 1890 13463 1892
rect 13176 1880 13228 1890
rect 14110 1878 14170 1892
rect 14568 1794 14596 1970
rect 14846 1967 14858 1970
rect 14892 1967 14904 2001
rect 14846 1961 14904 1967
rect 16078 2001 16136 2007
rect 16078 1967 16090 2001
rect 16124 1998 16136 2001
rect 16538 2001 16596 2007
rect 16538 1998 16550 2001
rect 16124 1970 16550 1998
rect 16124 1967 16136 1970
rect 16078 1961 16136 1967
rect 16538 1967 16550 1970
rect 16584 1998 16596 2001
rect 16910 2001 16968 2007
rect 16910 1998 16922 2001
rect 16584 1970 16922 1998
rect 16584 1967 16596 1970
rect 16538 1961 16596 1967
rect 15128 1928 15180 1946
rect 16174 1934 16234 1940
rect 16174 1930 16188 1934
rect 15538 1928 16188 1930
rect 15126 1892 15140 1928
rect 15174 1900 16188 1928
rect 16222 1900 16234 1934
rect 15174 1892 16234 1900
rect 15126 1890 15575 1892
rect 15128 1880 15180 1890
rect 16174 1878 16234 1892
rect 16632 1794 16660 1970
rect 16910 1967 16922 1970
rect 16956 1967 16968 2001
rect 16910 1961 16968 1967
rect 17192 1928 17244 1946
rect 17362 1930 17488 1982
rect 17362 1928 17402 1930
rect 17190 1892 17204 1928
rect 17238 1892 17402 1928
rect 17190 1890 17402 1892
rect 17192 1880 17244 1890
rect 17362 1876 17402 1890
rect 17454 1876 17488 1930
rect 17362 1828 17488 1876
rect 1806 1761 2604 1778
rect 2656 1761 3278 1778
rect 1806 1727 1835 1761
rect 1869 1727 1927 1761
rect 1961 1727 2019 1761
rect 2053 1727 2111 1761
rect 2145 1727 2203 1761
rect 2237 1727 2295 1761
rect 2329 1727 2387 1761
rect 2421 1727 2479 1761
rect 2513 1727 2571 1761
rect 2656 1727 2663 1761
rect 2697 1727 2755 1761
rect 2789 1727 2847 1761
rect 2881 1727 2939 1761
rect 2973 1727 3031 1761
rect 3065 1727 3123 1761
rect 3157 1727 3215 1761
rect 3249 1727 3278 1761
rect 1806 1723 2604 1727
rect 1719 1720 2604 1723
rect 2656 1720 3278 1727
rect 3876 1768 5348 1788
rect 3876 1757 4596 1768
rect 4652 1757 5348 1768
rect 3876 1725 3905 1757
rect 1719 1696 3278 1720
rect 3783 1723 3905 1725
rect 3939 1723 3997 1757
rect 4031 1723 4089 1757
rect 4123 1723 4181 1757
rect 4215 1723 4273 1757
rect 4307 1723 4365 1757
rect 4399 1723 4457 1757
rect 4491 1723 4549 1757
rect 4583 1723 4596 1757
rect 4675 1723 4733 1757
rect 4767 1723 4825 1757
rect 4859 1723 4917 1757
rect 4951 1723 5009 1757
rect 5043 1723 5101 1757
rect 5135 1723 5193 1757
rect 5227 1723 5285 1757
rect 5319 1723 5348 1757
rect 5828 1768 7300 1788
rect 5828 1757 6548 1768
rect 6604 1757 7300 1768
rect 5828 1725 5857 1757
rect 3783 1710 4596 1723
rect 4652 1710 5348 1723
rect 1719 1692 1849 1696
rect 3783 1694 5348 1710
rect 5738 1723 5857 1725
rect 5891 1723 5949 1757
rect 5983 1723 6041 1757
rect 6075 1723 6133 1757
rect 6167 1723 6225 1757
rect 6259 1723 6317 1757
rect 6351 1723 6409 1757
rect 6443 1723 6501 1757
rect 6535 1723 6548 1757
rect 6627 1723 6685 1757
rect 6719 1723 6777 1757
rect 6811 1723 6869 1757
rect 6903 1723 6961 1757
rect 6995 1723 7053 1757
rect 7087 1723 7145 1757
rect 7179 1723 7237 1757
rect 7271 1723 7300 1757
rect 7830 1774 9302 1794
rect 7830 1763 8550 1774
rect 8606 1763 9302 1774
rect 7830 1731 7859 1763
rect 5738 1710 6548 1723
rect 6604 1710 7300 1723
rect 5738 1694 7300 1710
rect 7749 1729 7859 1731
rect 7893 1729 7951 1763
rect 7985 1729 8043 1763
rect 8077 1729 8135 1763
rect 8169 1729 8227 1763
rect 8261 1729 8319 1763
rect 8353 1729 8411 1763
rect 8445 1729 8503 1763
rect 8537 1729 8550 1763
rect 8629 1729 8687 1763
rect 8721 1729 8779 1763
rect 8813 1729 8871 1763
rect 8905 1729 8963 1763
rect 8997 1729 9055 1763
rect 9089 1729 9147 1763
rect 9181 1729 9239 1763
rect 9273 1729 9302 1763
rect 9782 1774 11254 1794
rect 9782 1763 10502 1774
rect 10558 1763 11254 1774
rect 9782 1729 9811 1763
rect 9845 1729 9903 1763
rect 9937 1729 9995 1763
rect 10029 1729 10087 1763
rect 10121 1729 10179 1763
rect 10213 1729 10271 1763
rect 10305 1729 10363 1763
rect 10397 1729 10455 1763
rect 10489 1729 10502 1763
rect 10581 1729 10639 1763
rect 10673 1729 10731 1763
rect 10765 1729 10823 1763
rect 10857 1729 10915 1763
rect 10949 1729 11007 1763
rect 11041 1729 11099 1763
rect 11133 1729 11191 1763
rect 11225 1729 11254 1763
rect 11774 1774 13246 1794
rect 11774 1763 12494 1774
rect 12550 1763 13246 1774
rect 11774 1731 11803 1763
rect 7749 1716 8550 1729
rect 8606 1716 9302 1729
rect 7749 1700 9302 1716
rect 7830 1698 9302 1700
rect 9697 1716 10502 1729
rect 10558 1716 11254 1729
rect 9697 1698 11254 1716
rect 11692 1729 11803 1731
rect 11837 1729 11895 1763
rect 11929 1729 11987 1763
rect 12021 1729 12079 1763
rect 12113 1729 12171 1763
rect 12205 1729 12263 1763
rect 12297 1729 12355 1763
rect 12389 1729 12447 1763
rect 12481 1729 12494 1763
rect 12573 1729 12631 1763
rect 12665 1729 12723 1763
rect 12757 1729 12815 1763
rect 12849 1729 12907 1763
rect 12941 1729 12999 1763
rect 13033 1729 13091 1763
rect 13125 1729 13183 1763
rect 13217 1729 13246 1763
rect 13726 1774 15198 1794
rect 13726 1763 14446 1774
rect 14502 1763 15198 1774
rect 13726 1731 13755 1763
rect 11692 1716 12494 1729
rect 12550 1716 13246 1729
rect 11692 1700 13246 1716
rect 13645 1729 13755 1731
rect 13789 1729 13847 1763
rect 13881 1729 13939 1763
rect 13973 1729 14031 1763
rect 14065 1729 14123 1763
rect 14157 1729 14215 1763
rect 14249 1729 14307 1763
rect 14341 1729 14399 1763
rect 14433 1729 14446 1763
rect 14525 1729 14583 1763
rect 14617 1729 14675 1763
rect 14709 1729 14767 1763
rect 14801 1729 14859 1763
rect 14893 1729 14951 1763
rect 14985 1729 15043 1763
rect 15077 1729 15135 1763
rect 15169 1729 15198 1763
rect 15790 1774 17262 1794
rect 15790 1763 16510 1774
rect 16566 1763 17262 1774
rect 15790 1731 15819 1763
rect 13645 1716 14446 1729
rect 14502 1716 15198 1729
rect 13645 1700 15198 1716
rect 15681 1729 15819 1731
rect 15853 1729 15911 1763
rect 15945 1729 16003 1763
rect 16037 1729 16095 1763
rect 16129 1729 16187 1763
rect 16221 1729 16279 1763
rect 16313 1729 16371 1763
rect 16405 1729 16463 1763
rect 16497 1729 16510 1763
rect 16589 1729 16647 1763
rect 16681 1729 16739 1763
rect 16773 1729 16831 1763
rect 16865 1729 16923 1763
rect 16957 1729 17015 1763
rect 17049 1729 17107 1763
rect 17141 1729 17199 1763
rect 17233 1729 17262 1763
rect 15681 1716 16510 1729
rect 16566 1716 17262 1729
rect 15681 1700 17262 1716
rect 11774 1698 13246 1700
rect 13726 1698 15198 1700
rect 15790 1698 17262 1700
rect 3876 1692 5348 1694
rect 5828 1692 7300 1694
<< via1 >>
rect 18768 43898 18962 44096
rect 18562 42762 18624 42820
rect 19124 42724 19186 42782
rect 18540 40890 18602 40948
rect 19106 40882 19168 40940
rect 18564 39262 18626 39320
rect 19106 39258 19168 39316
rect 18572 38066 18634 38124
rect 19122 38082 19184 38140
rect 18580 36996 18642 37054
rect 19128 36986 19190 37044
rect 18598 36200 18652 36256
rect 19142 36228 19200 36284
rect 18424 34427 18449 34454
rect 18449 34427 18483 34454
rect 18483 34427 18504 34454
rect 18424 34372 18504 34427
rect 18972 34427 18993 34458
rect 18993 34427 19027 34458
rect 19027 34427 19052 34458
rect 18972 34376 19052 34427
rect 18432 32121 18457 32148
rect 18457 32121 18491 32148
rect 18491 32121 18512 32148
rect 18432 32066 18512 32121
rect 18980 32121 19001 32152
rect 19001 32121 19035 32152
rect 19035 32121 19060 32152
rect 18980 32070 19060 32121
rect 18440 29907 18465 29934
rect 18465 29907 18499 29934
rect 18499 29907 18520 29934
rect 18440 29852 18520 29907
rect 18988 29907 19009 29938
rect 19009 29907 19043 29938
rect 19043 29907 19068 29938
rect 18988 29856 19068 29907
rect 18422 27707 18447 27734
rect 18447 27707 18481 27734
rect 18481 27707 18502 27734
rect 18422 27652 18502 27707
rect 18970 27707 18991 27738
rect 18991 27707 19025 27738
rect 19025 27707 19050 27738
rect 18970 27656 19050 27707
rect 18430 25493 18455 25520
rect 18455 25493 18489 25520
rect 18489 25493 18510 25520
rect 18430 25438 18510 25493
rect 18978 25493 18999 25524
rect 18999 25493 19033 25524
rect 19033 25493 19058 25524
rect 18978 25442 19058 25493
rect 8532 23405 8614 23430
rect 8532 23371 8587 23405
rect 8587 23371 8614 23405
rect 8532 23350 8614 23371
rect 10746 23413 10828 23438
rect 10746 23379 10801 23413
rect 10801 23379 10828 23413
rect 10746 23358 10828 23379
rect 12946 23395 13028 23420
rect 12946 23361 13001 23395
rect 13001 23361 13028 23395
rect 12946 23340 13028 23361
rect 15160 23403 15242 23428
rect 15160 23369 15215 23403
rect 15215 23369 15242 23403
rect 15160 23348 15242 23369
rect 17466 23411 17548 23436
rect 17466 23377 17521 23411
rect 17521 23377 17548 23411
rect 17466 23356 17548 23377
rect 8536 22861 8618 22882
rect 8536 22827 8587 22861
rect 8587 22827 8618 22861
rect 8536 22802 8618 22827
rect 10750 22869 10832 22890
rect 10750 22835 10801 22869
rect 10801 22835 10832 22869
rect 10750 22810 10832 22835
rect 12950 22851 13032 22872
rect 12950 22817 13001 22851
rect 13001 22817 13032 22851
rect 12950 22792 13032 22817
rect 15164 22859 15246 22880
rect 15164 22825 15215 22859
rect 15215 22825 15246 22859
rect 15164 22800 15246 22825
rect 17470 22867 17552 22888
rect 17470 22833 17521 22867
rect 17521 22833 17552 22867
rect 17470 22808 17552 22833
rect 9540 17762 9600 17822
rect 16455 17701 16523 17714
rect 15683 17663 15751 17674
rect 15683 17629 15688 17663
rect 15688 17629 15722 17663
rect 15722 17629 15751 17663
rect 16455 17667 16466 17701
rect 16466 17667 16500 17701
rect 16500 17667 16523 17701
rect 16455 17652 16523 17667
rect 17335 17703 17403 17714
rect 17335 17669 17340 17703
rect 17340 17669 17374 17703
rect 17374 17669 17403 17703
rect 17335 17652 17403 17669
rect 18121 17693 18189 17704
rect 18121 17659 18142 17693
rect 18142 17659 18189 17693
rect 18121 17642 18189 17659
rect 19219 17695 19287 17708
rect 19219 17661 19230 17695
rect 19230 17661 19264 17695
rect 19264 17661 19287 17695
rect 19219 17646 19287 17661
rect 15683 17612 15751 17629
rect 20099 17697 20167 17708
rect 20099 17663 20104 17697
rect 20104 17663 20138 17697
rect 20138 17663 20167 17697
rect 20099 17646 20167 17663
rect 20885 17687 20953 17698
rect 20885 17653 20906 17687
rect 20906 17653 20953 17687
rect 20885 17636 20953 17653
rect 21475 17685 21543 17698
rect 21475 17651 21486 17685
rect 21486 17651 21520 17685
rect 21520 17651 21543 17685
rect 21475 17636 21543 17651
rect 22355 17687 22423 17698
rect 22355 17653 22360 17687
rect 22360 17653 22394 17687
rect 22394 17653 22423 17687
rect 22355 17636 22423 17653
rect 23141 17677 23209 17688
rect 23141 17643 23162 17677
rect 23162 17643 23209 17677
rect 23141 17626 23209 17643
rect 6646 17504 6722 17576
rect 9536 17218 9594 17278
rect 11414 16986 11474 17042
rect 4590 16570 4642 16624
rect 4976 16020 5034 16074
rect 4746 15814 4808 15874
rect 6712 15706 6780 15768
rect 6608 15356 6660 15408
rect 4898 15270 4966 15332
rect 6130 15202 6198 15264
rect 7114 15156 7182 15218
rect 4582 14986 4648 15052
rect 5794 14654 5862 14716
rect 5012 14442 5078 14508
rect 4682 14244 4754 14314
rect 6350 14232 6418 14294
rect 7916 14222 7984 14284
rect 9456 16607 9508 16628
rect 9456 16574 9489 16607
rect 9489 16574 9508 16607
rect 10872 16344 10942 16410
rect 9842 16063 9900 16078
rect 9842 16029 9857 16063
rect 9857 16029 9900 16063
rect 9842 16024 9900 16029
rect 9612 15863 9674 15878
rect 9612 15829 9645 15863
rect 9645 15829 9674 15863
rect 9612 15818 9674 15829
rect 11578 15753 11646 15772
rect 11578 15719 11595 15753
rect 11595 15719 11629 15753
rect 11629 15719 11646 15753
rect 11578 15710 11646 15719
rect 9842 15494 9896 15506
rect 9842 15460 9872 15494
rect 9872 15460 9896 15494
rect 9842 15452 9896 15460
rect 9764 15319 9832 15336
rect 9764 15285 9771 15319
rect 9771 15285 9829 15319
rect 9829 15285 9832 15319
rect 9764 15274 9832 15285
rect 9448 15043 9514 15056
rect 9448 15009 9465 15043
rect 9465 15009 9499 15043
rect 9499 15009 9514 15043
rect 9448 14990 9514 15009
rect 11474 15404 11526 15412
rect 11474 15368 11498 15404
rect 11498 15368 11526 15404
rect 11474 15360 11526 15368
rect 10996 15253 11064 15268
rect 10996 15219 11013 15253
rect 11013 15219 11047 15253
rect 11047 15219 11064 15253
rect 10996 15206 11064 15219
rect 11980 15209 12048 15222
rect 11980 15175 11997 15209
rect 11997 15175 12048 15209
rect 11980 15160 12048 15175
rect 9878 14499 9944 14512
rect 9878 14465 9925 14499
rect 9925 14465 9944 14499
rect 9878 14446 9944 14465
rect 9548 14299 9620 14318
rect 9548 14265 9563 14299
rect 9563 14265 9597 14299
rect 9597 14265 9620 14299
rect 9548 14248 9620 14265
rect 6828 13856 6896 13918
rect 7652 13882 7704 13936
rect 9896 13842 9956 13904
rect 4884 13700 4956 13770
rect 9750 13755 9822 13774
rect 5862 13692 5930 13754
rect 7656 13676 7724 13738
rect 9750 13721 9781 13755
rect 9781 13721 9822 13755
rect 9750 13704 9822 13721
rect 5984 13390 6052 13450
rect 4576 13318 4648 13384
rect 7136 13316 7204 13378
rect 9442 13375 9514 13388
rect 9442 13341 9457 13375
rect 9457 13341 9491 13375
rect 9491 13341 9514 13375
rect 9442 13322 9514 13341
rect 10660 14709 10728 14720
rect 10660 14675 10679 14709
rect 10679 14675 10728 14709
rect 16453 17157 16521 17172
rect 15691 17119 15759 17134
rect 15691 17085 15722 17119
rect 15722 17085 15759 17119
rect 16453 17123 16466 17157
rect 16466 17123 16500 17157
rect 16500 17123 16521 17157
rect 16453 17110 16521 17123
rect 17343 17159 17411 17174
rect 17343 17125 17374 17159
rect 17374 17125 17411 17159
rect 17343 17112 17411 17125
rect 18101 17149 18169 17166
rect 18101 17115 18108 17149
rect 18108 17115 18142 17149
rect 18142 17115 18169 17149
rect 18101 17104 18169 17115
rect 15691 17072 15759 17085
rect 19217 17151 19285 17166
rect 19217 17117 19230 17151
rect 19230 17117 19264 17151
rect 19264 17117 19285 17151
rect 19217 17104 19285 17117
rect 20107 17153 20175 17168
rect 20107 17119 20138 17153
rect 20138 17119 20175 17153
rect 20107 17106 20175 17119
rect 20865 17143 20933 17160
rect 20865 17109 20872 17143
rect 20872 17109 20906 17143
rect 20906 17109 20933 17143
rect 20865 17098 20933 17109
rect 21473 17141 21541 17156
rect 21473 17107 21486 17141
rect 21486 17107 21520 17141
rect 21520 17107 21541 17141
rect 21473 17094 21541 17107
rect 22363 17143 22431 17158
rect 22363 17109 22394 17143
rect 22394 17109 22431 17143
rect 22363 17096 22431 17109
rect 23121 17133 23189 17150
rect 23121 17099 23128 17133
rect 23128 17099 23162 17133
rect 23162 17099 23189 17133
rect 23121 17088 23189 17099
rect 16430 16660 16498 16722
rect 17188 16652 17256 16714
rect 18078 16654 18146 16716
rect 18686 16650 18754 16712
rect 19444 16642 19512 16704
rect 20334 16644 20402 16706
rect 21450 16644 21518 16706
rect 22208 16636 22276 16698
rect 23098 16638 23166 16700
rect 16410 16122 16478 16184
rect 17196 16112 17264 16174
rect 18076 16112 18144 16174
rect 18666 16112 18734 16174
rect 19452 16102 19520 16164
rect 20332 16102 20400 16164
rect 21430 16106 21498 16168
rect 22216 16096 22284 16158
rect 23096 16096 23164 16158
rect 24400 14810 24462 14870
rect 10660 14658 10728 14675
rect 11216 14287 11284 14298
rect 11216 14253 11271 14287
rect 11271 14253 11284 14287
rect 11216 14236 11284 14253
rect 24144 14662 24196 14714
rect 12782 14271 12850 14288
rect 12782 14237 12801 14271
rect 12801 14237 12835 14271
rect 12835 14237 12850 14271
rect 12782 14226 12850 14237
rect 24452 14552 24504 14564
rect 24452 14518 24456 14552
rect 24456 14518 24492 14552
rect 24492 14518 24504 14552
rect 24452 14512 24504 14518
rect 24552 14554 24556 14578
rect 24556 14554 24592 14578
rect 24592 14554 24604 14578
rect 24552 14526 24604 14554
rect 24698 14562 24750 14602
rect 24698 14550 24712 14562
rect 24712 14550 24746 14562
rect 24746 14550 24750 14562
rect 23992 14258 24054 14318
rect 10164 13308 10226 13360
rect 10878 13884 10930 13894
rect 10878 13850 10886 13884
rect 10886 13850 10920 13884
rect 10920 13850 10930 13884
rect 10878 13842 10930 13850
rect 10976 13924 11028 13934
rect 10976 13890 10984 13924
rect 10984 13890 11018 13924
rect 11018 13890 11028 13924
rect 10976 13882 11028 13890
rect 11074 13834 11126 13890
rect 11694 13913 11762 13922
rect 11694 13879 11723 13913
rect 11723 13879 11762 13913
rect 11694 13860 11762 13879
rect 12518 13886 12570 13940
rect 12732 13964 12812 13984
rect 12732 13922 12746 13964
rect 12746 13922 12796 13964
rect 12796 13922 12812 13964
rect 12732 13908 12812 13922
rect 10728 13743 10796 13758
rect 10728 13709 10753 13743
rect 10753 13709 10796 13743
rect 10728 13696 10796 13709
rect 12522 13680 12590 13742
rect 10850 13445 10918 13454
rect 10850 13411 10877 13445
rect 10877 13411 10918 13445
rect 10850 13394 10918 13411
rect 11006 13338 11060 13342
rect 11006 13302 11012 13338
rect 11012 13302 11048 13338
rect 11048 13302 11060 13338
rect 11006 13290 11060 13302
rect 12002 13369 12070 13382
rect 12002 13335 12057 13369
rect 12057 13335 12070 13369
rect 12002 13320 12070 13335
rect 5996 12856 6064 12916
rect 11062 13070 11114 13086
rect 11062 13036 11098 13070
rect 11098 13036 11114 13070
rect 11062 13032 11114 13036
rect 4990 12778 5062 12844
rect 9856 12831 9928 12848
rect 9856 12797 9859 12831
rect 9859 12797 9917 12831
rect 9917 12797 9928 12831
rect 9856 12782 9928 12797
rect 4634 12576 4708 12642
rect 9500 12631 9574 12646
rect 9500 12597 9555 12631
rect 9555 12597 9574 12631
rect 9500 12580 9574 12597
rect 6280 12370 6348 12432
rect 9872 12326 9934 12394
rect 10862 12901 10930 12920
rect 10862 12867 10877 12901
rect 10877 12867 10930 12901
rect 10862 12860 10930 12867
rect 11146 12425 11214 12436
rect 11146 12391 11149 12425
rect 11149 12391 11207 12425
rect 11207 12391 11214 12425
rect 11146 12374 11214 12391
rect 11206 12200 11258 12212
rect 11206 12166 11212 12200
rect 11212 12166 11246 12200
rect 11246 12166 11258 12200
rect 11206 12160 11258 12166
rect 4906 12034 4980 12100
rect 9772 12087 9846 12104
rect 9772 12053 9773 12087
rect 9773 12053 9831 12087
rect 9831 12053 9846 12087
rect 9772 12038 9846 12053
rect 11016 12114 11068 12122
rect 11016 12080 11024 12114
rect 11024 12080 11060 12114
rect 11060 12080 11068 12114
rect 11016 12070 11068 12080
rect 6002 11830 6070 11892
rect 4560 11756 4640 11820
rect 9426 11811 9506 11824
rect 9426 11777 9467 11811
rect 9467 11777 9501 11811
rect 9501 11777 9506 11811
rect 9426 11760 9506 11777
rect 10868 11881 10936 11896
rect 10868 11847 10873 11881
rect 10873 11847 10931 11881
rect 10931 11847 10936 11881
rect 10868 11834 10936 11847
rect 4994 11214 5074 11278
rect 9860 11267 9940 11282
rect 9860 11233 9869 11267
rect 9869 11233 9927 11267
rect 9927 11233 9940 11267
rect 9860 11218 9940 11233
rect 4626 11010 4706 11074
rect 9492 11067 9572 11078
rect 9492 11033 9507 11067
rect 9507 11033 9565 11067
rect 9565 11033 9572 11067
rect 9492 11014 9572 11033
rect 5054 10676 5108 10732
rect 9920 10680 9974 10736
rect 4904 10476 4984 10540
rect 9770 10523 9850 10544
rect 9770 10489 9783 10523
rect 9783 10489 9841 10523
rect 9841 10489 9850 10523
rect 9770 10480 9850 10489
rect 6226 6617 6282 6638
rect 6226 6583 6233 6617
rect 6233 6583 6267 6617
rect 6267 6583 6282 6617
rect 6226 6580 6282 6583
rect 6168 6382 6220 6390
rect 6168 6348 6178 6382
rect 6178 6348 6212 6382
rect 6212 6348 6220 6382
rect 6168 6338 6220 6348
rect 6268 6384 6320 6396
rect 6268 6350 6274 6384
rect 6274 6350 6308 6384
rect 6308 6350 6320 6384
rect 6268 6344 6320 6350
rect 6170 6073 6226 6088
rect 6170 6039 6175 6073
rect 6175 6039 6226 6073
rect 6170 6030 6226 6039
rect 10406 5985 10464 6002
rect 10774 5985 10832 6000
rect 10406 5951 10415 5985
rect 10415 5951 10449 5985
rect 10449 5951 10464 5985
rect 10774 5951 10783 5985
rect 10783 5951 10817 5985
rect 10817 5951 10832 5985
rect 10406 5940 10464 5951
rect 10774 5936 10832 5951
rect 12796 5973 12852 5986
rect 12796 5939 12845 5973
rect 12845 5939 12852 5973
rect 12796 5928 12852 5939
rect 14754 5981 14810 5994
rect 14754 5947 14803 5981
rect 14803 5947 14810 5981
rect 14754 5936 14810 5947
rect 16748 5987 16804 6000
rect 16748 5953 16797 5987
rect 16797 5953 16804 5987
rect 16748 5942 16804 5953
rect 2564 5565 2620 5578
rect 2564 5531 2601 5565
rect 2601 5531 2620 5565
rect 2564 5520 2620 5531
rect 4686 5557 4742 5570
rect 4686 5523 4735 5557
rect 4735 5523 4742 5557
rect 4686 5512 4742 5523
rect 6638 5557 6694 5570
rect 6638 5523 6687 5557
rect 6687 5523 6694 5557
rect 6638 5512 6694 5523
rect 8640 5563 8696 5576
rect 8640 5529 8689 5563
rect 8689 5529 8696 5563
rect 10410 5614 10462 5618
rect 10410 5580 10418 5614
rect 10418 5580 10452 5614
rect 10452 5580 10462 5614
rect 10410 5566 10462 5580
rect 8640 5518 8696 5529
rect 11214 5441 11270 5452
rect 11214 5407 11243 5441
rect 11243 5407 11270 5441
rect 11214 5394 11270 5407
rect 12800 5429 12856 5440
rect 12800 5395 12845 5429
rect 12845 5395 12856 5429
rect 12800 5382 12856 5395
rect 14758 5437 14814 5448
rect 14758 5403 14803 5437
rect 14803 5403 14814 5437
rect 14758 5390 14814 5403
rect 16752 5443 16808 5454
rect 16752 5409 16797 5443
rect 16797 5409 16808 5443
rect 16752 5396 16808 5409
rect 18726 5364 18784 5428
rect 2228 5194 2280 5198
rect 2228 5160 2236 5194
rect 2236 5160 2270 5194
rect 2270 5160 2280 5194
rect 2228 5146 2280 5160
rect 10188 5111 10244 5120
rect 10188 5077 10201 5111
rect 10201 5077 10244 5111
rect 10188 5062 10244 5077
rect 13032 5067 13088 5080
rect 2584 5021 2640 5040
rect 2584 4987 2601 5021
rect 2601 4987 2635 5021
rect 2635 4987 2640 5021
rect 2584 4982 2640 4987
rect 4690 5013 4746 5024
rect 4690 4979 4735 5013
rect 4735 4979 4746 5013
rect 4690 4966 4746 4979
rect 6642 5013 6698 5024
rect 6642 4979 6687 5013
rect 6687 4979 6698 5013
rect 6642 4966 6698 4979
rect 8644 5019 8700 5030
rect 8644 4985 8689 5019
rect 8689 4985 8700 5019
rect 8644 4972 8700 4985
rect 13032 5033 13081 5067
rect 13081 5033 13088 5067
rect 13032 5022 13088 5033
rect 15034 5061 15090 5074
rect 15034 5027 15083 5061
rect 15083 5027 15090 5061
rect 15034 5016 15090 5027
rect 10438 4740 10490 4744
rect 10438 4706 10446 4740
rect 10446 4706 10480 4740
rect 10480 4706 10490 4740
rect 10438 4692 10490 4706
rect 17056 5043 17112 5056
rect 17056 5009 17105 5043
rect 17105 5009 17112 5043
rect 17056 4998 17112 5009
rect 19056 5042 19108 5050
rect 19056 5004 19064 5042
rect 19064 5004 19102 5042
rect 19102 5004 19108 5042
rect 19056 4998 19108 5004
rect 10788 4567 10844 4580
rect 10440 4533 10443 4566
rect 10443 4533 10477 4566
rect 10477 4533 10492 4566
rect 10788 4533 10811 4567
rect 10811 4533 10844 4567
rect 10440 4512 10492 4533
rect 10788 4522 10844 4533
rect 13036 4523 13092 4534
rect 13036 4489 13081 4523
rect 13081 4489 13092 4523
rect 13036 4476 13092 4489
rect 18720 4816 18778 4880
rect 15038 4517 15094 4528
rect 15038 4483 15083 4517
rect 15083 4483 15094 4517
rect 15038 4470 15094 4483
rect 17060 4499 17116 4510
rect 17060 4465 17105 4499
rect 17105 4465 17116 4499
rect 17060 4452 17116 4465
rect 6194 3320 6254 3382
rect 6138 3122 6190 3130
rect 6138 3088 6148 3122
rect 6148 3088 6182 3122
rect 6182 3088 6190 3122
rect 6138 3078 6190 3088
rect 6238 3124 6290 3136
rect 6238 3090 6244 3124
rect 6244 3090 6278 3124
rect 6278 3090 6290 3124
rect 6238 3084 6290 3090
rect 6176 2766 6236 2828
rect 2604 2305 2660 2318
rect 2604 2271 2605 2305
rect 2605 2271 2660 2305
rect 2604 2260 2660 2271
rect 4592 2301 4648 2314
rect 4592 2267 4641 2301
rect 4641 2267 4648 2301
rect 4592 2256 4648 2267
rect 6544 2301 6600 2314
rect 6544 2267 6593 2301
rect 6593 2267 6600 2301
rect 6544 2256 6600 2267
rect 8546 2307 8602 2320
rect 8546 2273 8595 2307
rect 8595 2273 8602 2307
rect 8546 2262 8602 2273
rect 10498 2307 10554 2320
rect 10498 2273 10547 2307
rect 10547 2273 10554 2307
rect 10498 2262 10554 2273
rect 12490 2307 12546 2320
rect 12490 2273 12539 2307
rect 12539 2273 12546 2307
rect 12490 2262 12546 2273
rect 14442 2307 14498 2320
rect 14442 2273 14491 2307
rect 14491 2273 14498 2307
rect 14442 2262 14498 2273
rect 16506 2307 16562 2320
rect 16506 2273 16555 2307
rect 16555 2273 16562 2307
rect 16506 2262 16562 2273
rect 2198 1934 2250 1938
rect 2198 1900 2206 1934
rect 2206 1900 2240 1934
rect 2240 1900 2250 1934
rect 2198 1886 2250 1900
rect 17402 1876 17454 1930
rect 2604 1761 2656 1778
rect 2604 1727 2605 1761
rect 2605 1727 2656 1761
rect 2604 1720 2656 1727
rect 4596 1757 4652 1768
rect 4596 1723 4641 1757
rect 4641 1723 4652 1757
rect 6548 1757 6604 1768
rect 4596 1710 4652 1723
rect 6548 1723 6593 1757
rect 6593 1723 6604 1757
rect 8550 1763 8606 1774
rect 6548 1710 6604 1723
rect 8550 1729 8595 1763
rect 8595 1729 8606 1763
rect 10502 1763 10558 1774
rect 10502 1729 10547 1763
rect 10547 1729 10558 1763
rect 12494 1763 12550 1774
rect 8550 1716 8606 1729
rect 10502 1716 10558 1729
rect 12494 1729 12539 1763
rect 12539 1729 12550 1763
rect 14446 1763 14502 1774
rect 12494 1716 12550 1729
rect 14446 1729 14491 1763
rect 14491 1729 14502 1763
rect 16510 1763 16566 1774
rect 14446 1716 14502 1729
rect 16510 1729 16555 1763
rect 16555 1729 16566 1763
rect 16510 1716 16566 1729
<< metal2 >>
rect 18590 44096 19128 44168
rect 18590 43898 18768 44096
rect 18962 43898 19128 44096
rect 18590 43828 19128 43898
rect 18554 42820 18644 43002
rect 18554 42762 18562 42820
rect 18624 42762 18644 42820
rect 18554 42576 18644 42762
rect 19118 42782 19208 42956
rect 19118 42724 19124 42782
rect 19186 42724 19208 42782
rect 19118 42530 19208 42724
rect 18530 40948 18620 41118
rect 18530 40890 18540 40948
rect 18602 40890 18620 40948
rect 18530 40692 18620 40890
rect 19090 40940 19180 41096
rect 19090 40882 19106 40940
rect 19168 40882 19180 40940
rect 19090 40670 19180 40882
rect 18548 39320 18638 39512
rect 18548 39262 18564 39320
rect 18626 39262 18638 39320
rect 18548 39086 18638 39262
rect 19092 39316 19182 39484
rect 19092 39258 19106 39316
rect 19168 39258 19182 39316
rect 19092 39058 19182 39258
rect 18558 38124 18648 38298
rect 18558 38066 18572 38124
rect 18634 38066 18648 38124
rect 18558 37872 18648 38066
rect 19106 38140 19196 38320
rect 19106 38082 19122 38140
rect 19184 38082 19196 38140
rect 19106 37894 19196 38082
rect 18568 37054 18658 37240
rect 18568 36996 18580 37054
rect 18642 36996 18658 37054
rect 18568 36814 18658 36996
rect 19114 37044 19204 37230
rect 19114 36986 19128 37044
rect 19190 36986 19204 37044
rect 19114 36804 19204 36986
rect 19120 36284 19218 36320
rect 18574 36256 18670 36272
rect 18574 36200 18598 36256
rect 18656 36200 18670 36256
rect 18574 36178 18670 36200
rect 19120 36228 19142 36284
rect 19200 36228 19218 36284
rect 19120 36180 19218 36228
rect 18340 34458 18512 34648
rect 18340 34376 18374 34458
rect 18454 34454 18512 34458
rect 18340 34372 18424 34376
rect 18504 34372 18512 34454
rect 18340 34220 18512 34372
rect 18960 34458 19116 34626
rect 18960 34376 18972 34458
rect 19052 34376 19116 34458
rect 18960 34204 19116 34376
rect 18348 32152 18520 32342
rect 18348 32070 18382 32152
rect 18462 32148 18520 32152
rect 18348 32066 18432 32070
rect 18512 32066 18520 32148
rect 18348 31914 18520 32066
rect 18968 32152 19124 32320
rect 18968 32070 18980 32152
rect 19060 32070 19124 32152
rect 18968 31898 19124 32070
rect 18356 29938 18528 30128
rect 18356 29856 18390 29938
rect 18470 29934 18528 29938
rect 18356 29852 18440 29856
rect 18520 29852 18528 29934
rect 18356 29700 18528 29852
rect 18976 29938 19132 30106
rect 18976 29856 18988 29938
rect 19068 29856 19132 29938
rect 18976 29684 19132 29856
rect 18338 27738 18510 27928
rect 18338 27656 18372 27738
rect 18452 27734 18510 27738
rect 18338 27652 18422 27656
rect 18502 27652 18510 27734
rect 18338 27500 18510 27652
rect 18958 27738 19114 27906
rect 18958 27656 18970 27738
rect 19050 27656 19114 27738
rect 18958 27484 19114 27656
rect 18346 25524 18518 25714
rect 18346 25442 18380 25524
rect 18460 25520 18518 25524
rect 18346 25438 18430 25442
rect 18510 25438 18518 25520
rect 18346 25286 18518 25438
rect 18966 25524 19122 25692
rect 18966 25442 18978 25524
rect 19058 25442 19122 25524
rect 18966 25270 19122 25442
rect 8380 23480 8808 23514
rect 8380 23430 8536 23480
rect 8380 23350 8532 23430
rect 8618 23400 8808 23480
rect 8614 23350 8808 23400
rect 10594 23488 11022 23522
rect 10594 23438 10750 23488
rect 10594 23358 10746 23438
rect 10832 23408 11022 23488
rect 10828 23358 11022 23408
rect 10594 23350 11022 23358
rect 12794 23470 13222 23504
rect 12794 23420 12950 23470
rect 8380 23342 8808 23350
rect 12794 23340 12946 23420
rect 13032 23390 13222 23470
rect 13028 23340 13222 23390
rect 15008 23478 15436 23512
rect 15008 23428 15164 23478
rect 15008 23348 15160 23428
rect 15246 23398 15436 23478
rect 15242 23348 15436 23398
rect 17314 23486 17742 23520
rect 17314 23436 17470 23486
rect 17314 23356 17466 23436
rect 17552 23406 17742 23486
rect 17548 23356 17742 23406
rect 17314 23348 17742 23356
rect 15008 23340 15436 23348
rect 12794 23332 13222 23340
rect 8364 22882 8786 22894
rect 8364 22802 8536 22882
rect 8618 22802 8786 22882
rect 8364 22738 8786 22802
rect 10578 22890 11000 22902
rect 10578 22810 10750 22890
rect 10832 22810 11000 22890
rect 10578 22746 11000 22810
rect 12778 22872 13200 22884
rect 12778 22792 12950 22872
rect 13032 22792 13200 22872
rect 12778 22728 13200 22792
rect 14992 22880 15414 22892
rect 14992 22800 15164 22880
rect 15246 22800 15414 22880
rect 14992 22736 15414 22800
rect 17298 22888 17720 22900
rect 17298 22808 17470 22888
rect 17552 22808 17720 22888
rect 17298 22744 17720 22808
rect 9430 17822 9706 17844
rect 9430 17762 9540 17822
rect 9600 17762 9706 17822
rect 9430 17746 9706 17762
rect 16391 17714 16603 17732
rect 15609 17674 15821 17692
rect 15609 17612 15683 17674
rect 15751 17612 15821 17674
rect 16391 17652 16455 17714
rect 16523 17652 16603 17714
rect 16391 17640 16603 17652
rect 17261 17714 17473 17732
rect 17261 17652 17335 17714
rect 17403 17652 17473 17714
rect 17261 17640 17473 17652
rect 18051 17704 18263 17724
rect 18051 17642 18121 17704
rect 18189 17642 18263 17704
rect 18051 17632 18263 17642
rect 19155 17708 19367 17726
rect 19155 17646 19219 17708
rect 19287 17646 19367 17708
rect 19155 17634 19367 17646
rect 20025 17708 20237 17726
rect 20025 17646 20099 17708
rect 20167 17646 20237 17708
rect 20025 17634 20237 17646
rect 20815 17698 21027 17718
rect 20815 17636 20885 17698
rect 20953 17636 21027 17698
rect 20815 17626 21027 17636
rect 21411 17698 21623 17716
rect 21411 17636 21475 17698
rect 21543 17636 21623 17698
rect 21411 17624 21623 17636
rect 22281 17698 22493 17716
rect 22281 17636 22355 17698
rect 22423 17636 22493 17698
rect 22281 17624 22493 17636
rect 23071 17688 23283 17708
rect 23071 17626 23141 17688
rect 23209 17626 23283 17688
rect 23071 17616 23283 17626
rect 15609 17600 15821 17612
rect 6463 17587 6545 17588
rect 6463 17586 6759 17587
rect 6463 17576 6760 17586
rect 6463 17505 6646 17576
rect 4472 16624 4732 16636
rect 4472 16614 4590 16624
rect 4472 16558 4552 16614
rect 4642 16570 4732 16624
rect 4608 16558 4732 16570
rect 4472 16536 4732 16558
rect 4886 16076 5106 16090
rect 4886 16020 4976 16076
rect 5034 16020 5106 16076
rect 4886 15994 5106 16020
rect 4562 15874 4938 15880
rect 4562 15814 4746 15874
rect 4808 15814 4938 15874
rect 4562 15792 4938 15814
rect 6463 15424 6545 17505
rect 6604 17504 6646 17505
rect 6722 17504 6760 17576
rect 6604 17498 6760 17504
rect 9432 17278 9706 17302
rect 9432 17218 9536 17278
rect 9594 17218 9706 17278
rect 9432 17202 9706 17218
rect 16379 17172 16591 17186
rect 15619 17134 15831 17146
rect 15619 17072 15691 17134
rect 15759 17072 15831 17134
rect 16379 17110 16453 17172
rect 16521 17110 16591 17172
rect 16379 17094 16591 17110
rect 17271 17174 17483 17186
rect 17271 17112 17343 17174
rect 17411 17112 17483 17174
rect 17271 17094 17483 17112
rect 18041 17166 18253 17180
rect 18041 17104 18101 17166
rect 18169 17104 18253 17166
rect 18041 17088 18253 17104
rect 19143 17166 19355 17180
rect 19143 17104 19217 17166
rect 19285 17104 19355 17166
rect 19143 17088 19355 17104
rect 20035 17168 20247 17180
rect 20035 17106 20107 17168
rect 20175 17106 20247 17168
rect 20035 17088 20247 17106
rect 20805 17160 21017 17174
rect 20805 17098 20865 17160
rect 20933 17098 21017 17160
rect 20805 17082 21017 17098
rect 21399 17156 21611 17170
rect 21399 17094 21473 17156
rect 21541 17094 21611 17156
rect 21399 17078 21611 17094
rect 22291 17158 22503 17170
rect 22291 17096 22363 17158
rect 22431 17096 22503 17158
rect 22291 17078 22503 17096
rect 23061 17150 23273 17164
rect 23061 17088 23121 17150
rect 23189 17088 23273 17150
rect 23061 17072 23273 17088
rect 11401 17054 11483 17055
rect 15619 17054 15831 17072
rect 11400 17042 11506 17054
rect 11400 16986 11414 17042
rect 11474 17033 11506 17042
rect 11474 16986 11507 17033
rect 11400 16812 11507 16986
rect 11329 16730 11507 16812
rect 9338 16628 9598 16640
rect 9338 16618 9456 16628
rect 9338 16562 9418 16618
rect 9508 16574 9598 16628
rect 9474 16562 9598 16574
rect 9338 16540 9598 16562
rect 10812 16410 11014 16442
rect 10812 16344 10872 16410
rect 10942 16344 11014 16410
rect 10812 16316 11014 16344
rect 9752 16080 9972 16094
rect 9752 16024 9842 16080
rect 9900 16024 9972 16080
rect 9752 15998 9972 16024
rect 9428 15878 9804 15884
rect 9428 15818 9612 15878
rect 9674 15818 9804 15878
rect 9428 15796 9804 15818
rect 6608 15768 6894 15780
rect 6608 15706 6712 15768
rect 6780 15706 6894 15768
rect 6608 15684 6894 15706
rect 9824 15506 9932 15514
rect 9824 15452 9842 15506
rect 9896 15476 9932 15506
rect 9896 15452 10324 15476
rect 9824 15440 10324 15452
rect 6463 15408 6682 15424
rect 6463 15356 6608 15408
rect 6660 15356 6682 15408
rect 4836 15332 5028 15350
rect 6463 15342 6682 15356
rect 4836 15270 4898 15332
rect 4966 15270 5028 15332
rect 9702 15336 9894 15354
rect 4836 15254 5028 15270
rect 6108 15264 6254 15280
rect 6108 15202 6130 15264
rect 6198 15202 6254 15264
rect 9702 15274 9764 15336
rect 9832 15274 9894 15336
rect 9702 15258 9894 15274
rect 6108 15184 6254 15202
rect 7046 15218 7252 15238
rect 7046 15156 7114 15218
rect 7182 15156 7252 15218
rect 7046 15140 7252 15156
rect 4476 15052 4750 15070
rect 4476 14986 4582 15052
rect 4648 14986 4750 15052
rect 4476 14978 4750 14986
rect 9342 15056 9616 15074
rect 9342 14990 9448 15056
rect 9514 14990 9616 15056
rect 9342 14982 9616 14990
rect 5748 14716 5908 14736
rect 5748 14654 5794 14716
rect 5862 14654 5908 14716
rect 5748 14640 5908 14654
rect 4946 14508 5118 14524
rect 4946 14442 5012 14508
rect 5078 14442 5118 14508
rect 4946 14434 5118 14442
rect 7635 14487 8531 14581
rect 4576 14314 4870 14320
rect 4576 14244 4682 14314
rect 4754 14244 4870 14314
rect 4576 14232 4870 14244
rect 6322 14294 6470 14316
rect 6322 14232 6350 14294
rect 6418 14232 6470 14294
rect 6322 14218 6470 14232
rect 7635 13974 7729 14487
rect 7840 14284 8072 14296
rect 7840 14222 7916 14284
rect 7984 14222 8072 14284
rect 7840 14204 8072 14222
rect 6794 13918 6946 13938
rect 6794 13856 6828 13918
rect 6896 13856 6946 13918
rect 7635 13936 7806 13974
rect 7635 13882 7652 13936
rect 7704 13882 7806 13936
rect 7635 13857 7806 13882
rect 7724 13856 7806 13857
rect 6794 13842 6946 13856
rect 4820 13770 5040 13780
rect 4820 13700 4884 13770
rect 4956 13700 5040 13770
rect 4820 13684 5040 13700
rect 5824 13754 5974 13770
rect 5824 13692 5862 13754
rect 5930 13692 5974 13754
rect 5824 13672 5974 13692
rect 7642 13738 7744 13754
rect 7642 13676 7656 13738
rect 7724 13676 7744 13738
rect 7642 13658 7744 13676
rect 5950 13450 6084 13470
rect 4468 13384 4738 13396
rect 4468 13318 4576 13384
rect 4648 13318 4738 13384
rect 5950 13390 5984 13450
rect 6052 13390 6084 13450
rect 5950 13378 6084 13390
rect 7096 13378 7248 13396
rect 4468 13310 4738 13318
rect 7096 13316 7136 13378
rect 7204 13316 7248 13378
rect 7096 13300 7248 13316
rect 5948 12916 6100 12928
rect 5948 12856 5996 12916
rect 6064 12856 6100 12916
rect 4922 12844 5112 12854
rect 4922 12778 4990 12844
rect 5062 12778 5112 12844
rect 5948 12834 6100 12856
rect 4922 12766 5112 12778
rect 4574 12642 4780 12654
rect 4574 12576 4634 12642
rect 4708 12576 4780 12642
rect 4574 12560 4780 12576
rect 6230 12432 6402 12452
rect 6230 12370 6280 12432
rect 6348 12370 6402 12432
rect 6230 12356 6402 12370
rect 4858 12100 5024 12116
rect 4858 12034 4906 12100
rect 4980 12034 5024 12100
rect 4858 12022 5024 12034
rect 5944 11892 6100 11908
rect 4510 11820 4690 11834
rect 4510 11756 4560 11820
rect 4640 11756 4690 11820
rect 5944 11830 6002 11892
rect 6070 11830 6100 11892
rect 5944 11812 6100 11830
rect 4510 11746 4690 11756
rect 4938 11278 5118 11292
rect 4938 11214 4994 11278
rect 5074 11214 5118 11278
rect 4938 11204 5118 11214
rect 4580 11074 4776 11092
rect 4580 11010 4626 11074
rect 4706 11010 4776 11074
rect 4580 10996 4776 11010
rect 8437 10762 8531 14487
rect 9812 14512 9984 14528
rect 9812 14446 9878 14512
rect 9944 14446 9984 14512
rect 9812 14438 9984 14446
rect 9442 14318 9736 14324
rect 9442 14248 9548 14318
rect 9620 14248 9736 14318
rect 9442 14236 9736 14248
rect 10288 14102 10324 15440
rect 10614 14720 10774 14740
rect 10614 14658 10660 14720
rect 10728 14658 10774 14720
rect 10614 14644 10774 14658
rect 10876 14514 10944 16316
rect 11329 15428 11411 16730
rect 16346 16722 16558 16738
rect 16346 16660 16430 16722
rect 16498 16660 16558 16722
rect 16346 16646 16558 16660
rect 17116 16714 17328 16732
rect 17116 16652 17188 16714
rect 17256 16652 17328 16714
rect 17116 16640 17328 16652
rect 18008 16716 18220 16732
rect 18008 16654 18078 16716
rect 18146 16654 18220 16716
rect 18008 16640 18220 16654
rect 18602 16712 18814 16728
rect 18602 16650 18686 16712
rect 18754 16650 18814 16712
rect 18602 16636 18814 16650
rect 19372 16704 19584 16722
rect 19372 16642 19444 16704
rect 19512 16642 19584 16704
rect 19372 16630 19584 16642
rect 20264 16706 20476 16722
rect 20264 16644 20334 16706
rect 20402 16644 20476 16706
rect 20264 16630 20476 16644
rect 21366 16706 21578 16722
rect 21366 16644 21450 16706
rect 21518 16644 21578 16706
rect 21366 16630 21578 16644
rect 22136 16698 22348 16716
rect 22136 16636 22208 16698
rect 22276 16636 22348 16698
rect 22136 16624 22348 16636
rect 23028 16700 23240 16716
rect 23028 16638 23098 16700
rect 23166 16638 23240 16700
rect 23028 16624 23240 16638
rect 16336 16184 16548 16194
rect 16336 16122 16410 16184
rect 16478 16122 16548 16184
rect 16336 16102 16548 16122
rect 17126 16174 17338 16186
rect 17126 16112 17196 16174
rect 17264 16112 17338 16174
rect 17126 16094 17338 16112
rect 17996 16174 18208 16186
rect 17996 16112 18076 16174
rect 18144 16112 18208 16174
rect 17996 16094 18208 16112
rect 18592 16174 18804 16184
rect 18592 16112 18666 16174
rect 18734 16112 18804 16174
rect 18592 16092 18804 16112
rect 19382 16164 19594 16176
rect 19382 16102 19452 16164
rect 19520 16102 19594 16164
rect 19382 16084 19594 16102
rect 20252 16164 20464 16176
rect 20252 16102 20332 16164
rect 20400 16102 20464 16164
rect 20252 16084 20464 16102
rect 21356 16168 21568 16178
rect 21356 16106 21430 16168
rect 21498 16106 21568 16168
rect 21356 16086 21568 16106
rect 22146 16158 22358 16170
rect 22146 16096 22216 16158
rect 22284 16096 22358 16158
rect 22146 16078 22358 16096
rect 23016 16158 23228 16170
rect 23016 16096 23096 16158
rect 23164 16096 23228 16158
rect 23016 16078 23228 16096
rect 11474 15772 11760 15784
rect 11474 15710 11578 15772
rect 11646 15710 11760 15772
rect 11474 15688 11760 15710
rect 11329 15412 11548 15428
rect 11329 15360 11474 15412
rect 11526 15360 11548 15412
rect 11329 15346 11548 15360
rect 10974 15268 11120 15284
rect 10974 15206 10996 15268
rect 11064 15206 11120 15268
rect 10974 15188 11120 15206
rect 11912 15222 12118 15242
rect 11912 15160 11980 15222
rect 12048 15160 12118 15222
rect 11912 15144 12118 15160
rect 24312 14870 24542 14880
rect 24312 14810 24400 14870
rect 24462 14810 24542 14870
rect 24312 14788 24542 14810
rect 26389 14843 27464 14921
rect 26389 14740 26467 14843
rect 26948 14766 27172 14794
rect 26389 14726 26466 14740
rect 24138 14714 26466 14726
rect 24138 14662 24144 14714
rect 24196 14662 26466 14714
rect 24138 14658 26466 14662
rect 10876 14446 11034 14514
rect 10288 14066 10898 14102
rect 10862 13940 10898 14066
rect 9834 13904 10004 13916
rect 9834 13842 9896 13904
rect 9956 13884 10004 13904
rect 10862 13894 10938 13940
rect 10862 13884 10878 13894
rect 9956 13842 10580 13884
rect 9834 13836 10580 13842
rect 10860 13842 10878 13884
rect 10930 13842 10938 13894
rect 10860 13836 10938 13842
rect 9834 13822 10004 13836
rect 9686 13774 9906 13784
rect 9686 13704 9750 13774
rect 9822 13704 9906 13774
rect 9686 13688 9906 13704
rect 10530 13596 10578 13836
rect 10868 13798 10938 13836
rect 10966 13934 11034 14446
rect 12501 14491 13397 14585
rect 24138 14578 24198 14658
rect 26389 14657 26466 14658
rect 26948 14646 27000 14766
rect 27122 14726 27172 14766
rect 27122 14658 27176 14726
rect 27122 14646 27172 14658
rect 11188 14298 11336 14320
rect 11188 14236 11216 14298
rect 11284 14236 11336 14298
rect 11188 14222 11336 14236
rect 10966 13882 10976 13934
rect 11028 13882 11034 13934
rect 10966 13796 11034 13882
rect 11067 13890 11141 13989
rect 12501 13978 12595 14491
rect 12706 14288 12938 14300
rect 12706 14226 12782 14288
rect 12850 14226 12938 14288
rect 12706 14208 12938 14226
rect 12704 13984 12842 13996
rect 11067 13834 11074 13890
rect 11126 13834 11141 13890
rect 11660 13922 11812 13942
rect 11660 13860 11694 13922
rect 11762 13860 11812 13922
rect 12501 13940 12672 13978
rect 12501 13886 12518 13940
rect 12570 13886 12672 13940
rect 12704 13908 12732 13984
rect 12812 13908 12842 13984
rect 12704 13894 12842 13908
rect 12501 13861 12672 13886
rect 12590 13860 12672 13861
rect 11660 13846 11812 13860
rect 11067 13805 11141 13834
rect 10690 13758 10840 13774
rect 10690 13696 10728 13758
rect 10796 13696 10840 13758
rect 11067 13731 11209 13805
rect 10690 13676 10840 13696
rect 10530 13548 11040 13596
rect 10816 13454 10950 13474
rect 9334 13388 9604 13400
rect 9334 13322 9442 13388
rect 9514 13322 9604 13388
rect 10816 13394 10850 13454
rect 10918 13394 10950 13454
rect 10816 13382 10950 13394
rect 10992 13376 11040 13548
rect 10226 13370 10632 13372
rect 9334 13314 9604 13322
rect 10156 13360 10632 13370
rect 10156 13308 10164 13360
rect 10226 13308 10632 13360
rect 10156 13300 10632 13308
rect 10560 13174 10632 13300
rect 10986 13342 11084 13376
rect 10986 13290 11006 13342
rect 11060 13290 11084 13342
rect 10986 13272 11084 13290
rect 11135 13176 11209 13731
rect 12508 13742 12610 13758
rect 12508 13680 12522 13742
rect 12590 13680 12610 13742
rect 12508 13662 12610 13680
rect 12724 13660 12792 13894
rect 12704 13658 12792 13660
rect 12644 13590 12792 13658
rect 11962 13382 12114 13400
rect 11962 13320 12002 13382
rect 12070 13320 12114 13382
rect 11962 13304 12114 13320
rect 11006 13174 11209 13176
rect 10560 13102 11209 13174
rect 11052 13086 11124 13102
rect 11052 13032 11062 13086
rect 11114 13032 11124 13086
rect 11052 12948 11124 13032
rect 10814 12920 10966 12932
rect 10814 12860 10862 12920
rect 10930 12860 10966 12920
rect 9788 12848 9978 12858
rect 9788 12782 9856 12848
rect 9928 12782 9978 12848
rect 10814 12838 10966 12860
rect 9788 12770 9978 12782
rect 9440 12646 9646 12658
rect 9440 12580 9500 12646
rect 9574 12580 9646 12646
rect 9440 12564 9646 12580
rect 11096 12436 11268 12456
rect 9826 12394 9976 12408
rect 9826 12326 9872 12394
rect 9934 12342 9976 12394
rect 11096 12374 11146 12436
rect 11214 12374 11268 12436
rect 11096 12360 11268 12374
rect 9934 12326 11056 12342
rect 9826 12310 11056 12326
rect 11024 12130 11056 12310
rect 12644 12222 12712 13590
rect 11200 12212 12712 12222
rect 11200 12160 11206 12212
rect 11258 12160 12712 12212
rect 11200 12154 12712 12160
rect 11008 12122 11078 12130
rect 9724 12104 9890 12120
rect 9724 12038 9772 12104
rect 9846 12038 9890 12104
rect 11008 12070 11016 12122
rect 11068 12070 11078 12122
rect 11008 12064 11078 12070
rect 9724 12026 9890 12038
rect 10810 11896 10966 11912
rect 9376 11824 9556 11838
rect 9376 11760 9426 11824
rect 9506 11760 9556 11824
rect 10810 11834 10868 11896
rect 10936 11834 10966 11896
rect 10810 11816 10966 11834
rect 9376 11750 9556 11760
rect 9804 11282 9984 11296
rect 9804 11218 9860 11282
rect 9940 11218 9984 11282
rect 9804 11208 9984 11218
rect 9446 11078 9642 11096
rect 9446 11014 9492 11078
rect 9572 11014 9642 11078
rect 9446 11000 9642 11014
rect 13303 10766 13397 14491
rect 24448 14564 24504 14620
rect 24448 14512 24452 14564
rect 23850 14318 24212 14334
rect 23850 14258 23992 14318
rect 24054 14258 24212 14318
rect 23850 14240 24212 14258
rect 24448 14112 24504 14512
rect 24546 14578 24606 14622
rect 24546 14526 24552 14578
rect 24604 14526 24606 14578
rect 24448 14056 24502 14112
rect 4970 10732 8531 10762
rect 4970 10676 5054 10732
rect 5108 10676 8531 10732
rect 4970 10668 8531 10676
rect 9836 10736 13397 10766
rect 9836 10680 9920 10736
rect 9974 10680 13397 10736
rect 9836 10672 13397 10680
rect 23258 14000 24502 14056
rect 4970 10652 5202 10668
rect 9836 10656 10068 10672
rect 4856 10540 5036 10546
rect 4856 10476 4904 10540
rect 4984 10476 5036 10540
rect 4856 10458 5036 10476
rect 9722 10544 9902 10550
rect 9722 10480 9770 10544
rect 9850 10480 9902 10544
rect 9722 10462 9902 10480
rect 6112 6638 6388 6648
rect 6112 6580 6226 6638
rect 6282 6580 6388 6638
rect 6112 6558 6388 6580
rect 5585 6398 5651 6404
rect 2222 6390 6228 6398
rect 2222 6338 6168 6390
rect 6220 6338 6228 6390
rect 6262 6396 13156 6398
rect 6262 6344 6268 6396
rect 6320 6394 13156 6396
rect 23258 6394 23314 14000
rect 24546 13290 24606 14526
rect 24685 14602 24870 14619
rect 26948 14604 27172 14646
rect 24685 14550 24698 14602
rect 24750 14550 24870 14602
rect 24685 14541 24870 14550
rect 24685 14499 24763 14541
rect 24792 14514 24870 14541
rect 26993 14514 27071 14604
rect 24792 14436 27071 14514
rect 27386 14514 27464 14843
rect 27386 14510 27604 14514
rect 27386 14492 27730 14510
rect 27386 14436 27550 14492
rect 27512 14372 27550 14436
rect 27682 14372 27730 14492
rect 27512 14336 27730 14372
rect 6320 6344 23314 6394
rect 6262 6340 23314 6344
rect 6262 6338 16050 6340
rect 17150 6338 23314 6340
rect 24252 13230 24608 13290
rect 2222 6332 6228 6338
rect 18793 6336 18848 6338
rect 2222 5198 2290 6332
rect 6110 6088 6274 6104
rect 6110 6030 6170 6088
rect 6226 6030 6274 6088
rect 6110 6018 6274 6030
rect 10404 6002 10472 6018
rect 10404 5940 10406 6002
rect 10464 5940 10472 6002
rect 10404 5618 10472 5940
rect 10708 6000 10888 6016
rect 10708 5936 10774 6000
rect 10832 5936 10888 6000
rect 10708 5922 10888 5936
rect 12738 5986 12918 6002
rect 12738 5928 12796 5986
rect 12852 5928 12918 5986
rect 12738 5908 12918 5928
rect 14696 5994 14876 6010
rect 14696 5936 14754 5994
rect 14810 5936 14876 5994
rect 14696 5916 14876 5936
rect 16690 6000 16870 6016
rect 16690 5942 16748 6000
rect 16804 5942 16870 6000
rect 16690 5922 16870 5942
rect 2510 5578 2690 5596
rect 2510 5520 2564 5578
rect 2620 5520 2690 5578
rect 2510 5502 2690 5520
rect 4628 5570 4808 5586
rect 4628 5512 4686 5570
rect 4742 5512 4808 5570
rect 4628 5492 4808 5512
rect 6580 5570 6760 5586
rect 6580 5512 6638 5570
rect 6694 5512 6760 5570
rect 6580 5492 6760 5512
rect 8582 5576 8762 5592
rect 8582 5518 8640 5576
rect 8696 5518 8762 5576
rect 10404 5566 10410 5618
rect 10462 5566 10472 5618
rect 10404 5562 10472 5566
rect 8582 5498 8762 5518
rect 11142 5452 11324 5474
rect 11142 5394 11214 5452
rect 11270 5394 11324 5452
rect 11142 5378 11324 5394
rect 12738 5440 12918 5458
rect 12738 5382 12800 5440
rect 12856 5382 12918 5440
rect 12738 5364 12918 5382
rect 14696 5448 14876 5466
rect 14696 5390 14758 5448
rect 14814 5390 14876 5448
rect 14696 5372 14876 5390
rect 16690 5454 16870 5472
rect 16690 5396 16752 5454
rect 16808 5396 16870 5454
rect 16690 5378 16870 5396
rect 18658 5428 18838 5444
rect 18658 5364 18726 5428
rect 18784 5364 18838 5428
rect 18658 5348 18838 5364
rect 2222 5146 2228 5198
rect 2280 5146 2290 5198
rect 19193 5175 19248 6338
rect 2222 5142 2290 5146
rect 10128 5120 10308 5142
rect 10128 5062 10188 5120
rect 10244 5062 10308 5120
rect 19196 5098 19244 5175
rect 2520 5040 2700 5050
rect 2520 4982 2584 5040
rect 2640 4982 2700 5040
rect 2520 4956 2700 4982
rect 4628 5024 4808 5042
rect 4628 4966 4690 5024
rect 4746 4966 4808 5024
rect 4628 4948 4808 4966
rect 6580 5024 6760 5042
rect 6580 4966 6642 5024
rect 6698 4966 6760 5024
rect 6580 4948 6760 4966
rect 8582 5030 8762 5048
rect 10128 5046 10308 5062
rect 12974 5080 13154 5096
rect 8582 4972 8644 5030
rect 8700 4972 8762 5030
rect 12974 5022 13032 5080
rect 13088 5022 13154 5080
rect 12974 5002 13154 5022
rect 14976 5074 15156 5090
rect 14976 5016 15034 5074
rect 15090 5016 15156 5074
rect 14976 4996 15156 5016
rect 16998 5056 17178 5072
rect 16998 4998 17056 5056
rect 17112 4998 17178 5056
rect 16998 4978 17178 4998
rect 19048 5050 19244 5098
rect 19048 4998 19056 5050
rect 19108 4998 19112 5050
rect 8582 4954 8762 4972
rect 19048 4942 19112 4998
rect 18662 4880 18842 4894
rect 18662 4816 18720 4880
rect 18778 4816 18842 4880
rect 10432 4744 10500 4802
rect 18662 4798 18842 4816
rect 10432 4692 10438 4744
rect 10490 4692 10500 4744
rect 10432 4566 10500 4692
rect 10432 4512 10440 4566
rect 10492 4512 10500 4566
rect 10432 4502 10500 4512
rect 10734 4580 10914 4594
rect 10734 4522 10788 4580
rect 10844 4522 10914 4580
rect 10734 4498 10914 4522
rect 12974 4534 13154 4552
rect 12974 4476 13036 4534
rect 13092 4476 13154 4534
rect 12974 4458 13154 4476
rect 14976 4528 15156 4546
rect 14976 4470 15038 4528
rect 15094 4470 15156 4528
rect 14976 4452 15156 4470
rect 16998 4510 17178 4528
rect 16998 4452 17060 4510
rect 17116 4452 17178 4510
rect 16998 4434 17178 4452
rect 6082 3382 6354 3386
rect 6082 3320 6194 3382
rect 6254 3320 6354 3382
rect 6082 3292 6354 3320
rect 24252 3138 24312 13230
rect 2192 3130 6198 3138
rect 2192 3078 6138 3130
rect 6190 3078 6198 3130
rect 6232 3136 24312 3138
rect 6232 3084 6238 3136
rect 6290 3084 24312 3136
rect 6232 3078 24312 3084
rect 2192 3072 6198 3078
rect 2192 1938 2260 3072
rect 6080 2828 6300 2842
rect 6080 2766 6176 2828
rect 6236 2766 6300 2828
rect 6080 2752 6300 2766
rect 2540 2318 2720 2336
rect 2540 2260 2604 2318
rect 2660 2260 2720 2318
rect 2540 2242 2720 2260
rect 4534 2314 4714 2330
rect 4534 2256 4592 2314
rect 4648 2256 4714 2314
rect 4534 2236 4714 2256
rect 6486 2314 6666 2330
rect 6486 2256 6544 2314
rect 6600 2256 6666 2314
rect 6486 2236 6666 2256
rect 8488 2320 8668 2336
rect 8488 2262 8546 2320
rect 8602 2262 8668 2320
rect 8488 2242 8668 2262
rect 10440 2320 10620 2336
rect 10440 2262 10498 2320
rect 10554 2262 10620 2320
rect 10440 2242 10620 2262
rect 12432 2320 12612 2336
rect 12432 2262 12490 2320
rect 12546 2262 12612 2320
rect 12432 2242 12612 2262
rect 14384 2320 14564 2336
rect 14384 2262 14442 2320
rect 14498 2262 14564 2320
rect 14384 2242 14564 2262
rect 16448 2320 16628 2336
rect 16448 2262 16506 2320
rect 16562 2262 16628 2320
rect 16448 2242 16628 2262
rect 17390 1982 17450 3078
rect 2192 1886 2198 1938
rect 2250 1886 2260 1938
rect 2192 1882 2260 1886
rect 17362 1930 17488 1982
rect 17362 1876 17402 1930
rect 17454 1876 17488 1930
rect 17362 1828 17488 1876
rect 2538 1778 2718 1794
rect 2538 1720 2604 1778
rect 2660 1720 2718 1778
rect 2538 1700 2718 1720
rect 4534 1768 4714 1786
rect 4534 1710 4596 1768
rect 4652 1710 4714 1768
rect 4534 1692 4714 1710
rect 6486 1768 6666 1786
rect 6486 1710 6548 1768
rect 6604 1710 6666 1768
rect 6486 1692 6666 1710
rect 8488 1774 8668 1792
rect 8488 1716 8550 1774
rect 8606 1716 8668 1774
rect 8488 1698 8668 1716
rect 10440 1774 10620 1792
rect 10440 1716 10502 1774
rect 10558 1716 10620 1774
rect 10440 1698 10620 1716
rect 12432 1774 12612 1792
rect 12432 1716 12494 1774
rect 12550 1716 12612 1774
rect 12432 1698 12612 1716
rect 14384 1774 14564 1792
rect 14384 1716 14446 1774
rect 14502 1716 14564 1774
rect 14384 1698 14564 1716
rect 16448 1774 16628 1792
rect 16448 1716 16510 1774
rect 16566 1716 16628 1774
rect 16448 1698 16628 1716
<< via2 >>
rect 18768 43898 18962 44096
rect 18562 42762 18624 42820
rect 19124 42724 19186 42782
rect 18540 40890 18602 40948
rect 19106 40882 19168 40940
rect 18564 39262 18626 39320
rect 19106 39258 19168 39316
rect 18572 38066 18634 38124
rect 19122 38082 19184 38140
rect 18580 36996 18642 37054
rect 19128 36986 19190 37044
rect 18598 36200 18652 36256
rect 18652 36200 18656 36256
rect 19142 36228 19200 36284
rect 18374 34454 18454 34458
rect 18374 34376 18424 34454
rect 18424 34376 18454 34454
rect 18972 34376 19052 34458
rect 18382 32148 18462 32152
rect 18382 32070 18432 32148
rect 18432 32070 18462 32148
rect 18980 32070 19060 32152
rect 18390 29934 18470 29938
rect 18390 29856 18440 29934
rect 18440 29856 18470 29934
rect 18988 29856 19068 29938
rect 18372 27734 18452 27738
rect 18372 27656 18422 27734
rect 18422 27656 18452 27734
rect 18970 27656 19050 27738
rect 18380 25520 18460 25524
rect 18380 25442 18430 25520
rect 18430 25442 18460 25520
rect 18978 25442 19058 25524
rect 8536 23430 8618 23480
rect 8536 23400 8614 23430
rect 8614 23400 8618 23430
rect 10750 23438 10832 23488
rect 10750 23408 10828 23438
rect 10828 23408 10832 23438
rect 12950 23420 13032 23470
rect 12950 23390 13028 23420
rect 13028 23390 13032 23420
rect 15164 23428 15246 23478
rect 15164 23398 15242 23428
rect 15242 23398 15246 23428
rect 17470 23436 17552 23486
rect 17470 23406 17548 23436
rect 17548 23406 17552 23436
rect 8536 22802 8618 22882
rect 10750 22810 10832 22890
rect 12950 22792 13032 22872
rect 15164 22800 15246 22880
rect 17470 22808 17552 22888
rect 9540 17762 9600 17822
rect 15683 17612 15751 17674
rect 16455 17652 16523 17714
rect 17335 17652 17403 17714
rect 18121 17642 18189 17704
rect 19219 17646 19287 17708
rect 20099 17646 20167 17708
rect 20885 17636 20953 17698
rect 21475 17636 21543 17698
rect 22355 17636 22423 17698
rect 23141 17626 23209 17688
rect 4552 16570 4590 16614
rect 4590 16570 4608 16614
rect 4552 16558 4608 16570
rect 4976 16074 5034 16076
rect 4976 16020 5034 16074
rect 4746 15814 4808 15874
rect 9536 17218 9594 17278
rect 15691 17072 15759 17134
rect 16453 17110 16521 17172
rect 17343 17112 17411 17174
rect 18101 17104 18169 17166
rect 19217 17104 19285 17166
rect 20107 17106 20175 17168
rect 20865 17098 20933 17160
rect 21473 17094 21541 17156
rect 22363 17096 22431 17158
rect 23121 17088 23189 17150
rect 9418 16574 9456 16618
rect 9456 16574 9474 16618
rect 9418 16562 9474 16574
rect 9842 16078 9900 16080
rect 9842 16024 9900 16078
rect 9612 15818 9674 15878
rect 6712 15706 6780 15768
rect 4898 15270 4966 15332
rect 6130 15202 6198 15264
rect 9764 15274 9832 15336
rect 7114 15156 7182 15218
rect 4582 14986 4648 15052
rect 9448 14990 9514 15056
rect 5794 14654 5862 14716
rect 5012 14442 5078 14508
rect 4682 14244 4754 14314
rect 6350 14232 6418 14294
rect 7916 14222 7984 14284
rect 6828 13856 6896 13918
rect 4884 13700 4956 13770
rect 5862 13692 5930 13754
rect 7656 13676 7724 13738
rect 4576 13318 4648 13384
rect 5984 13390 6052 13450
rect 7136 13316 7204 13378
rect 5996 12856 6064 12916
rect 4990 12778 5062 12844
rect 4634 12576 4708 12642
rect 6280 12370 6348 12432
rect 4906 12034 4980 12100
rect 4560 11756 4640 11820
rect 6002 11830 6070 11892
rect 4994 11214 5074 11278
rect 4626 11010 4706 11074
rect 9878 14446 9944 14512
rect 9548 14248 9620 14318
rect 10660 14658 10728 14720
rect 16430 16660 16498 16722
rect 17188 16652 17256 16714
rect 18078 16654 18146 16716
rect 18686 16650 18754 16712
rect 19444 16642 19512 16704
rect 20334 16644 20402 16706
rect 21450 16644 21518 16706
rect 22208 16636 22276 16698
rect 23098 16638 23166 16700
rect 16410 16122 16478 16184
rect 17196 16112 17264 16174
rect 18076 16112 18144 16174
rect 18666 16112 18734 16174
rect 19452 16102 19520 16164
rect 20332 16102 20400 16164
rect 21430 16106 21498 16168
rect 22216 16096 22284 16158
rect 23096 16096 23164 16158
rect 11578 15710 11646 15772
rect 10996 15206 11064 15268
rect 11980 15160 12048 15222
rect 24400 14810 24462 14870
rect 9750 13704 9822 13774
rect 27000 14646 27122 14766
rect 11216 14236 11284 14298
rect 12782 14226 12850 14288
rect 11694 13860 11762 13922
rect 10728 13696 10796 13758
rect 9442 13322 9514 13388
rect 10850 13394 10918 13454
rect 12522 13680 12590 13742
rect 12002 13320 12070 13382
rect 10862 12860 10930 12920
rect 9856 12782 9928 12848
rect 9500 12580 9574 12646
rect 11146 12374 11214 12436
rect 9772 12038 9846 12104
rect 9426 11760 9506 11824
rect 10868 11834 10936 11896
rect 9860 11218 9940 11282
rect 9492 11014 9572 11078
rect 23992 14258 24054 14318
rect 4904 10476 4984 10540
rect 9770 10480 9850 10544
rect 6226 6580 6282 6638
rect 27550 14372 27682 14492
rect 6170 6030 6226 6088
rect 10774 5936 10832 6000
rect 12796 5928 12852 5986
rect 14754 5936 14810 5994
rect 16748 5942 16804 6000
rect 2564 5520 2620 5578
rect 4686 5512 4742 5570
rect 6638 5512 6694 5570
rect 8640 5518 8696 5576
rect 11214 5394 11270 5452
rect 12800 5382 12856 5440
rect 14758 5390 14814 5448
rect 16752 5396 16808 5454
rect 18726 5364 18784 5428
rect 10188 5062 10244 5120
rect 2584 4982 2640 5040
rect 4690 4966 4746 5024
rect 6642 4966 6698 5024
rect 8644 4972 8700 5030
rect 13032 5022 13088 5080
rect 15034 5016 15090 5074
rect 17056 4998 17112 5056
rect 18720 4816 18778 4880
rect 10788 4522 10844 4580
rect 13036 4476 13092 4534
rect 15038 4470 15094 4528
rect 17060 4452 17116 4510
rect 6194 3320 6254 3382
rect 6176 2766 6236 2828
rect 2604 2260 2660 2318
rect 4592 2256 4648 2314
rect 6544 2256 6600 2314
rect 8546 2262 8602 2320
rect 10498 2262 10554 2320
rect 12490 2262 12546 2320
rect 14442 2262 14498 2320
rect 16506 2262 16562 2320
rect 2604 1720 2656 1778
rect 2656 1720 2660 1778
rect 4596 1710 4652 1768
rect 6548 1710 6604 1768
rect 8550 1716 8606 1774
rect 10502 1716 10558 1774
rect 12494 1716 12550 1774
rect 14446 1716 14502 1774
rect 16510 1716 16566 1774
<< metal3 >>
rect 18590 44096 19128 44168
rect 18590 43898 18768 44096
rect 18962 43898 19128 44096
rect 18590 43828 19128 43898
rect 17652 43002 18076 43406
rect 17652 42820 18672 43002
rect 19448 42956 19880 43622
rect 17652 42762 18562 42820
rect 18624 42762 18672 42820
rect 17652 42578 18672 42762
rect 19102 42782 19880 42956
rect 19102 42724 19124 42782
rect 19186 42724 19880 42782
rect 17652 41110 18076 42578
rect 19102 42524 19880 42724
rect 18530 41110 18620 41118
rect 17652 40948 18636 41110
rect 19448 41102 19880 42524
rect 19116 41096 19880 41102
rect 17652 40890 18540 40948
rect 18602 40890 18636 40948
rect 17652 40686 18636 40890
rect 19090 40940 19880 41096
rect 19090 40882 19106 40940
rect 19168 40882 19880 40940
rect 17652 39508 18076 40686
rect 19090 40670 19880 40882
rect 17652 39320 18636 39508
rect 19448 39486 19880 40670
rect 19116 39484 19880 39486
rect 17652 39262 18564 39320
rect 18626 39262 18636 39320
rect 17652 39084 18636 39262
rect 19092 39316 19880 39484
rect 19092 39258 19106 39316
rect 19168 39258 19880 39316
rect 17652 38286 18076 39084
rect 19092 39058 19880 39258
rect 19116 39054 19880 39058
rect 19448 38310 19880 39054
rect 18558 38286 18648 38298
rect 17652 38124 18658 38286
rect 17652 38066 18572 38124
rect 18634 38066 18658 38124
rect 17652 37862 18658 38066
rect 19094 38140 19880 38310
rect 19094 38082 19122 38140
rect 19184 38082 19880 38140
rect 19094 37878 19880 38082
rect 17652 37228 18076 37862
rect 17652 37054 18656 37228
rect 19448 37222 19880 37878
rect 17652 36996 18580 37054
rect 18642 36996 18656 37054
rect 17652 36804 18656 36996
rect 19116 37044 19880 37222
rect 19116 36986 19128 37044
rect 19190 36986 19880 37044
rect 17652 36446 18076 36804
rect 19116 36790 19880 36986
rect 19448 36448 19880 36790
rect 17652 36256 18674 36446
rect 17652 36200 18598 36256
rect 18656 36200 18674 36256
rect 17652 36022 18674 36200
rect 19120 36284 19880 36448
rect 19120 36228 19142 36284
rect 19200 36228 19880 36284
rect 17652 34644 18076 36022
rect 19120 36016 19880 36228
rect 17652 34458 18512 34644
rect 19448 34628 19880 36016
rect 17652 34376 18374 34458
rect 18454 34376 18512 34458
rect 17652 34220 18512 34376
rect 18960 34458 19880 34628
rect 18960 34376 18972 34458
rect 19052 34376 19880 34458
rect 17652 33912 17888 34220
rect 18960 34204 19880 34376
rect 17652 32338 18076 33912
rect 17652 32152 18520 32338
rect 19448 32322 19880 34204
rect 17652 32070 18382 32152
rect 18462 32070 18520 32152
rect 17652 31914 18520 32070
rect 18968 32152 19880 32322
rect 18968 32070 18980 32152
rect 19060 32070 19880 32152
rect 17652 31698 17888 31914
rect 18968 31898 19880 32070
rect 17652 30124 18076 31698
rect 17652 29938 18528 30124
rect 19448 30108 19880 31898
rect 17652 29856 18390 29938
rect 18470 29856 18528 29938
rect 17652 29700 18528 29856
rect 18976 29938 19880 30108
rect 18976 29856 18988 29938
rect 19068 29856 19880 29938
rect 17652 29498 17888 29700
rect 18976 29684 19880 29856
rect 17652 27924 18076 29498
rect 17652 27738 18510 27924
rect 19448 27908 19880 29684
rect 17652 27656 18372 27738
rect 18452 27656 18510 27738
rect 17652 27500 18510 27656
rect 18958 27738 19880 27908
rect 18958 27656 18970 27738
rect 19050 27656 19880 27738
rect 17652 27284 17888 27500
rect 18958 27484 19880 27656
rect 17652 25710 18076 27284
rect 17652 25524 18518 25710
rect 19448 25694 19880 27484
rect 17652 25442 18380 25524
rect 18460 25442 18518 25524
rect 17652 25286 18518 25442
rect 18966 25524 19880 25694
rect 18966 25442 18978 25524
rect 19058 25442 19880 25524
rect 17652 24978 17888 25286
rect 18966 25270 19880 25442
rect 17652 24396 18076 24978
rect 228 24272 18076 24396
rect 228 24092 300 24272
rect 488 24092 18076 24272
rect 228 23972 18076 24092
rect 8380 23480 8804 23972
rect 8380 23400 8536 23480
rect 8618 23400 8804 23480
rect 8380 23342 8804 23400
rect 10594 23488 11018 23972
rect 10594 23408 10750 23488
rect 10832 23408 11018 23488
rect 10594 23350 11018 23408
rect 12794 23470 13218 23972
rect 12794 23390 12950 23470
rect 13032 23390 13218 23470
rect 12794 23332 13218 23390
rect 15008 23478 15432 23972
rect 15008 23398 15164 23478
rect 15246 23398 15432 23478
rect 15008 23340 15432 23398
rect 17314 23486 17738 23972
rect 17314 23406 17470 23486
rect 17552 23406 17738 23486
rect 17314 23348 17738 23406
rect 8364 22882 8788 22894
rect 8364 22802 8536 22882
rect 8618 22802 8788 22882
rect 8364 22244 8788 22802
rect 10578 22890 11002 22902
rect 10578 22810 10750 22890
rect 10832 22810 11002 22890
rect 10578 22244 11002 22810
rect 12778 22872 13202 22884
rect 12778 22792 12950 22872
rect 13032 22792 13202 22872
rect 12778 22244 13202 22792
rect 14992 22880 15416 22892
rect 14992 22800 15164 22880
rect 15246 22800 15416 22880
rect 14992 22244 15416 22800
rect 17298 22888 17722 22900
rect 17298 22808 17470 22888
rect 17552 22808 17722 22888
rect 17298 22252 17722 22808
rect 19448 22252 19880 25270
rect 16310 22244 19880 22252
rect 898 22150 19880 22244
rect 898 21970 978 22150
rect 1166 21970 19880 22150
rect 898 21820 19880 21970
rect 814 17848 23871 17936
rect 814 17780 996 17848
rect 1066 17822 23871 17848
rect 1066 17780 9540 17822
rect 814 17762 9540 17780
rect 9600 17762 23871 17822
rect 814 17722 23871 17762
rect 15360 17674 15904 17722
rect 16084 17718 23871 17722
rect 15360 17646 15683 17674
rect 15606 17612 15683 17646
rect 15751 17646 15904 17674
rect 16392 17714 16606 17718
rect 16392 17652 16455 17714
rect 16523 17652 16606 17714
rect 15751 17612 15820 17646
rect 16392 17635 16606 17652
rect 17258 17714 17472 17718
rect 17258 17652 17335 17714
rect 17403 17652 17472 17714
rect 17258 17641 17472 17652
rect 18052 17704 18266 17718
rect 18052 17642 18121 17704
rect 18189 17642 18266 17704
rect 18052 17627 18266 17642
rect 19156 17708 19370 17718
rect 19156 17646 19219 17708
rect 19287 17646 19370 17708
rect 19156 17629 19370 17646
rect 20022 17708 20236 17718
rect 20022 17646 20099 17708
rect 20167 17646 20236 17708
rect 20022 17635 20236 17646
rect 20816 17698 21030 17718
rect 20816 17636 20885 17698
rect 20953 17636 21030 17698
rect 20816 17621 21030 17636
rect 21412 17698 21626 17718
rect 21412 17636 21475 17698
rect 21543 17636 21626 17698
rect 21412 17619 21626 17636
rect 22278 17698 22492 17718
rect 22278 17636 22355 17698
rect 22423 17636 22492 17698
rect 22278 17625 22492 17636
rect 23072 17688 23286 17718
rect 23072 17626 23141 17688
rect 23209 17626 23286 17688
rect 15606 17601 15820 17612
rect 23072 17611 23286 17626
rect 200 17278 13306 17330
rect 200 17218 9536 17278
rect 9594 17218 13306 17278
rect 200 17104 13306 17218
rect 16373 17172 16601 17188
rect 200 16942 322 17104
rect 474 17038 13306 17104
rect 15611 17134 15839 17144
rect 15611 17072 15691 17134
rect 15759 17072 15839 17134
rect 16373 17110 16453 17172
rect 16521 17110 16601 17172
rect 16373 17074 16601 17110
rect 17263 17174 17491 17184
rect 17263 17112 17343 17174
rect 17411 17112 17491 17174
rect 17263 17074 17491 17112
rect 18031 17166 18259 17174
rect 18031 17104 18101 17166
rect 18169 17104 18259 17166
rect 18031 17074 18259 17104
rect 19137 17166 19365 17182
rect 19137 17104 19217 17166
rect 19285 17104 19365 17166
rect 19137 17074 19365 17104
rect 20027 17168 20255 17178
rect 20027 17106 20107 17168
rect 20175 17106 20255 17168
rect 20027 17074 20255 17106
rect 20795 17160 21023 17168
rect 20795 17098 20865 17160
rect 20933 17098 21023 17160
rect 20795 17074 21023 17098
rect 21393 17156 21621 17172
rect 21393 17094 21473 17156
rect 21541 17094 21621 17156
rect 21393 17074 21621 17094
rect 22283 17158 22511 17168
rect 22283 17096 22363 17158
rect 22431 17096 22511 17158
rect 22283 17074 22511 17096
rect 23051 17150 23279 17158
rect 23051 17088 23121 17150
rect 23189 17088 23279 17150
rect 23051 17074 23279 17088
rect 15611 17038 15839 17072
rect 16134 17038 23388 17074
rect 474 16942 23388 17038
rect 200 16810 23388 16942
rect 200 16808 13306 16810
rect 4036 16628 4280 16808
rect 4036 16614 4844 16628
rect 4036 16558 4552 16614
rect 4608 16558 4844 16614
rect 4036 16536 4844 16558
rect 4036 15884 4280 16536
rect 4880 16076 5584 16082
rect 4880 16020 4976 16076
rect 5034 16020 5584 16076
rect 4880 15994 5584 16020
rect 5342 15912 5584 15994
rect 4036 15874 4938 15884
rect 4036 15814 4746 15874
rect 4808 15814 4938 15874
rect 4036 15792 4938 15814
rect 4036 15066 4280 15792
rect 5340 15344 5584 15912
rect 4834 15332 5584 15344
rect 4834 15270 4898 15332
rect 4966 15270 5584 15332
rect 6320 15780 6502 16808
rect 6320 15768 6896 15780
rect 6320 15706 6712 15768
rect 6780 15706 6896 15768
rect 6320 15684 6896 15706
rect 6320 15278 6502 15684
rect 4834 15256 5584 15270
rect 4036 15052 4900 15066
rect 4036 14986 4582 15052
rect 4648 14986 4900 15052
rect 4036 14974 4900 14986
rect 4036 14324 4280 14974
rect 5340 14738 5584 15256
rect 6088 15264 6502 15278
rect 6088 15202 6130 15264
rect 6198 15202 6502 15264
rect 6088 15180 6502 15202
rect 5340 14716 6026 14738
rect 5340 14654 5794 14716
rect 5862 14654 6026 14716
rect 5340 14642 6026 14654
rect 5340 14522 5584 14642
rect 4942 14508 5584 14522
rect 4942 14442 5012 14508
rect 5078 14442 5584 14508
rect 4942 14434 5584 14442
rect 4036 14314 4880 14324
rect 4036 14244 4682 14314
rect 4754 14244 4880 14314
rect 4036 14232 4880 14244
rect 4036 13404 4280 14232
rect 5340 13776 5584 14434
rect 6320 14433 6502 15180
rect 7050 15218 7552 15236
rect 7050 15156 7114 15218
rect 7182 15156 7552 15218
rect 7050 15140 7552 15156
rect 6321 14430 6502 14433
rect 6321 14334 6684 14430
rect 6321 14328 6502 14334
rect 6320 14294 6502 14328
rect 6320 14232 6350 14294
rect 6418 14232 6502 14294
rect 6320 14213 6502 14232
rect 6589 13938 6684 14334
rect 6584 13918 6948 13938
rect 6584 13856 6828 13918
rect 6896 13856 6948 13918
rect 6584 13846 6948 13856
rect 4822 13772 5584 13776
rect 4822 13770 6086 13772
rect 4822 13700 4884 13770
rect 4956 13754 6086 13770
rect 4956 13700 5862 13754
rect 4822 13692 5862 13700
rect 5930 13692 6086 13754
rect 4822 13688 6086 13692
rect 5340 13676 6086 13688
rect 4036 13384 4884 13404
rect 4036 13318 4576 13384
rect 4648 13318 4884 13384
rect 4036 13312 4884 13318
rect 4036 12658 4280 13312
rect 5340 12928 5584 13676
rect 6589 13470 6684 13846
rect 5948 13450 6684 13470
rect 5948 13390 5984 13450
rect 6052 13390 6684 13450
rect 7348 13752 7552 15140
rect 7838 14284 8072 16808
rect 7838 14222 7916 14284
rect 7984 14222 8072 14284
rect 7838 14188 8072 14222
rect 8902 16792 9242 16808
rect 11186 16792 11464 16808
rect 12704 16792 13034 16808
rect 8902 16632 9146 16792
rect 8902 16618 9710 16632
rect 8902 16562 9418 16618
rect 9474 16562 9710 16618
rect 8902 16540 9710 16562
rect 8902 15888 9146 16540
rect 9746 16080 10450 16086
rect 9746 16024 9842 16080
rect 9900 16024 10450 16080
rect 9746 15998 10450 16024
rect 10208 15916 10450 15998
rect 8902 15878 9804 15888
rect 8902 15818 9612 15878
rect 9674 15818 9804 15878
rect 8902 15796 9804 15818
rect 8902 15070 9146 15796
rect 10206 15348 10450 15916
rect 9700 15336 10450 15348
rect 9700 15274 9764 15336
rect 9832 15274 10450 15336
rect 11186 15784 11368 16792
rect 11186 15772 11762 15784
rect 11186 15710 11578 15772
rect 11646 15710 11762 15772
rect 11186 15688 11762 15710
rect 11186 15282 11368 15688
rect 9700 15260 10450 15274
rect 8902 15056 9766 15070
rect 8902 14990 9448 15056
rect 9514 14990 9766 15056
rect 8902 14978 9766 14990
rect 8902 14328 9146 14978
rect 10206 14742 10450 15260
rect 10954 15268 11368 15282
rect 10954 15206 10996 15268
rect 11064 15206 11368 15268
rect 10954 15184 11368 15206
rect 10206 14720 10892 14742
rect 10206 14658 10660 14720
rect 10728 14658 10892 14720
rect 10206 14646 10892 14658
rect 10206 14526 10450 14646
rect 9808 14512 10450 14526
rect 9808 14446 9878 14512
rect 9944 14446 10450 14512
rect 9808 14438 10450 14446
rect 8902 14318 9746 14328
rect 8902 14248 9548 14318
rect 9620 14248 9746 14318
rect 8902 14236 9746 14248
rect 7348 13738 7746 13752
rect 7348 13676 7656 13738
rect 7724 13676 7746 13738
rect 7348 13656 7746 13676
rect 7348 13394 7552 13656
rect 5948 13378 6684 13390
rect 5340 12916 6098 12928
rect 5340 12856 5996 12916
rect 6064 12856 6098 12916
rect 5340 12854 6098 12856
rect 4926 12844 6098 12854
rect 4926 12778 4990 12844
rect 5062 12832 6098 12844
rect 5062 12778 5584 12832
rect 4926 12766 5584 12778
rect 4036 12642 4952 12658
rect 4036 12576 4634 12642
rect 4708 12576 4952 12642
rect 4036 12566 4952 12576
rect 4036 11840 4280 12566
rect 5340 12110 5584 12766
rect 6589 12454 6684 13378
rect 7092 13378 7552 13394
rect 7092 13316 7136 13378
rect 7204 13316 7552 13378
rect 7092 13298 7552 13316
rect 6193 12432 6684 12454
rect 6193 12370 6280 12432
rect 6348 12370 6684 12432
rect 6193 12359 6684 12370
rect 4850 12100 5584 12110
rect 4850 12034 4906 12100
rect 4980 12034 5584 12100
rect 4850 12022 5584 12034
rect 5340 11906 5584 12022
rect 5340 11892 6100 11906
rect 4036 11820 4838 11840
rect 4036 11756 4560 11820
rect 4640 11756 4838 11820
rect 4036 11748 4838 11756
rect 5340 11830 6002 11892
rect 6070 11830 6100 11892
rect 5340 11810 6100 11830
rect 4036 11090 4280 11748
rect 5340 11294 5584 11810
rect 4936 11278 5584 11294
rect 4936 11214 4994 11278
rect 5074 11214 5584 11278
rect 4936 11200 5584 11214
rect 4036 11074 4904 11090
rect 4036 11010 4626 11074
rect 4706 11010 4904 11074
rect 4036 10998 4904 11010
rect 4036 10996 4280 10998
rect 5340 10554 5584 11200
rect 4852 10540 5584 10554
rect 4852 10476 4904 10540
rect 4984 10476 5584 10540
rect 4852 10448 5584 10476
rect 5340 9882 5584 10448
rect 7348 9882 7552 13298
rect 8902 13408 9146 14236
rect 10206 13780 10450 14438
rect 11186 14437 11368 15184
rect 11916 15222 12418 15240
rect 11916 15160 11980 15222
rect 12048 15160 12418 15222
rect 11916 15144 12418 15160
rect 11187 14434 11368 14437
rect 11187 14338 11550 14434
rect 11187 14332 11368 14338
rect 11186 14298 11368 14332
rect 11186 14236 11216 14298
rect 11284 14236 11368 14298
rect 11186 14217 11368 14236
rect 11455 13942 11550 14338
rect 11450 13922 11814 13942
rect 11450 13860 11694 13922
rect 11762 13860 11814 13922
rect 11450 13850 11814 13860
rect 9688 13776 10450 13780
rect 9688 13774 10952 13776
rect 9688 13704 9750 13774
rect 9822 13758 10952 13774
rect 9822 13704 10728 13758
rect 9688 13696 10728 13704
rect 10796 13696 10952 13758
rect 9688 13692 10952 13696
rect 10206 13680 10952 13692
rect 8902 13388 9750 13408
rect 8902 13322 9442 13388
rect 9514 13322 9750 13388
rect 8902 13316 9750 13322
rect 8902 12662 9146 13316
rect 10206 12932 10450 13680
rect 11455 13474 11550 13850
rect 10814 13454 11550 13474
rect 10814 13394 10850 13454
rect 10918 13394 11550 13454
rect 12214 13756 12418 15144
rect 12704 14288 12938 16792
rect 15198 15406 15426 16810
rect 16134 16794 23388 16810
rect 16340 16722 16568 16794
rect 16340 16660 16430 16722
rect 16498 16660 16568 16722
rect 16340 16652 16568 16660
rect 17108 16714 17336 16794
rect 17108 16652 17188 16714
rect 17256 16652 17336 16714
rect 17108 16642 17336 16652
rect 17998 16716 18226 16794
rect 17998 16654 18078 16716
rect 18146 16654 18226 16716
rect 17998 16638 18226 16654
rect 18596 16712 18824 16794
rect 18596 16650 18686 16712
rect 18754 16650 18824 16712
rect 18596 16642 18824 16650
rect 19364 16704 19592 16794
rect 19364 16642 19444 16704
rect 19512 16642 19592 16704
rect 19364 16632 19592 16642
rect 20254 16706 20482 16794
rect 20254 16644 20334 16706
rect 20402 16644 20482 16706
rect 20254 16628 20482 16644
rect 21360 16706 21588 16794
rect 21360 16644 21450 16706
rect 21518 16644 21588 16706
rect 21360 16636 21588 16644
rect 22128 16698 22356 16794
rect 22128 16636 22208 16698
rect 22276 16636 22356 16698
rect 22128 16626 22356 16636
rect 23018 16700 23246 16794
rect 23018 16638 23098 16700
rect 23166 16638 23246 16700
rect 23018 16622 23246 16638
rect 16333 16184 16547 16199
rect 16333 16122 16410 16184
rect 16478 16122 16547 16184
rect 16333 16027 16547 16122
rect 17127 16174 17341 16185
rect 17127 16112 17196 16174
rect 17264 16112 17341 16174
rect 17127 16027 17341 16112
rect 17993 16174 18207 16191
rect 17993 16112 18076 16174
rect 18144 16112 18207 16174
rect 17993 16027 18207 16112
rect 18589 16174 18803 16189
rect 18589 16112 18666 16174
rect 18734 16112 18803 16174
rect 16197 16018 18300 16027
rect 16197 16017 18510 16018
rect 18589 16017 18803 16112
rect 19383 16164 19597 16175
rect 19383 16102 19452 16164
rect 19520 16102 19597 16164
rect 19383 16017 19597 16102
rect 20249 16164 20463 16181
rect 20249 16102 20332 16164
rect 20400 16102 20463 16164
rect 20249 16017 20463 16102
rect 21353 16168 21567 16183
rect 21353 16106 21430 16168
rect 21498 16106 21567 16168
rect 21353 16017 21567 16106
rect 16197 16011 21567 16017
rect 22147 16158 22361 16169
rect 22147 16096 22216 16158
rect 22284 16096 22361 16158
rect 22147 16011 22361 16096
rect 23013 16158 23227 16175
rect 23013 16096 23096 16158
rect 23164 16096 23227 16158
rect 23013 16027 23227 16096
rect 23657 16027 23871 17718
rect 22627 16011 23871 16027
rect 16197 16010 21710 16011
rect 21790 16010 21966 16011
rect 16197 16006 21966 16010
rect 22094 16006 23871 16011
rect 16197 15896 23871 16006
rect 16197 15813 23874 15896
rect 18292 15803 23874 15813
rect 20597 15797 23874 15803
rect 23270 15794 23874 15797
rect 15198 15178 24536 15406
rect 24310 15150 24536 15178
rect 24310 14870 24538 15150
rect 24310 14810 24400 14870
rect 24462 14810 24538 14870
rect 24310 14790 24538 14810
rect 26956 14766 27174 14788
rect 26956 14646 27000 14766
rect 27122 14646 27174 14766
rect 26956 14604 27174 14646
rect 27512 14492 27730 14510
rect 27512 14372 27550 14492
rect 27682 14372 27730 14492
rect 27512 14336 27730 14372
rect 12704 14226 12782 14288
rect 12850 14226 12938 14288
rect 12704 14192 12938 14226
rect 23852 14318 24212 14334
rect 23852 14258 23992 14318
rect 24054 14258 24212 14318
rect 23852 14128 24212 14258
rect 23852 13946 24204 14128
rect 12214 13742 12612 13756
rect 12214 13680 12522 13742
rect 12590 13680 12612 13742
rect 12214 13660 12612 13680
rect 15110 13726 24204 13946
rect 12214 13398 12418 13660
rect 10814 13382 11550 13394
rect 10206 12920 10964 12932
rect 10206 12860 10862 12920
rect 10930 12860 10964 12920
rect 10206 12858 10964 12860
rect 9792 12848 10964 12858
rect 9792 12782 9856 12848
rect 9928 12836 10964 12848
rect 9928 12782 10450 12836
rect 9792 12770 10450 12782
rect 8902 12646 9818 12662
rect 8902 12580 9500 12646
rect 9574 12580 9818 12646
rect 8902 12570 9818 12580
rect 8902 11844 9146 12570
rect 10206 12114 10450 12770
rect 11455 12458 11550 13382
rect 11958 13382 12418 13398
rect 11958 13320 12002 13382
rect 12070 13320 12418 13382
rect 11958 13302 12418 13320
rect 11059 12436 11550 12458
rect 11059 12374 11146 12436
rect 11214 12374 11550 12436
rect 11059 12363 11550 12374
rect 9716 12104 10450 12114
rect 9716 12038 9772 12104
rect 9846 12038 10450 12104
rect 9716 12026 10450 12038
rect 10206 11910 10450 12026
rect 10206 11896 10966 11910
rect 8902 11824 9704 11844
rect 8902 11760 9426 11824
rect 9506 11760 9704 11824
rect 8902 11752 9704 11760
rect 10206 11834 10868 11896
rect 10936 11834 10966 11896
rect 10206 11814 10966 11834
rect 8902 11094 9146 11752
rect 10206 11298 10450 11814
rect 9802 11282 10450 11298
rect 9802 11218 9860 11282
rect 9940 11218 10450 11282
rect 9802 11204 10450 11218
rect 8902 11078 9770 11094
rect 8902 11014 9492 11078
rect 9572 11014 9770 11078
rect 8902 11002 9770 11014
rect 8902 11000 9146 11002
rect 10206 10558 10450 11204
rect 9718 10544 10450 10558
rect 9718 10480 9770 10544
rect 9850 10480 10450 10544
rect 9718 10452 10450 10480
rect 10206 9944 10450 10452
rect 12214 9944 12418 13302
rect 15110 13586 24208 13726
rect 10206 9922 10540 9944
rect 12214 9922 12508 9944
rect 13258 9922 13626 9926
rect 8392 9890 14696 9922
rect 15110 9890 15470 13586
rect 8392 9886 15470 9890
rect 8312 9882 15470 9886
rect 800 9724 15470 9882
rect 800 9562 994 9724
rect 1146 9562 15470 9724
rect 800 9530 15470 9562
rect 800 9376 13253 9530
rect 6108 6638 6646 6736
rect 6108 6580 6226 6638
rect 6282 6580 6646 6638
rect 6108 6556 6646 6580
rect 372 6088 6274 6108
rect 372 6074 6170 6088
rect 372 5986 392 6074
rect 498 6030 6170 6074
rect 6226 6030 6274 6088
rect 498 5986 6274 6030
rect 372 5954 6274 5986
rect 6466 5814 6646 6556
rect 9652 6050 18838 6222
rect 9652 6042 11818 6050
rect 9652 5814 9832 6042
rect 802 5774 9844 5814
rect 802 5670 936 5774
rect 1052 5670 9844 5774
rect 802 5634 9844 5670
rect 2512 5578 2692 5634
rect 4378 5620 4558 5634
rect 2512 5520 2564 5578
rect 2620 5520 2692 5578
rect 2512 5506 2692 5520
rect 4628 5574 4808 5634
rect 6104 5620 6284 5634
rect 6572 5602 6766 5634
rect 8010 5620 8190 5634
rect 6572 5574 6762 5602
rect 4628 5570 4810 5574
rect 4628 5512 4686 5570
rect 4742 5512 4810 5570
rect 4628 5492 4810 5512
rect 6570 5570 6762 5574
rect 6570 5512 6638 5570
rect 6694 5512 6762 5570
rect 6570 5492 6762 5512
rect 8584 5576 8762 5634
rect 8584 5518 8640 5576
rect 8696 5574 8762 5576
rect 8696 5518 8764 5574
rect 8584 5498 8764 5518
rect 4628 5478 4808 5492
rect 6570 5488 6750 5492
rect 10128 5120 10308 6042
rect 10708 6000 10888 6042
rect 10708 5936 10774 6000
rect 10832 5936 10888 6000
rect 10708 5924 10888 5936
rect 12736 5986 12922 6050
rect 12736 5928 12796 5986
rect 12852 5928 12922 5986
rect 12736 5922 12922 5928
rect 12740 5908 12920 5922
rect 10972 5452 12936 5480
rect 10972 5394 11214 5452
rect 11270 5440 12936 5452
rect 11270 5394 12800 5440
rect 10972 5382 12800 5394
rect 12856 5382 12936 5440
rect 10972 5300 12936 5382
rect 10128 5062 10188 5120
rect 10244 5062 10308 5120
rect 2520 5040 2700 5048
rect 2520 4982 2584 5040
rect 2640 4982 2700 5040
rect 2520 4850 2700 4982
rect 4628 5024 4808 5048
rect 4628 4966 4690 5024
rect 4746 4966 4808 5024
rect 4380 4850 4560 4858
rect 4628 4850 4808 4966
rect 6580 5024 6760 5048
rect 6580 4966 6642 5024
rect 6698 4966 6760 5024
rect 6580 4948 6760 4966
rect 6092 4850 6272 4858
rect 6574 4850 6760 4948
rect 8582 5030 8762 5054
rect 10128 5046 10308 5062
rect 8582 4972 8644 5030
rect 8700 4972 8762 5030
rect 8002 4852 8182 4858
rect 8582 4852 8762 4972
rect 7674 4850 9835 4852
rect 198 4814 9835 4850
rect 198 4710 330 4814
rect 446 4710 9835 4814
rect 198 4670 9835 4710
rect 9652 4496 9832 4670
rect 10732 4580 10912 4598
rect 10732 4522 10788 4580
rect 10844 4522 10912 4580
rect 9652 4376 9834 4496
rect 10732 4376 10912 4522
rect 11576 4376 11756 5300
rect 13626 5174 13798 6050
rect 14696 5994 14882 6050
rect 14696 5952 14754 5994
rect 14698 5936 14754 5952
rect 14810 5952 14882 5994
rect 16690 6000 16876 6050
rect 17510 6042 18838 6050
rect 16690 5958 16748 6000
rect 14810 5936 14878 5952
rect 14698 5916 14878 5936
rect 16692 5942 16748 5958
rect 16804 5958 16876 6000
rect 16804 5942 16872 5958
rect 16692 5922 16872 5942
rect 14688 5454 16890 5480
rect 14688 5448 16752 5454
rect 14688 5390 14758 5448
rect 14814 5396 16752 5448
rect 16808 5396 16890 5454
rect 14814 5390 16890 5396
rect 14688 5308 16890 5390
rect 12976 5124 15154 5174
rect 12976 5080 15156 5124
rect 12976 5022 13032 5080
rect 13088 5074 15156 5080
rect 13088 5022 15034 5074
rect 12976 5016 15034 5022
rect 15090 5072 15156 5074
rect 15090 5016 15158 5072
rect 12976 5002 15158 5016
rect 14978 4996 15158 5002
rect 12974 4534 13154 4558
rect 12974 4476 13036 4534
rect 13092 4476 13154 4534
rect 9652 4368 11818 4376
rect 12974 4368 13154 4476
rect 14976 4528 15156 4552
rect 14976 4470 15038 4528
rect 15094 4470 15156 4528
rect 14976 4368 15156 4470
rect 15878 4368 16050 5308
rect 17648 5168 17828 6042
rect 18658 5428 18838 6042
rect 18658 5364 18726 5428
rect 18784 5364 18838 5428
rect 18658 5354 18838 5364
rect 17002 5106 17828 5168
rect 17000 5056 17828 5106
rect 17000 4998 17056 5056
rect 17112 4998 17828 5056
rect 17000 4988 17828 4998
rect 17000 4978 17180 4988
rect 18662 4880 18842 4888
rect 18662 4816 18720 4880
rect 18778 4816 18842 4880
rect 9652 4352 16050 4368
rect 16998 4510 17178 4534
rect 16998 4452 17060 4510
rect 17116 4452 17178 4510
rect 16998 4368 17178 4452
rect 18662 4376 18842 4816
rect 17510 4368 18840 4376
rect 16998 4352 18840 4368
rect 9652 4328 18840 4352
rect 9656 4196 18840 4328
rect 6082 3382 6656 3408
rect 6082 3320 6194 3382
rect 6254 3320 6656 3382
rect 6082 3228 6656 3320
rect 294 2828 6298 2858
rect 294 2808 6176 2828
rect 294 2714 384 2808
rect 484 2766 6176 2808
rect 6236 2766 6298 2828
rect 484 2714 6298 2766
rect 294 2664 6298 2714
rect 6476 2554 6656 3228
rect 794 2518 16633 2554
rect 794 2410 936 2518
rect 1068 2410 16633 2518
rect 794 2380 16633 2410
rect 794 2374 3426 2380
rect 3626 2374 5476 2380
rect 5676 2376 16633 2380
rect 2540 2318 2720 2374
rect 2540 2260 2604 2318
rect 2660 2260 2720 2318
rect 2540 2244 2720 2260
rect 4536 2314 4716 2374
rect 4536 2256 4592 2314
rect 4648 2256 4716 2314
rect 4536 2236 4716 2256
rect 6476 2314 6668 2376
rect 6476 2256 6544 2314
rect 6600 2256 6668 2314
rect 6476 2236 6668 2256
rect 8490 2320 8670 2376
rect 8490 2262 8546 2320
rect 8602 2262 8670 2320
rect 8490 2242 8670 2262
rect 10430 2320 10622 2376
rect 10430 2262 10498 2320
rect 10554 2262 10622 2320
rect 10430 2242 10622 2262
rect 12434 2320 12614 2376
rect 12434 2262 12490 2320
rect 12546 2262 12614 2320
rect 12434 2242 12614 2262
rect 14374 2320 14566 2376
rect 14374 2262 14442 2320
rect 14498 2262 14566 2320
rect 14374 2242 14566 2262
rect 16438 2320 16630 2376
rect 16438 2262 16506 2320
rect 16562 2262 16630 2320
rect 16438 2242 16630 2262
rect 10430 2238 10610 2242
rect 14374 2238 14554 2242
rect 16438 2238 16618 2242
rect 6476 2232 6656 2236
rect 2542 1778 2722 1790
rect 2542 1720 2604 1778
rect 2660 1720 2722 1778
rect 2542 1590 2722 1720
rect 4534 1768 4714 1792
rect 4534 1710 4596 1768
rect 4652 1710 4714 1768
rect 4534 1590 4714 1710
rect 6486 1768 6666 1792
rect 6486 1710 6548 1768
rect 6604 1710 6666 1768
rect 6486 1692 6666 1710
rect 6480 1590 6666 1692
rect 8488 1774 8668 1798
rect 8488 1716 8550 1774
rect 8606 1716 8668 1774
rect 8488 1596 8668 1716
rect 10440 1774 10620 1798
rect 10440 1716 10502 1774
rect 10558 1716 10620 1774
rect 10440 1698 10620 1716
rect 10434 1596 10620 1698
rect 12432 1774 12612 1798
rect 12432 1716 12494 1774
rect 12550 1716 12612 1774
rect 12432 1596 12612 1716
rect 14384 1774 14564 1798
rect 14384 1716 14446 1774
rect 14502 1716 14564 1774
rect 16448 1774 16628 1798
rect 16448 1716 16510 1774
rect 16566 1716 16628 1774
rect 14384 1698 14564 1716
rect 14378 1596 14564 1698
rect 16442 1686 16628 1716
rect 16442 1656 16626 1686
rect 7580 1592 9430 1596
rect 9630 1592 11402 1596
rect 11524 1592 13374 1596
rect 13574 1592 15346 1596
rect 7456 1590 15346 1592
rect 210 1586 3426 1590
rect 3626 1586 5476 1590
rect 5676 1588 15630 1590
rect 16446 1588 16626 1656
rect 5676 1586 16626 1588
rect 210 1548 16626 1586
rect 210 1438 336 1548
rect 456 1438 16626 1548
rect 210 1410 16626 1438
<< via3 >>
rect 18768 43898 18962 44096
rect 300 24092 488 24272
rect 978 21970 1166 22150
rect 996 17780 1066 17848
rect 322 16942 474 17104
rect 27000 14646 27122 14766
rect 27550 14372 27682 14492
rect 994 9562 1146 9724
rect 392 5986 498 6074
rect 936 5670 1052 5774
rect 330 4710 446 4814
rect 384 2714 484 2808
rect 936 2410 1068 2518
rect 336 1438 456 1548
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44168 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 200 24272 600 44152
rect 200 24092 300 24272
rect 488 24092 600 24272
rect 200 17104 600 24092
rect 200 16942 322 17104
rect 474 16942 600 17104
rect 200 6074 600 16942
rect 200 5986 392 6074
rect 498 5986 600 6074
rect 200 4814 600 5986
rect 200 4710 330 4814
rect 446 4710 600 4814
rect 200 2808 600 4710
rect 200 2714 384 2808
rect 484 2714 600 2808
rect 200 1548 600 2714
rect 200 1438 336 1548
rect 456 1438 600 1548
rect 200 1000 600 1438
rect 800 22150 1200 44152
rect 18590 44096 19130 44168
rect 18590 43898 18768 44096
rect 18962 43898 19130 44096
rect 18590 43830 19130 43898
rect 800 21970 978 22150
rect 1166 21970 1200 22150
rect 800 17848 1200 21970
rect 800 17780 996 17848
rect 1066 17780 1200 17848
rect 800 9724 1200 17780
rect 27110 14788 27170 45152
rect 26956 14766 27174 14788
rect 26956 14646 27000 14766
rect 27122 14646 27174 14766
rect 26956 14604 27174 14646
rect 27662 14510 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 27512 14492 27730 14510
rect 27512 14372 27550 14492
rect 27682 14372 27730 14492
rect 27512 14336 27730 14372
rect 800 9562 994 9724
rect 1146 9562 1200 9724
rect 800 5774 1200 9562
rect 800 5670 936 5774
rect 1052 5670 1200 5774
rect 800 2518 1200 5670
rect 800 2410 936 2518
rect 1068 2410 1200 2518
rect 800 1000 1200 2410
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 0 30542 196
use CLA  CLA_0
timestamp 1755018483
transform 1 0 4568 0 1 15292
box -138 -4838 3744 1342
use CLA  CLA_1
timestamp 1755018483
transform 1 0 9434 0 1 15296
box -138 -4838 3744 1342
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 9760 0 1 22852
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_1
timestamp 1723858470
transform 1 0 11960 0 1 22834
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_2
timestamp 1723858470
transform 1 0 14174 0 1 22842
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_3
timestamp 1723858470
transform 1 0 16480 0 1 22850
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_4
timestamp 1723858470
transform 0 -1 19010 1 0 33386
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_5
timestamp 1723858470
transform 1 0 7546 0 1 22844
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_6
timestamp 1723858470
transform 0 -1 19018 1 0 31080
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_7
timestamp 1723858470
transform 0 -1 19026 1 0 28866
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_8
timestamp 1723858470
transform 0 -1 19008 1 0 26666
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_9
timestamp 1723858470
transform 0 -1 19016 1 0 24452
box -38 -48 1786 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 3278 0 -1 2288
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_1
timestamp 1723858470
transform -1 0 5348 0 -1 2284
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_2
timestamp 1723858470
transform -1 0 7300 0 -1 2284
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_3
timestamp 1723858470
transform -1 0 9302 0 -1 2290
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_4
timestamp 1723858470
transform -1 0 11254 0 -1 2290
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_5
timestamp 1723858470
transform -1 0 13246 0 -1 2290
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_6
timestamp 1723858470
transform -1 0 15198 0 -1 2290
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_7
timestamp 1723858470
transform -1 0 17262 0 -1 2290
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_8
timestamp 1723858470
transform -1 0 5442 0 -1 5540
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_9
timestamp 1723858470
transform -1 0 7394 0 -1 5540
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_10
timestamp 1723858470
transform -1 0 3308 0 -1 5548
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_11
timestamp 1723858470
transform -1 0 9396 0 -1 5546
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_12
timestamp 1723858470
transform -1 0 13552 0 -1 5956
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_13
timestamp 1723858470
transform -1 0 11490 0 -1 5968
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_14
timestamp 1723858470
transform -1 0 15510 0 -1 5964
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_15
timestamp 1723858470
transform -1 0 17504 0 -1 5970
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_16
timestamp 1723858470
transform -1 0 13788 0 -1 5050
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_17
timestamp 1723858470
transform -1 0 11518 0 -1 5094
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_18
timestamp 1723858470
transform -1 0 15790 0 -1 5044
box -38 -48 1510 592
use sky130_fd_sc_hd__fa_1  sky130_fd_sc_hd__fa_1_19
timestamp 1723858470
transform -1 0 17812 0 -1 5026
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1755028488
transform -1 0 6358 0 -1 3340
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1755028488
transform -1 0 6388 0 -1 6600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1755028488
transform -1 0 9706 0 -1 17794
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1755028488
transform 1 0 16336 0 1 16150
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_4
timestamp 1755028488
transform 1 0 17104 0 1 16140
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_5
timestamp 1755028488
transform 1 0 17978 0 1 16142
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_6
timestamp 1755028488
transform 1 0 18592 0 1 16140
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_7
timestamp 1755028488
transform 1 0 19360 0 1 16130
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_8
timestamp 1755028488
transform 1 0 20234 0 1 16132
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_9
timestamp 1755028488
transform 1 0 21356 0 1 16134
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_10
timestamp 1755028488
transform 1 0 22124 0 1 16124
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_11
timestamp 1755028488
transform 1 0 22998 0 1 16126
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_12
timestamp 1755028488
transform -1 0 23283 0 -1 17660
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_13
timestamp 1755028488
transform -1 0 22515 0 -1 17670
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_14
timestamp 1755028488
transform -1 0 21641 0 -1 17668
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_15
timestamp 1755028488
transform -1 0 21027 0 -1 17670
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_16
timestamp 1755028488
transform -1 0 20259 0 -1 17680
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_17
timestamp 1755028488
transform -1 0 19385 0 -1 17678
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_18
timestamp 1755028488
transform -1 0 18263 0 -1 17676
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_19
timestamp 1755028488
transform -1 0 17495 0 -1 17686
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_20
timestamp 1755028488
transform -1 0 16621 0 -1 17684
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_21
timestamp 1755028488
transform -1 0 15843 0 -1 17646
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 0 -1 19166 1 0 36060
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 0 -1 19158 1 0 36764
box -38 -48 498 592
use sky130_fd_sc_hd__inv_6  sky130_fd_sc_hd__inv_6_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 0 -1 19146 1 0 37730
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  sky130_fd_sc_hd__inv_8_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 0 -1 19132 1 0 38808
box -38 -48 866 592
use sky130_fd_sc_hd__inv_12  sky130_fd_sc_hd__inv_12_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 0 -1 19124 1 0 40236
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_16  sky130_fd_sc_hd__inv_16_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 0 -1 19140 1 0 41948
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  sky130_fd_sc_hd__mux2_1_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 19130 0 -1 5396
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  sky130_fd_sc_hd__mux4_1_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 23484 0 1 14288
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 1808 0 -1 2288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1723858470
transform -1 0 3878 0 -1 2284
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1723858470
transform -1 0 5834 0 -1 2284
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1723858470
transform -1 0 7832 0 -1 2290
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1723858470
transform -1 0 9788 0 -1 2290
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1723858470
transform -1 0 11776 0 -1 2290
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1723858470
transform -1 0 13730 0 -1 2290
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1723858470
transform -1 0 19222 0 -1 5396
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1723858470
transform -1 0 6086 0 -1 3340
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1723858470
transform 1 0 25416 0 1 14288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_10
timestamp 1723858470
transform 1 0 23260 0 1 16126
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_11
timestamp 1723858470
transform 1 0 22394 0 1 16124
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_12
timestamp 1723858470
transform 1 0 21616 0 1 16134
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_13
timestamp 1723858470
transform 1 0 20500 0 1 16132
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_14
timestamp 1723858470
transform 1 0 19634 0 1 16130
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_15
timestamp 1723858470
transform 1 0 18864 0 1 16140
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_16
timestamp 1723858470
transform 1 0 17886 0 1 16142
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_17
timestamp 1723858470
transform 1 0 17378 0 1 16140
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_18
timestamp 1723858470
transform 1 0 16246 0 1 16150
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_19
timestamp 1723858470
transform -1 0 6470 0 -1 6600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_20
timestamp 1723858470
transform -1 0 9782 0 -1 17794
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_21
timestamp 1723858470
transform 1 0 4376 0 1 16042
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_22
timestamp 1723858470
transform 1 0 4476 0 1 15298
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_23
timestamp 1723858470
transform 1 0 4386 0 1 14478
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_24
timestamp 1723858470
transform 1 0 4486 0 1 13734
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_25
timestamp 1723858470
transform 1 0 4378 0 1 12810
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_26
timestamp 1723858470
transform 1 0 4478 0 1 12066
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_27
timestamp 1723858470
transform 1 0 4388 0 1 11246
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_28
timestamp 1723858470
transform 1 0 4486 0 1 10502
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_29
timestamp 1723858470
transform 1 0 5852 0 1 11860
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_30
timestamp 1723858470
transform 1 0 5856 0 1 12880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_31
timestamp 1723858470
transform 1 0 5732 0 1 13722
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_32
timestamp 1723858470
transform -1 0 6302 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_33
timestamp 1723858470
transform 1 0 7252 0 1 15188
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_34
timestamp 1723858470
transform 1 0 7250 0 1 13348
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_35
timestamp 1723858470
transform 1 0 8274 0 1 13706
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_36
timestamp 1723858470
transform 1 0 12118 0 1 13352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_37
timestamp 1723858470
transform 1 0 13140 0 1 13710
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_38
timestamp 1723858470
transform 1 0 12118 0 1 15192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_39
timestamp 1723858470
transform 1 0 11076 0 1 14692
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_40
timestamp 1723858470
transform 1 0 9252 0 1 14482
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_41
timestamp 1723858470
transform 1 0 9342 0 1 15302
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_42
timestamp 1723858470
transform 1 0 9242 0 1 16046
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_43
timestamp 1723858470
transform 1 0 10598 0 1 13726
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_44
timestamp 1723858470
transform 1 0 9350 0 1 13738
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_45
timestamp 1723858470
transform 1 0 10722 0 1 12884
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_46
timestamp 1723858470
transform 1 0 10718 0 1 11864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_47
timestamp 1723858470
transform 1 0 9352 0 1 10506
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_48
timestamp 1723858470
transform 1 0 9254 0 1 11250
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_49
timestamp 1723858470
transform 1 0 9342 0 1 12070
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_50
timestamp 1723858470
transform 1 0 9244 0 1 12814
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_51
timestamp 1723858470
transform -1 0 1838 0 -1 5548
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_52
timestamp 1723858470
transform -1 0 15792 0 -1 2290
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_53
timestamp 1723858470
transform -1 0 10020 0 -1 5968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_54
timestamp 1723858470
transform -1 0 11610 0 -1 5094
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_55
timestamp 1723858470
transform -1 0 3972 0 -1 5540
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_56
timestamp 1723858470
transform -1 0 5922 0 -1 5540
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_57
timestamp 1723858470
transform -1 0 7924 0 -1 5546
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_58
timestamp 1723858470
transform -1 0 12080 0 -1 5956
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_59
timestamp 1723858470
transform -1 0 14038 0 -1 5964
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_60
timestamp 1723858470
transform -1 0 16034 0 -1 5970
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_61
timestamp 1723858470
transform -1 0 12320 0 -1 5050
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_62
timestamp 1723858470
transform -1 0 14320 0 -1 5044
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_63
timestamp 1723858470
transform -1 0 16344 0 -1 5026
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_64
timestamp 1723858470
transform -1 0 23373 0 -1 17660
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_65
timestamp 1723858470
transform -1 0 19119 0 -1 17678
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_66
timestamp 1723858470
transform -1 0 19985 0 -1 17680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_67
timestamp 1723858470
transform -1 0 21733 0 -1 17668
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_68
timestamp 1723858470
transform -1 0 20755 0 -1 17670
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_69
timestamp 1723858470
transform -1 0 22241 0 -1 17670
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_70
timestamp 1723858470
transform -1 0 16359 0 -1 17684
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_71
timestamp 1723858470
transform -1 0 17225 0 -1 17686
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_72
timestamp 1723858470
transform -1 0 18003 0 -1 17676
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_73
timestamp 1723858470
transform 1 0 11508 0 1 22852
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_74
timestamp 1723858470
transform 1 0 13708 0 1 22834
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_75
timestamp 1723858470
transform 1 0 15922 0 1 22842
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_76
timestamp 1723858470
transform 1 0 18228 0 1 22850
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_77
timestamp 1723858470
transform 1 0 9294 0 1 22844
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_78
timestamp 1723858470
transform 0 -1 19010 1 0 35134
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_79
timestamp 1723858470
transform 0 -1 19018 1 0 32828
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_80
timestamp 1723858470
transform 0 -1 19026 1 0 30614
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_81
timestamp 1723858470
transform 0 -1 19008 1 0 28414
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_82
timestamp 1723858470
transform 0 -1 19016 1 0 26200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_84
timestamp 1723858470
transform 0 -1 19166 1 0 36336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_85
timestamp 1723858470
transform 0 -1 19158 1 0 37220
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_86
timestamp 1723858470
transform 0 -1 19146 1 0 38374
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_87
timestamp 1723858470
transform 0 -1 19132 1 0 39636
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_88
timestamp 1723858470
transform 0 -1 19124 1 0 41432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_89
timestamp 1723858470
transform 0 -1 19140 1 0 43418
box -38 -48 130 592
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
rlabel metal1 s 16345 17092 16621 17188 5 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 16345 17636 16621 17732 5 VGND
port 2 nsew ground bidirectional abutment
rlabel comment s 16621 17684 16621 17684 8 inv_1
flabel metal1 s 16558 17123 16592 17157 0 FreeSans 200 180 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel metal1 s 16558 17667 16592 17701 0 FreeSans 200 180 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel pwell s 16558 17667 16592 17701 0 FreeSans 200 180 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 16558 17123 16592 17157 0 FreeSans 200 180 0 0 VPB
port 4 nsew power bidirectional
flabel locali s 16515 17429 16549 17463 0 FreeSans 340 180 0 0 A
port 1 nsew signal input
flabel locali s 16423 17429 16457 17463 0 FreeSans 340 180 0 0 Y
port 6 nsew signal output
flabel locali s 16423 17361 16457 17395 0 FreeSans 340 180 0 0 Y
port 6 nsew signal output
rlabel metal1 s 17219 17094 17495 17190 5 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 17219 17638 17495 17734 5 VGND
port 2 nsew ground bidirectional abutment
rlabel comment s 17495 17686 17495 17686 8 inv_1
flabel metal1 s 17432 17125 17466 17159 0 FreeSans 200 180 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel metal1 s 17432 17669 17466 17703 0 FreeSans 200 180 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel pwell s 17432 17669 17466 17703 0 FreeSans 200 180 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 17432 17125 17466 17159 0 FreeSans 200 180 0 0 VPB
port 4 nsew power bidirectional
flabel locali s 17389 17431 17423 17465 0 FreeSans 340 180 0 0 A
port 1 nsew signal input
flabel locali s 17297 17431 17331 17465 0 FreeSans 340 180 0 0 Y
port 6 nsew signal output
flabel locali s 17297 17363 17331 17397 0 FreeSans 340 180 0 0 Y
port 6 nsew signal output
rlabel metal1 s 17987 17084 18263 17180 5 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 17987 17628 18263 17724 5 VGND
port 2 nsew ground bidirectional abutment
rlabel comment s 18263 17676 18263 17676 8 inv_1
flabel metal1 s 18200 17115 18234 17149 0 FreeSans 200 180 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel metal1 s 18200 17659 18234 17693 0 FreeSans 200 180 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel pwell s 18200 17659 18234 17693 0 FreeSans 200 180 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 18200 17115 18234 17149 0 FreeSans 200 180 0 0 VPB
port 4 nsew power bidirectional
flabel locali s 18157 17421 18191 17455 0 FreeSans 340 180 0 0 A
port 1 nsew signal input
flabel locali s 18065 17421 18099 17455 0 FreeSans 340 180 0 0 Y
port 6 nsew signal output
flabel locali s 18065 17353 18099 17387 0 FreeSans 340 180 0 0 Y
port 6 nsew signal output
rlabel metal1 s 17911 17084 18003 17180 5 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 17911 17628 18003 17724 5 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 18003 17676 18003 17676 8 tapvpwrvgnd_1
flabel metal1 s 17931 17656 17982 17694 0 FreeSans 200 180 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 17928 17123 17981 17152 0 FreeSans 200 180 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 17133 17094 17225 17190 5 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 17133 17638 17225 17734 5 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 17225 17686 17225 17686 8 tapvpwrvgnd_1
flabel metal1 s 17153 17666 17204 17704 0 FreeSans 200 180 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 17150 17133 17203 17162 0 FreeSans 200 180 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 16267 17092 16359 17188 5 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 16267 17636 16359 17732 5 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 16359 17684 16359 17684 8 tapvpwrvgnd_1
flabel metal1 s 16287 17664 16338 17702 0 FreeSans 200 180 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 16284 17131 16337 17160 0 FreeSans 200 180 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 19109 17086 19385 17182 5 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 19109 17630 19385 17726 5 VGND
port 2 nsew ground bidirectional abutment
rlabel comment s 19385 17678 19385 17678 8 inv_1
flabel metal1 s 19322 17117 19356 17151 0 FreeSans 200 180 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel metal1 s 19322 17661 19356 17695 0 FreeSans 200 180 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel pwell s 19322 17661 19356 17695 0 FreeSans 200 180 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 19322 17117 19356 17151 0 FreeSans 200 180 0 0 VPB
port 4 nsew power bidirectional
flabel locali s 19279 17423 19313 17457 0 FreeSans 340 180 0 0 A
port 1 nsew signal input
flabel locali s 19187 17423 19221 17457 0 FreeSans 340 180 0 0 Y
port 6 nsew signal output
flabel locali s 19187 17355 19221 17389 0 FreeSans 340 180 0 0 Y
port 6 nsew signal output
rlabel metal1 s 19983 17088 20259 17184 5 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 19983 17632 20259 17728 5 VGND
port 2 nsew ground bidirectional abutment
rlabel comment s 20259 17680 20259 17680 8 inv_1
flabel metal1 s 20196 17119 20230 17153 0 FreeSans 200 180 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel metal1 s 20196 17663 20230 17697 0 FreeSans 200 180 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel pwell s 20196 17663 20230 17697 0 FreeSans 200 180 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 20196 17119 20230 17153 0 FreeSans 200 180 0 0 VPB
port 4 nsew power bidirectional
flabel locali s 20153 17425 20187 17459 0 FreeSans 340 180 0 0 A
port 1 nsew signal input
flabel locali s 20061 17425 20095 17459 0 FreeSans 340 180 0 0 Y
port 6 nsew signal output
flabel locali s 20061 17357 20095 17391 0 FreeSans 340 180 0 0 Y
port 6 nsew signal output
rlabel metal1 s 20751 17078 21027 17174 5 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 20751 17622 21027 17718 5 VGND
port 2 nsew ground bidirectional abutment
rlabel comment s 21027 17670 21027 17670 8 inv_1
flabel metal1 s 20964 17109 20998 17143 0 FreeSans 200 180 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel metal1 s 20964 17653 20998 17687 0 FreeSans 200 180 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel pwell s 20964 17653 20998 17687 0 FreeSans 200 180 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 20964 17109 20998 17143 0 FreeSans 200 180 0 0 VPB
port 4 nsew power bidirectional
flabel locali s 20921 17415 20955 17449 0 FreeSans 340 180 0 0 A
port 1 nsew signal input
flabel locali s 20829 17415 20863 17449 0 FreeSans 340 180 0 0 Y
port 6 nsew signal output
flabel locali s 20829 17347 20863 17381 0 FreeSans 340 180 0 0 Y
port 6 nsew signal output
rlabel metal1 s 21365 17076 21641 17172 5 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 21365 17620 21641 17716 5 VGND
port 2 nsew ground bidirectional abutment
rlabel comment s 21641 17668 21641 17668 8 inv_1
flabel metal1 s 21578 17107 21612 17141 0 FreeSans 200 180 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel metal1 s 21578 17651 21612 17685 0 FreeSans 200 180 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel pwell s 21578 17651 21612 17685 0 FreeSans 200 180 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 21578 17107 21612 17141 0 FreeSans 200 180 0 0 VPB
port 4 nsew power bidirectional
flabel locali s 21535 17413 21569 17447 0 FreeSans 340 180 0 0 A
port 1 nsew signal input
flabel locali s 21443 17413 21477 17447 0 FreeSans 340 180 0 0 Y
port 6 nsew signal output
flabel locali s 21443 17345 21477 17379 0 FreeSans 340 180 0 0 Y
port 6 nsew signal output
rlabel metal1 s 22149 17078 22241 17174 5 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 22149 17622 22241 17718 5 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 22241 17670 22241 17670 8 tapvpwrvgnd_1
flabel metal1 s 22169 17650 22220 17688 0 FreeSans 200 180 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 22166 17117 22219 17146 0 FreeSans 200 180 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 20663 17078 20755 17174 5 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 20663 17622 20755 17718 5 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 20755 17670 20755 17670 8 tapvpwrvgnd_1
flabel metal1 s 20683 17650 20734 17688 0 FreeSans 200 180 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 20680 17117 20733 17146 0 FreeSans 200 180 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 21641 17076 21733 17172 5 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 21641 17620 21733 17716 5 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 21733 17668 21733 17668 8 tapvpwrvgnd_1
flabel metal1 s 21661 17648 21712 17686 0 FreeSans 200 180 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 21658 17115 21711 17144 0 FreeSans 200 180 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 19893 17088 19985 17184 5 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 19893 17632 19985 17728 5 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 19985 17680 19985 17680 8 tapvpwrvgnd_1
flabel metal1 s 19913 17660 19964 17698 0 FreeSans 200 180 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 19910 17127 19963 17156 0 FreeSans 200 180 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 19027 17086 19119 17182 5 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 19027 17630 19119 17726 5 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 19119 17678 19119 17678 8 tapvpwrvgnd_1
flabel metal1 s 19047 17658 19098 17696 0 FreeSans 200 180 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 19044 17125 19097 17154 0 FreeSans 200 180 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 22239 17078 22515 17174 5 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 22239 17622 22515 17718 5 VGND
port 2 nsew ground bidirectional abutment
rlabel comment s 22515 17670 22515 17670 8 inv_1
flabel metal1 s 22452 17109 22486 17143 0 FreeSans 200 180 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel metal1 s 22452 17653 22486 17687 0 FreeSans 200 180 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel pwell s 22452 17653 22486 17687 0 FreeSans 200 180 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 22452 17109 22486 17143 0 FreeSans 200 180 0 0 VPB
port 4 nsew power bidirectional
flabel locali s 22409 17415 22443 17449 0 FreeSans 340 180 0 0 A
port 1 nsew signal input
flabel locali s 22317 17415 22351 17449 0 FreeSans 340 180 0 0 Y
port 6 nsew signal output
flabel locali s 22317 17347 22351 17381 0 FreeSans 340 180 0 0 Y
port 6 nsew signal output
rlabel metal1 s 23007 17068 23283 17164 5 VPWR
port 5 nsew power bidirectional abutment
rlabel metal1 s 23007 17612 23283 17708 5 VGND
port 2 nsew ground bidirectional abutment
rlabel comment s 23283 17660 23283 17660 8 inv_1
flabel metal1 s 23220 17099 23254 17133 0 FreeSans 200 180 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel metal1 s 23220 17643 23254 17677 0 FreeSans 200 180 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel pwell s 23220 17643 23254 17677 0 FreeSans 200 180 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 23220 17099 23254 17133 0 FreeSans 200 180 0 0 VPB
port 4 nsew power bidirectional
flabel locali s 23177 17405 23211 17439 0 FreeSans 340 180 0 0 A
port 1 nsew signal input
flabel locali s 23085 17405 23119 17439 0 FreeSans 340 180 0 0 Y
port 6 nsew signal output
flabel locali s 23085 17337 23119 17371 0 FreeSans 340 180 0 0 Y
port 6 nsew signal output
rlabel metal1 s 23281 17068 23373 17164 5 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 23281 17612 23373 17708 5 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 23373 17660 23373 17660 8 tapvpwrvgnd_1
flabel metal1 s 23301 17640 23352 17678 0 FreeSans 200 180 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 23298 17107 23351 17136 0 FreeSans 200 180 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel locali s 15645 17323 15679 17357 0 FreeSans 340 180 0 0 Y
port 6 nsew signal output
flabel locali s 15645 17391 15679 17425 0 FreeSans 340 180 0 0 Y
port 6 nsew signal output
flabel locali s 15737 17391 15771 17425 0 FreeSans 340 180 0 0 A
port 1 nsew signal input
flabel nwell s 15780 17085 15814 17119 0 FreeSans 200 180 0 0 VPB
port 4 nsew power bidirectional
flabel pwell s 15780 17629 15814 17663 0 FreeSans 200 180 0 0 VNB
port 3 nsew ground bidirectional
flabel metal1 s 15780 17629 15814 17663 0 FreeSans 200 180 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel metal1 s 15780 17085 15814 17119 0 FreeSans 200 180 0 0 VPWR
port 5 nsew power bidirectional abutment
rlabel comment s 15843 17646 15843 17646 8 inv_1
rlabel metal1 s 15567 17598 15843 17694 5 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 15567 17054 15843 17150 5 VPWR
port 5 nsew power bidirectional abutment
flabel metal1 s 15498 17093 15551 17122 0 FreeSans 200 180 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 15501 17626 15552 17664 0 FreeSans 200 180 0 0 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 15573 17646 15573 17646 8 tapvpwrvgnd_1
rlabel metal1 s 15481 17598 15573 17694 5 VGND
port 1 nsew ground bidirectional abutment
rlabel metal1 s 15481 17054 15573 17150 5 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 7575 22827 7609 22861 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 7575 23371 7609 23405 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel locali s 9231 23148 9265 23182 0 FreeSans 400 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 7835 23065 7869 23099 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 7575 23065 7609 23099 0 FreeSans 400 0 0 0 CLK
port 1 nsew clock input
flabel locali s 8936 22929 8970 22963 0 FreeSans 400 0 0 0 Q
port 7 nsew signal output
flabel pwell s 7575 22827 7609 22861 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel pwell s 7592 22844 7592 22844 0 FreeSans 200 0 0 0 VNB
flabel nwell s 7575 23371 7609 23405 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel nwell s 7592 23388 7592 23388 0 FreeSans 200 0 0 0 VPB
rlabel comment s 7546 22844 7546 22844 4 dfxbp_1
rlabel metal1 s 7546 22796 9294 22892 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 7546 23340 9294 23436 1 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 9316 23368 9369 23397 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 9315 22826 9366 22864 0 FreeSans 200 0 0 0 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 9294 22844 9294 22844 4 tapvpwrvgnd_1
rlabel metal1 s 9294 22796 9386 22892 1 VGND
port 1 nsew ground bidirectional abutment
rlabel metal1 s 9294 23340 9386 23436 1 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 9760 23348 11508 23444 1 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 9760 22804 11508 22900 1 VGND
port 3 nsew ground bidirectional abutment
rlabel comment s 9760 22852 9760 22852 4 dfxbp_1
flabel nwell s 9806 23396 9806 23396 0 FreeSans 200 0 0 0 VPB
flabel nwell s 9789 23379 9823 23413 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 9806 22852 9806 22852 0 FreeSans 200 0 0 0 VNB
flabel pwell s 9789 22835 9823 22869 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel locali s 11150 22937 11184 22971 0 FreeSans 400 0 0 0 Q
port 7 nsew signal output
flabel locali s 9789 23073 9823 23107 0 FreeSans 400 0 0 0 CLK
port 1 nsew clock input
flabel locali s 10049 23073 10083 23107 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 11445 23156 11479 23190 0 FreeSans 400 0 0 0 Q_N
port 8 nsew signal output
flabel metal1 s 9789 23379 9823 23413 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 9789 22835 9823 22869 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 11508 23348 11600 23444 1 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 11508 22804 11600 22900 1 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 11508 22852 11508 22852 4 tapvpwrvgnd_1
flabel metal1 s 11529 22834 11580 22872 0 FreeSans 200 0 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 11530 23376 11583 23405 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 13730 23358 13783 23387 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 13729 22816 13780 22854 0 FreeSans 200 0 0 0 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 13708 22834 13708 22834 4 tapvpwrvgnd_1
rlabel metal1 s 13708 22786 13800 22882 1 VGND
port 1 nsew ground bidirectional abutment
rlabel metal1 s 13708 23330 13800 23426 1 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 11989 22817 12023 22851 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 11989 23361 12023 23395 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel locali s 13645 23138 13679 23172 0 FreeSans 400 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 12249 23055 12283 23089 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 11989 23055 12023 23089 0 FreeSans 400 0 0 0 CLK
port 1 nsew clock input
flabel locali s 13350 22919 13384 22953 0 FreeSans 400 0 0 0 Q
port 7 nsew signal output
flabel pwell s 11989 22817 12023 22851 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel pwell s 12006 22834 12006 22834 0 FreeSans 200 0 0 0 VNB
flabel nwell s 11989 23361 12023 23395 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel nwell s 12006 23378 12006 23378 0 FreeSans 200 0 0 0 VPB
rlabel comment s 11960 22834 11960 22834 4 dfxbp_1
rlabel metal1 s 11960 22786 13708 22882 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 11960 23330 13708 23426 1 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 14203 22825 14237 22859 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 14203 23369 14237 23403 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel locali s 15859 23146 15893 23180 0 FreeSans 400 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 14463 23063 14497 23097 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 14203 23063 14237 23097 0 FreeSans 400 0 0 0 CLK
port 1 nsew clock input
flabel locali s 15564 22927 15598 22961 0 FreeSans 400 0 0 0 Q
port 7 nsew signal output
flabel pwell s 14203 22825 14237 22859 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel pwell s 14220 22842 14220 22842 0 FreeSans 200 0 0 0 VNB
flabel nwell s 14203 23369 14237 23403 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel nwell s 14220 23386 14220 23386 0 FreeSans 200 0 0 0 VPB
rlabel comment s 14174 22842 14174 22842 4 dfxbp_1
rlabel metal1 s 14174 22794 15922 22890 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 14174 23338 15922 23434 1 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 15944 23366 15997 23395 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 15943 22824 15994 22862 0 FreeSans 200 0 0 0 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 15922 22842 15922 22842 4 tapvpwrvgnd_1
rlabel metal1 s 15922 22794 16014 22890 1 VGND
port 1 nsew ground bidirectional abutment
rlabel metal1 s 15922 23338 16014 23434 1 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 18250 23374 18303 23403 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 18249 22832 18300 22870 0 FreeSans 200 0 0 0 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 18228 22850 18228 22850 4 tapvpwrvgnd_1
rlabel metal1 s 18228 22802 18320 22898 1 VGND
port 1 nsew ground bidirectional abutment
rlabel metal1 s 18228 23346 18320 23442 1 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 16509 22833 16543 22867 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 16509 23377 16543 23411 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel locali s 18165 23154 18199 23188 0 FreeSans 400 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 16769 23071 16803 23105 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 16509 23071 16543 23105 0 FreeSans 400 0 0 0 CLK
port 1 nsew clock input
flabel locali s 17870 22935 17904 22969 0 FreeSans 400 0 0 0 Q
port 7 nsew signal output
flabel pwell s 16509 22833 16543 22867 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel pwell s 16526 22850 16526 22850 0 FreeSans 200 0 0 0 VNB
flabel nwell s 16509 23377 16543 23411 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel nwell s 16526 23394 16526 23394 0 FreeSans 200 0 0 0 VPB
rlabel comment s 16480 22850 16480 22850 4 dfxbp_1
rlabel metal1 s 16480 22802 18228 22898 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 16480 23346 18228 23442 1 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 18418 35134 18514 35226 7 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 18962 35134 19058 35226 7 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 19010 35134 19010 35134 2 tapvpwrvgnd_1
flabel metal1 s 18990 35155 19028 35206 0 FreeSans 200 270 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 18457 35156 18486 35209 0 FreeSans 200 270 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 18434 30614 18530 30706 7 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 18978 30614 19074 30706 7 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 19026 30614 19026 30614 2 tapvpwrvgnd_1
flabel metal1 s 19006 30635 19044 30686 0 FreeSans 200 270 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 18473 30636 18502 30689 0 FreeSans 200 270 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 18426 31080 18522 32828 7 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 18970 31080 19066 32828 7 VGND
port 3 nsew ground bidirectional abutment
rlabel comment s 19018 31080 19018 31080 2 dfxbp_1
flabel nwell s 18474 31126 18474 31126 0 FreeSans 200 270 0 0 VPB
flabel nwell s 18457 31109 18491 31143 0 FreeSans 200 270 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 19018 31126 19018 31126 0 FreeSans 200 270 0 0 VNB
flabel pwell s 19001 31109 19035 31143 0 FreeSans 200 270 0 0 VNB
port 4 nsew ground bidirectional
flabel locali s 18899 32470 18933 32504 0 FreeSans 400 270 0 0 Q
port 7 nsew signal output
flabel locali s 18763 31109 18797 31143 0 FreeSans 400 270 0 0 CLK
port 1 nsew clock input
flabel locali s 18763 31369 18797 31403 0 FreeSans 200 270 0 0 D
port 2 nsew signal input
flabel locali s 18680 32765 18714 32799 0 FreeSans 400 270 0 0 Q_N
port 8 nsew signal output
flabel metal1 s 18457 31109 18491 31143 0 FreeSans 200 270 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 19001 31109 19035 31143 0 FreeSans 200 270 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 18426 32828 18522 32920 7 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 18970 32828 19066 32920 7 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 19018 32828 19018 32828 2 tapvpwrvgnd_1
flabel metal1 s 18998 32849 19036 32900 0 FreeSans 200 270 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 18465 32850 18494 32903 0 FreeSans 200 270 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 18418 33386 18514 35134 7 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 18962 33386 19058 35134 7 VGND
port 3 nsew ground bidirectional abutment
rlabel comment s 19010 33386 19010 33386 2 dfxbp_1
flabel nwell s 18466 33432 18466 33432 0 FreeSans 200 270 0 0 VPB
flabel nwell s 18449 33415 18483 33449 0 FreeSans 200 270 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 19010 33432 19010 33432 0 FreeSans 200 270 0 0 VNB
flabel pwell s 18993 33415 19027 33449 0 FreeSans 200 270 0 0 VNB
port 4 nsew ground bidirectional
flabel locali s 18891 34776 18925 34810 0 FreeSans 400 270 0 0 Q
port 7 nsew signal output
flabel locali s 18755 33415 18789 33449 0 FreeSans 400 270 0 0 CLK
port 1 nsew clock input
flabel locali s 18755 33675 18789 33709 0 FreeSans 200 270 0 0 D
port 2 nsew signal input
flabel locali s 18672 35071 18706 35105 0 FreeSans 400 270 0 0 Q_N
port 8 nsew signal output
flabel metal1 s 18449 33415 18483 33449 0 FreeSans 200 270 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 18993 33415 19027 33449 0 FreeSans 200 270 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 18416 28414 18512 28506 7 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 18960 28414 19056 28506 7 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 19008 28414 19008 28414 2 tapvpwrvgnd_1
flabel metal1 s 18988 28435 19026 28486 0 FreeSans 200 270 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 18455 28436 18484 28489 0 FreeSans 200 270 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 18416 26666 18512 28414 7 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 18960 26666 19056 28414 7 VGND
port 3 nsew ground bidirectional abutment
rlabel comment s 19008 26666 19008 26666 2 dfxbp_1
flabel nwell s 18464 26712 18464 26712 0 FreeSans 200 270 0 0 VPB
flabel nwell s 18447 26695 18481 26729 0 FreeSans 200 270 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 19008 26712 19008 26712 0 FreeSans 200 270 0 0 VNB
flabel pwell s 18991 26695 19025 26729 0 FreeSans 200 270 0 0 VNB
port 4 nsew ground bidirectional
flabel locali s 18889 28056 18923 28090 0 FreeSans 400 270 0 0 Q
port 7 nsew signal output
flabel locali s 18753 26695 18787 26729 0 FreeSans 400 270 0 0 CLK
port 1 nsew clock input
flabel locali s 18753 26955 18787 26989 0 FreeSans 200 270 0 0 D
port 2 nsew signal input
flabel locali s 18670 28351 18704 28385 0 FreeSans 400 270 0 0 Q_N
port 8 nsew signal output
flabel metal1 s 18447 26695 18481 26729 0 FreeSans 200 270 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 18991 26695 19025 26729 0 FreeSans 200 270 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 18434 28866 18530 30614 7 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 18978 28866 19074 30614 7 VGND
port 3 nsew ground bidirectional abutment
rlabel comment s 19026 28866 19026 28866 2 dfxbp_1
flabel nwell s 18482 28912 18482 28912 0 FreeSans 200 270 0 0 VPB
flabel nwell s 18465 28895 18499 28929 0 FreeSans 200 270 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 19026 28912 19026 28912 0 FreeSans 200 270 0 0 VNB
flabel pwell s 19009 28895 19043 28929 0 FreeSans 200 270 0 0 VNB
port 4 nsew ground bidirectional
flabel locali s 18907 30256 18941 30290 0 FreeSans 400 270 0 0 Q
port 7 nsew signal output
flabel locali s 18771 28895 18805 28929 0 FreeSans 400 270 0 0 CLK
port 1 nsew clock input
flabel locali s 18771 29155 18805 29189 0 FreeSans 200 270 0 0 D
port 2 nsew signal input
flabel locali s 18688 30551 18722 30585 0 FreeSans 400 270 0 0 Q_N
port 8 nsew signal output
flabel metal1 s 18465 28895 18499 28929 0 FreeSans 200 270 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 19009 28895 19043 28929 0 FreeSans 200 270 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 18424 24452 18520 26200 7 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 18968 24452 19064 26200 7 VGND
port 3 nsew ground bidirectional abutment
rlabel comment s 19016 24452 19016 24452 2 dfxbp_1
flabel nwell s 18472 24498 18472 24498 0 FreeSans 200 270 0 0 VPB
flabel nwell s 18455 24481 18489 24515 0 FreeSans 200 270 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 19016 24498 19016 24498 0 FreeSans 200 270 0 0 VNB
flabel pwell s 18999 24481 19033 24515 0 FreeSans 200 270 0 0 VNB
port 4 nsew ground bidirectional
flabel locali s 18897 25842 18931 25876 0 FreeSans 400 270 0 0 Q
port 7 nsew signal output
flabel locali s 18761 24481 18795 24515 0 FreeSans 400 270 0 0 CLK
port 1 nsew clock input
flabel locali s 18761 24741 18795 24775 0 FreeSans 200 270 0 0 D
port 2 nsew signal input
flabel locali s 18678 26137 18712 26171 0 FreeSans 400 270 0 0 Q_N
port 8 nsew signal output
flabel metal1 s 18455 24481 18489 24515 0 FreeSans 200 270 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 18999 24481 19033 24515 0 FreeSans 200 270 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 18424 26200 18520 26292 7 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 18968 26200 19064 26292 7 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 19016 26200 19016 26200 2 tapvpwrvgnd_1
flabel metal1 s 18996 26221 19034 26272 0 FreeSans 200 270 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 18463 26222 18492 26275 0 FreeSans 200 270 0 0 VPWR
port 2 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
