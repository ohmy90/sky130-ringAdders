VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_ohmy90_ringOscillator
  CLASS BLOCK ;
  FOREIGN tt_um_ohmy90_ringOscillator ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
    PORT
      LAYER li1 ;
        RECT 22.275 14.290 22.445 14.460 ;
    END
    PORT
      LAYER li1 ;
        RECT 11.965 14.310 12.135 14.480 ;
    END
    PORT
      LAYER li1 ;
        RECT 32.645 14.280 32.815 14.450 ;
    END
    PORT
      LAYER li1 ;
        RECT 42.955 14.260 43.125 14.430 ;
    END
    PORT
      LAYER li1 ;
        RECT 73.935 14.210 74.105 14.380 ;
    END
    PORT
      LAYER li1 ;
        RECT 84.245 14.190 84.415 14.360 ;
    END
    PORT
      LAYER li1 ;
        RECT 63.565 14.220 63.735 14.390 ;
    END
    PORT
      LAYER li1 ;
        RECT 53.255 14.240 53.425 14.410 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
    PORT
      LAYER li1 ;
        RECT 24.675 14.660 24.845 14.830 ;
    END
    PORT
      LAYER li1 ;
        RECT 14.365 14.680 14.535 14.850 ;
    END
    PORT
      LAYER li1 ;
        RECT 35.045 14.650 35.215 14.820 ;
    END
    PORT
      LAYER li1 ;
        RECT 45.355 14.630 45.525 14.800 ;
    END
    PORT
      LAYER li1 ;
        RECT 76.335 14.580 76.505 14.750 ;
    END
    PORT
      LAYER li1 ;
        RECT 86.645 14.560 86.815 14.730 ;
    END
    PORT
      LAYER li1 ;
        RECT 65.965 14.590 66.135 14.760 ;
    END
    PORT
      LAYER li1 ;
        RECT 55.655 14.610 55.825 14.780 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.541300 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 11.485 14.680 11.655 14.850 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.800 13.080 26.440 13.325 ;
    END
    PORT
      LAYER met1 ;
        RECT 7.490 13.100 16.130 13.345 ;
    END
    PORT
      LAYER met1 ;
        RECT 28.170 13.070 36.810 13.315 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.480 13.050 47.120 13.295 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.460 13.000 78.100 13.245 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.770 12.980 88.410 13.225 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.090 13.010 67.730 13.255 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.780 13.030 57.420 13.275 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
    PORT
      LAYER pwell ;
        RECT 17.800 13.080 26.440 13.325 ;
    END
    PORT
      LAYER pwell ;
        RECT 7.490 13.100 16.130 13.345 ;
    END
    PORT
      LAYER pwell ;
        RECT 28.170 13.070 36.810 13.315 ;
    END
    PORT
      LAYER pwell ;
        RECT 38.480 13.050 47.120 13.295 ;
    END
    PORT
      LAYER pwell ;
        RECT 69.460 13.000 78.100 13.245 ;
    END
    PORT
      LAYER pwell ;
        RECT 79.770 12.980 88.410 13.225 ;
    END
    PORT
      LAYER pwell ;
        RECT 59.090 13.010 67.730 13.255 ;
    END
    PORT
      LAYER pwell ;
        RECT 48.780 13.030 57.420 13.275 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
    PORT
      LAYER nwell ;
        RECT 17.800 16.165 26.440 16.410 ;
    END
    PORT
      LAYER nwell ;
        RECT 7.490 16.185 16.130 16.430 ;
    END
    PORT
      LAYER nwell ;
        RECT 28.170 16.155 36.810 16.400 ;
    END
    PORT
      LAYER nwell ;
        RECT 38.480 16.135 47.120 16.380 ;
    END
    PORT
      LAYER nwell ;
        RECT 69.460 16.085 78.100 16.330 ;
    END
    PORT
      LAYER nwell ;
        RECT 79.770 16.065 88.410 16.310 ;
    END
    PORT
      LAYER nwell ;
        RECT 59.090 16.095 67.730 16.340 ;
    END
    PORT
      LAYER nwell ;
        RECT 48.780 16.115 57.420 16.360 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
    PORT
      LAYER met1 ;
        RECT 17.800 16.165 26.440 16.410 ;
    END
    PORT
      LAYER met1 ;
        RECT 7.490 16.185 16.130 16.430 ;
    END
    PORT
      LAYER met1 ;
        RECT 28.170 16.155 36.810 16.400 ;
    END
    PORT
      LAYER met1 ;
        RECT 38.480 16.135 47.120 16.380 ;
    END
    PORT
      LAYER met1 ;
        RECT 69.460 16.085 78.100 16.330 ;
    END
    PORT
      LAYER met1 ;
        RECT 79.770 16.065 88.410 16.310 ;
    END
    PORT
      LAYER met1 ;
        RECT 59.090 16.095 67.730 16.340 ;
    END
    PORT
      LAYER met1 ;
        RECT 48.780 16.115 57.420 16.360 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
    PORT
      LAYER li1 ;
        RECT 88.085 13.450 88.255 13.620 ;
    END
    PORT
      LAYER li1 ;
        RECT 88.085 13.820 88.255 13.990 ;
    END
    PORT
      LAYER li1 ;
        RECT 88.085 14.190 88.255 14.360 ;
    END
    PORT
      LAYER li1 ;
        RECT 88.085 14.560 88.255 14.730 ;
    END
    PORT
      LAYER li1 ;
        RECT 88.085 14.930 88.255 15.100 ;
    END
    PORT
      LAYER li1 ;
        RECT 88.085 15.300 88.255 15.470 ;
    END
    PORT
      LAYER li1 ;
        RECT 88.085 15.670 88.255 15.840 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
    PORT
      LAYER li1 ;
        RECT 17.955 13.550 18.125 13.720 ;
    END
    PORT
      LAYER li1 ;
        RECT 17.955 13.920 18.125 14.090 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.645 13.570 7.815 13.740 ;
    END
    PORT
      LAYER li1 ;
        RECT 7.645 13.940 7.815 14.110 ;
    END
    PORT
      LAYER li1 ;
        RECT 28.325 13.910 28.495 14.080 ;
    END
    PORT
      LAYER li1 ;
        RECT 28.325 13.540 28.495 13.710 ;
    END
    PORT
      LAYER li1 ;
        RECT 38.635 13.890 38.805 14.060 ;
    END
    PORT
      LAYER li1 ;
        RECT 38.635 13.520 38.805 13.690 ;
    END
    PORT
      LAYER li1 ;
        RECT 69.615 13.470 69.785 13.640 ;
    END
    PORT
      LAYER li1 ;
        RECT 69.615 13.840 69.785 14.010 ;
    END
    PORT
      LAYER li1 ;
        RECT 79.925 13.450 80.095 13.620 ;
    END
    PORT
      LAYER li1 ;
        RECT 79.925 13.820 80.095 13.990 ;
    END
    PORT
      LAYER li1 ;
        RECT 59.245 13.480 59.415 13.650 ;
    END
    PORT
      LAYER li1 ;
        RECT 59.245 13.850 59.415 14.020 ;
    END
    PORT
      LAYER li1 ;
        RECT 48.935 13.500 49.105 13.670 ;
    END
    PORT
      LAYER li1 ;
        RECT 48.935 13.870 49.105 14.040 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.469500 ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 7.150 34.575 16.170 36.435 ;
        RECT 8.840 34.470 14.820 34.575 ;
        RECT 17.560 34.415 26.580 36.275 ;
        RECT 27.860 34.555 36.880 36.415 ;
        RECT 38.170 34.585 47.190 36.445 ;
        RECT 29.550 34.450 35.530 34.555 ;
        RECT 39.860 34.480 45.840 34.585 ;
        RECT 19.250 34.310 25.230 34.415 ;
      LAYER pwell ;
        RECT 7.345 34.060 8.290 34.155 ;
        RECT 15.030 34.060 15.975 34.155 ;
        RECT 7.345 33.160 15.975 34.060 ;
        RECT 28.055 34.040 29.000 34.135 ;
        RECT 35.740 34.040 36.685 34.135 ;
        RECT 17.755 33.900 18.700 33.995 ;
        RECT 25.440 33.900 26.385 33.995 ;
        RECT 7.340 32.915 15.980 33.160 ;
        RECT 17.755 33.000 26.385 33.900 ;
        RECT 28.055 33.140 36.685 34.040 ;
        RECT 38.365 34.070 39.310 34.165 ;
        RECT 46.050 34.070 46.995 34.165 ;
        RECT 38.365 33.170 46.995 34.070 ;
        RECT 17.750 32.755 26.390 33.000 ;
        RECT 28.050 32.895 36.690 33.140 ;
        RECT 38.360 32.925 47.000 33.170 ;
        RECT 46.145 32.120 46.390 32.140 ;
        RECT 46.145 30.710 47.385 32.120 ;
        RECT 46.145 30.700 46.390 30.710 ;
      LAYER nwell ;
        RECT 47.805 30.510 49.665 32.330 ;
      LAYER pwell ;
        RECT 7.260 30.070 15.900 30.315 ;
        RECT 17.580 30.150 26.220 30.395 ;
        RECT 7.265 29.170 15.895 30.070 ;
        RECT 7.265 29.075 8.210 29.170 ;
        RECT 14.950 29.075 15.895 29.170 ;
        RECT 17.585 29.250 26.215 30.150 ;
        RECT 27.890 29.990 36.530 30.235 ;
        RECT 17.585 29.155 18.530 29.250 ;
        RECT 25.270 29.155 26.215 29.250 ;
        RECT 27.895 29.090 36.525 29.990 ;
        RECT 38.260 29.960 46.900 30.205 ;
        RECT 27.895 28.995 28.840 29.090 ;
        RECT 35.580 28.995 36.525 29.090 ;
        RECT 38.265 29.060 46.895 29.960 ;
        RECT 38.265 28.965 39.210 29.060 ;
        RECT 45.950 28.965 46.895 29.060 ;
      LAYER nwell ;
        RECT 84.400 28.900 89.100 30.760 ;
        RECT 8.420 28.655 14.400 28.760 ;
        RECT 18.740 28.735 24.720 28.840 ;
        RECT 7.070 26.795 16.090 28.655 ;
        RECT 17.390 26.875 26.410 28.735 ;
        RECT 29.050 28.575 35.030 28.680 ;
        RECT 27.700 26.715 36.720 28.575 ;
        RECT 39.420 28.545 45.400 28.650 ;
        RECT 38.070 26.685 47.090 28.545 ;
      LAYER pwell ;
        RECT 84.595 27.485 88.895 28.480 ;
        RECT 84.590 27.240 88.910 27.485 ;
        RECT 40.490 22.015 41.930 22.260 ;
        RECT 40.500 21.020 41.910 22.015 ;
      LAYER nwell ;
        RECT 40.300 18.740 42.120 20.600 ;
        RECT 7.300 16.430 16.320 16.620 ;
        RECT 7.300 16.185 7.490 16.430 ;
        RECT 16.130 16.185 16.320 16.430 ;
        RECT 7.300 14.760 16.320 16.185 ;
        RECT 17.610 16.410 26.630 16.600 ;
        RECT 17.610 16.165 17.800 16.410 ;
        RECT 26.440 16.165 26.630 16.410 ;
        RECT 8.990 14.655 14.970 14.760 ;
        RECT 17.610 14.740 26.630 16.165 ;
        RECT 27.980 16.400 37.000 16.590 ;
        RECT 27.980 16.155 28.170 16.400 ;
        RECT 36.810 16.155 37.000 16.400 ;
        RECT 19.300 14.635 25.280 14.740 ;
        RECT 27.980 14.730 37.000 16.155 ;
        RECT 38.290 16.380 47.310 16.570 ;
        RECT 38.290 16.135 38.480 16.380 ;
        RECT 47.120 16.135 47.310 16.380 ;
        RECT 29.670 14.625 35.650 14.730 ;
        RECT 38.290 14.710 47.310 16.135 ;
        RECT 48.590 16.360 57.610 16.550 ;
        RECT 48.590 16.115 48.780 16.360 ;
        RECT 57.420 16.115 57.610 16.360 ;
        RECT 39.980 14.605 45.960 14.710 ;
        RECT 48.590 14.690 57.610 16.115 ;
        RECT 58.900 16.340 67.920 16.530 ;
        RECT 58.900 16.095 59.090 16.340 ;
        RECT 67.730 16.095 67.920 16.340 ;
        RECT 50.280 14.585 56.260 14.690 ;
        RECT 58.900 14.670 67.920 16.095 ;
        RECT 69.270 16.330 78.290 16.520 ;
        RECT 69.270 16.085 69.460 16.330 ;
        RECT 78.100 16.085 78.290 16.330 ;
        RECT 60.590 14.565 66.570 14.670 ;
        RECT 69.270 14.660 78.290 16.085 ;
        RECT 79.580 16.310 88.600 16.500 ;
        RECT 79.580 16.065 79.770 16.310 ;
        RECT 88.410 16.065 88.600 16.310 ;
        RECT 70.960 14.555 76.940 14.660 ;
        RECT 79.580 14.640 88.600 16.065 ;
        RECT 81.270 14.535 87.250 14.640 ;
      LAYER pwell ;
        RECT 7.495 14.245 8.440 14.340 ;
        RECT 15.180 14.245 16.125 14.340 ;
        RECT 7.495 13.345 16.125 14.245 ;
        RECT 17.805 14.225 18.750 14.320 ;
        RECT 25.490 14.225 26.435 14.320 ;
        RECT 17.805 13.325 26.435 14.225 ;
        RECT 28.175 14.215 29.120 14.310 ;
        RECT 35.860 14.215 36.805 14.310 ;
        RECT 28.175 13.315 36.805 14.215 ;
        RECT 38.485 14.195 39.430 14.290 ;
        RECT 46.170 14.195 47.115 14.290 ;
        RECT 38.485 13.295 47.115 14.195 ;
        RECT 48.785 14.175 49.730 14.270 ;
        RECT 56.470 14.175 57.415 14.270 ;
        RECT 48.785 13.275 57.415 14.175 ;
        RECT 59.095 14.155 60.040 14.250 ;
        RECT 66.780 14.155 67.725 14.250 ;
        RECT 59.095 13.255 67.725 14.155 ;
        RECT 69.465 14.145 70.410 14.240 ;
        RECT 77.150 14.145 78.095 14.240 ;
        RECT 69.465 13.245 78.095 14.145 ;
        RECT 79.775 14.125 80.720 14.220 ;
        RECT 87.460 14.125 88.405 14.220 ;
        RECT 79.775 13.225 88.405 14.125 ;
      LAYER li1 ;
        RECT 7.340 36.160 15.980 36.330 ;
        RECT 7.425 34.735 7.695 35.895 ;
        RECT 7.895 34.965 8.225 36.160 ;
        RECT 9.420 35.035 9.750 35.670 ;
        RECT 8.395 34.865 9.750 35.035 ;
        RECT 9.950 35.375 10.200 35.670 ;
        RECT 10.420 35.545 10.750 36.160 ;
        RECT 10.940 35.375 11.270 35.670 ;
        RECT 9.950 35.205 11.270 35.375 ;
        RECT 11.445 35.220 11.775 36.160 ;
        RECT 9.950 34.880 10.200 35.205 ;
        RECT 12.410 35.035 12.835 35.670 ;
        RECT 8.395 34.795 8.565 34.865 ;
        RECT 7.425 34.045 7.595 34.735 ;
        RECT 7.875 34.625 8.565 34.795 ;
        RECT 7.875 34.545 8.045 34.625 ;
        RECT 7.765 34.215 8.045 34.545 ;
        RECT 8.905 34.490 9.135 34.695 ;
        RECT 9.420 34.660 9.750 34.865 ;
        RECT 10.370 34.865 12.835 35.035 ;
        RECT 13.005 35.170 13.290 35.670 ;
        RECT 13.460 35.415 14.165 36.160 ;
        RECT 14.340 35.170 14.660 35.745 ;
        RECT 13.005 35.000 14.660 35.170 ;
        RECT 14.330 34.865 14.660 35.000 ;
        RECT 10.370 34.710 10.540 34.865 ;
        RECT 9.920 34.540 10.540 34.710 ;
        RECT 12.665 34.830 12.835 34.865 ;
        RECT 9.920 34.490 10.090 34.540 ;
        RECT 7.425 33.265 7.705 34.045 ;
        RECT 7.875 33.665 8.045 34.215 ;
        RECT 8.225 34.135 8.555 34.455 ;
        RECT 8.905 34.175 9.455 34.490 ;
        RECT 9.665 34.175 10.090 34.490 ;
        RECT 8.385 34.005 8.555 34.135 ;
        RECT 10.640 34.005 10.970 34.370 ;
        RECT 11.180 34.175 11.535 34.695 ;
        RECT 12.265 34.490 12.495 34.695 ;
        RECT 12.665 34.660 13.890 34.830 ;
        RECT 15.095 34.735 15.425 36.160 ;
        RECT 17.750 36.000 26.390 36.170 ;
        RECT 28.050 36.140 36.690 36.310 ;
        RECT 38.360 36.170 47.000 36.340 ;
        RECT 11.720 34.020 12.050 34.370 ;
        RECT 12.265 34.190 12.980 34.490 ;
        RECT 13.150 34.235 13.550 34.490 ;
        RECT 13.150 34.020 13.320 34.235 ;
        RECT 13.720 34.065 13.890 34.660 ;
        RECT 14.140 34.235 14.810 34.695 ;
        RECT 15.050 34.065 15.380 34.465 ;
        RECT 11.720 34.005 13.320 34.020 ;
        RECT 8.385 33.850 13.320 34.005 ;
        RECT 13.490 33.895 15.380 34.065 ;
        RECT 15.625 34.045 15.880 35.895 ;
        RECT 8.385 33.835 12.050 33.850 ;
        RECT 13.490 33.680 13.660 33.895 ;
        RECT 7.875 33.495 9.610 33.665 ;
        RECT 7.965 33.000 8.320 33.325 ;
        RECT 9.280 33.270 9.610 33.495 ;
        RECT 9.820 33.495 11.250 33.665 ;
        RECT 9.820 33.335 10.230 33.495 ;
        RECT 10.920 33.335 11.250 33.495 ;
        RECT 10.410 33.000 10.740 33.325 ;
        RECT 11.420 33.000 11.895 33.625 ;
        RECT 12.385 33.510 13.660 33.680 ;
        RECT 13.830 33.555 14.930 33.725 ;
        RECT 12.385 33.350 12.715 33.510 ;
        RECT 13.830 33.340 14.000 33.555 ;
        RECT 14.600 33.395 14.930 33.555 ;
        RECT 12.895 33.170 14.000 33.340 ;
        RECT 14.170 33.000 14.420 33.385 ;
        RECT 15.120 33.000 15.370 33.685 ;
        RECT 15.550 33.265 15.880 34.045 ;
        RECT 17.835 34.575 18.105 35.735 ;
        RECT 18.305 34.805 18.635 36.000 ;
        RECT 19.830 34.875 20.160 35.510 ;
        RECT 18.805 34.705 20.160 34.875 ;
        RECT 20.360 35.215 20.610 35.510 ;
        RECT 20.830 35.385 21.160 36.000 ;
        RECT 21.350 35.215 21.680 35.510 ;
        RECT 20.360 35.045 21.680 35.215 ;
        RECT 21.855 35.060 22.185 36.000 ;
        RECT 20.360 34.720 20.610 35.045 ;
        RECT 22.820 34.875 23.245 35.510 ;
        RECT 18.805 34.635 18.975 34.705 ;
        RECT 17.835 33.885 18.005 34.575 ;
        RECT 18.285 34.465 18.975 34.635 ;
        RECT 18.285 34.385 18.455 34.465 ;
        RECT 18.175 34.055 18.455 34.385 ;
        RECT 19.315 34.330 19.545 34.535 ;
        RECT 19.830 34.500 20.160 34.705 ;
        RECT 20.780 34.705 23.245 34.875 ;
        RECT 23.415 35.010 23.700 35.510 ;
        RECT 23.870 35.255 24.575 36.000 ;
        RECT 24.750 35.010 25.070 35.585 ;
        RECT 23.415 34.840 25.070 35.010 ;
        RECT 24.740 34.705 25.070 34.840 ;
        RECT 20.780 34.550 20.950 34.705 ;
        RECT 20.330 34.380 20.950 34.550 ;
        RECT 23.075 34.670 23.245 34.705 ;
        RECT 20.330 34.330 20.500 34.380 ;
        RECT 17.835 33.105 18.115 33.885 ;
        RECT 18.285 33.505 18.455 34.055 ;
        RECT 18.635 33.975 18.965 34.295 ;
        RECT 19.315 34.015 19.865 34.330 ;
        RECT 20.075 34.015 20.500 34.330 ;
        RECT 18.795 33.845 18.965 33.975 ;
        RECT 21.050 33.845 21.380 34.210 ;
        RECT 21.590 34.015 21.945 34.535 ;
        RECT 22.675 34.330 22.905 34.535 ;
        RECT 23.075 34.500 24.300 34.670 ;
        RECT 25.505 34.575 25.835 36.000 ;
        RECT 22.130 33.860 22.460 34.210 ;
        RECT 22.675 34.030 23.390 34.330 ;
        RECT 23.560 34.075 23.960 34.330 ;
        RECT 23.560 33.860 23.730 34.075 ;
        RECT 24.130 33.905 24.300 34.500 ;
        RECT 24.550 34.075 25.220 34.535 ;
        RECT 25.460 33.905 25.790 34.305 ;
        RECT 22.130 33.845 23.730 33.860 ;
        RECT 18.795 33.690 23.730 33.845 ;
        RECT 23.900 33.735 25.790 33.905 ;
        RECT 26.035 33.885 26.290 35.735 ;
        RECT 18.795 33.675 22.460 33.690 ;
        RECT 23.900 33.520 24.070 33.735 ;
        RECT 18.285 33.335 20.020 33.505 ;
        RECT 7.340 32.830 15.980 33.000 ;
        RECT 18.375 32.840 18.730 33.165 ;
        RECT 19.690 33.110 20.020 33.335 ;
        RECT 20.230 33.335 21.660 33.505 ;
        RECT 20.230 33.175 20.640 33.335 ;
        RECT 21.330 33.175 21.660 33.335 ;
        RECT 20.820 32.840 21.150 33.165 ;
        RECT 21.830 32.840 22.305 33.465 ;
        RECT 22.795 33.350 24.070 33.520 ;
        RECT 24.240 33.395 25.340 33.565 ;
        RECT 22.795 33.190 23.125 33.350 ;
        RECT 24.240 33.180 24.410 33.395 ;
        RECT 25.010 33.235 25.340 33.395 ;
        RECT 23.305 33.010 24.410 33.180 ;
        RECT 24.580 32.840 24.830 33.225 ;
        RECT 25.530 32.840 25.780 33.525 ;
        RECT 25.960 33.105 26.290 33.885 ;
        RECT 28.135 34.715 28.405 35.875 ;
        RECT 28.605 34.945 28.935 36.140 ;
        RECT 30.130 35.015 30.460 35.650 ;
        RECT 29.105 34.845 30.460 35.015 ;
        RECT 30.660 35.355 30.910 35.650 ;
        RECT 31.130 35.525 31.460 36.140 ;
        RECT 31.650 35.355 31.980 35.650 ;
        RECT 30.660 35.185 31.980 35.355 ;
        RECT 32.155 35.200 32.485 36.140 ;
        RECT 30.660 34.860 30.910 35.185 ;
        RECT 33.120 35.015 33.545 35.650 ;
        RECT 29.105 34.775 29.275 34.845 ;
        RECT 28.135 34.025 28.305 34.715 ;
        RECT 28.585 34.605 29.275 34.775 ;
        RECT 28.585 34.525 28.755 34.605 ;
        RECT 28.475 34.195 28.755 34.525 ;
        RECT 29.615 34.470 29.845 34.675 ;
        RECT 30.130 34.640 30.460 34.845 ;
        RECT 31.080 34.845 33.545 35.015 ;
        RECT 33.715 35.150 34.000 35.650 ;
        RECT 34.170 35.395 34.875 36.140 ;
        RECT 35.050 35.150 35.370 35.725 ;
        RECT 33.715 34.980 35.370 35.150 ;
        RECT 35.040 34.845 35.370 34.980 ;
        RECT 31.080 34.690 31.250 34.845 ;
        RECT 30.630 34.520 31.250 34.690 ;
        RECT 33.375 34.810 33.545 34.845 ;
        RECT 30.630 34.470 30.800 34.520 ;
        RECT 28.135 33.245 28.415 34.025 ;
        RECT 28.585 33.645 28.755 34.195 ;
        RECT 28.935 34.115 29.265 34.435 ;
        RECT 29.615 34.155 30.165 34.470 ;
        RECT 30.375 34.155 30.800 34.470 ;
        RECT 29.095 33.985 29.265 34.115 ;
        RECT 31.350 33.985 31.680 34.350 ;
        RECT 31.890 34.155 32.245 34.675 ;
        RECT 32.975 34.470 33.205 34.675 ;
        RECT 33.375 34.640 34.600 34.810 ;
        RECT 35.805 34.715 36.135 36.140 ;
        RECT 32.430 34.000 32.760 34.350 ;
        RECT 32.975 34.170 33.690 34.470 ;
        RECT 33.860 34.215 34.260 34.470 ;
        RECT 33.860 34.000 34.030 34.215 ;
        RECT 34.430 34.045 34.600 34.640 ;
        RECT 34.850 34.215 35.520 34.675 ;
        RECT 35.760 34.045 36.090 34.445 ;
        RECT 32.430 33.985 34.030 34.000 ;
        RECT 29.095 33.830 34.030 33.985 ;
        RECT 34.200 33.875 36.090 34.045 ;
        RECT 36.335 34.025 36.590 35.875 ;
        RECT 29.095 33.815 32.760 33.830 ;
        RECT 34.200 33.660 34.370 33.875 ;
        RECT 28.585 33.475 30.320 33.645 ;
        RECT 28.675 32.980 29.030 33.305 ;
        RECT 29.990 33.250 30.320 33.475 ;
        RECT 30.530 33.475 31.960 33.645 ;
        RECT 30.530 33.315 30.940 33.475 ;
        RECT 31.630 33.315 31.960 33.475 ;
        RECT 31.120 32.980 31.450 33.305 ;
        RECT 32.130 32.980 32.605 33.605 ;
        RECT 33.095 33.490 34.370 33.660 ;
        RECT 34.540 33.535 35.640 33.705 ;
        RECT 33.095 33.330 33.425 33.490 ;
        RECT 34.540 33.320 34.710 33.535 ;
        RECT 35.310 33.375 35.640 33.535 ;
        RECT 33.605 33.150 34.710 33.320 ;
        RECT 34.880 32.980 35.130 33.365 ;
        RECT 35.830 32.980 36.080 33.665 ;
        RECT 36.260 33.245 36.590 34.025 ;
        RECT 38.445 34.745 38.715 35.905 ;
        RECT 38.915 34.975 39.245 36.170 ;
        RECT 40.440 35.045 40.770 35.680 ;
        RECT 39.415 34.875 40.770 35.045 ;
        RECT 40.970 35.385 41.220 35.680 ;
        RECT 41.440 35.555 41.770 36.170 ;
        RECT 41.960 35.385 42.290 35.680 ;
        RECT 40.970 35.215 42.290 35.385 ;
        RECT 42.465 35.230 42.795 36.170 ;
        RECT 40.970 34.890 41.220 35.215 ;
        RECT 43.430 35.045 43.855 35.680 ;
        RECT 39.415 34.805 39.585 34.875 ;
        RECT 38.445 34.055 38.615 34.745 ;
        RECT 38.895 34.635 39.585 34.805 ;
        RECT 38.895 34.555 39.065 34.635 ;
        RECT 38.785 34.225 39.065 34.555 ;
        RECT 39.925 34.500 40.155 34.705 ;
        RECT 40.440 34.670 40.770 34.875 ;
        RECT 41.390 34.875 43.855 35.045 ;
        RECT 44.025 35.180 44.310 35.680 ;
        RECT 44.480 35.425 45.185 36.170 ;
        RECT 45.360 35.180 45.680 35.755 ;
        RECT 44.025 35.010 45.680 35.180 ;
        RECT 45.350 34.875 45.680 35.010 ;
        RECT 41.390 34.720 41.560 34.875 ;
        RECT 40.940 34.550 41.560 34.720 ;
        RECT 43.685 34.840 43.855 34.875 ;
        RECT 40.940 34.500 41.110 34.550 ;
        RECT 38.445 33.275 38.725 34.055 ;
        RECT 38.895 33.675 39.065 34.225 ;
        RECT 39.245 34.145 39.575 34.465 ;
        RECT 39.925 34.185 40.475 34.500 ;
        RECT 40.685 34.185 41.110 34.500 ;
        RECT 39.405 34.015 39.575 34.145 ;
        RECT 41.660 34.015 41.990 34.380 ;
        RECT 42.200 34.185 42.555 34.705 ;
        RECT 43.285 34.500 43.515 34.705 ;
        RECT 43.685 34.670 44.910 34.840 ;
        RECT 46.115 34.745 46.445 36.170 ;
        RECT 42.740 34.030 43.070 34.380 ;
        RECT 43.285 34.200 44.000 34.500 ;
        RECT 44.170 34.245 44.570 34.500 ;
        RECT 44.170 34.030 44.340 34.245 ;
        RECT 44.740 34.075 44.910 34.670 ;
        RECT 45.160 34.245 45.830 34.705 ;
        RECT 46.070 34.075 46.400 34.475 ;
        RECT 42.740 34.015 44.340 34.030 ;
        RECT 39.405 33.860 44.340 34.015 ;
        RECT 44.510 33.905 46.400 34.075 ;
        RECT 46.645 34.055 46.900 35.905 ;
        RECT 39.405 33.845 43.070 33.860 ;
        RECT 44.510 33.690 44.680 33.905 ;
        RECT 38.895 33.505 40.630 33.675 ;
        RECT 38.985 33.010 39.340 33.335 ;
        RECT 40.300 33.280 40.630 33.505 ;
        RECT 40.840 33.505 42.270 33.675 ;
        RECT 40.840 33.345 41.250 33.505 ;
        RECT 41.940 33.345 42.270 33.505 ;
        RECT 41.430 33.010 41.760 33.335 ;
        RECT 42.440 33.010 42.915 33.635 ;
        RECT 43.405 33.520 44.680 33.690 ;
        RECT 44.850 33.565 45.950 33.735 ;
        RECT 43.405 33.360 43.735 33.520 ;
        RECT 44.850 33.350 45.020 33.565 ;
        RECT 45.620 33.405 45.950 33.565 ;
        RECT 43.915 33.180 45.020 33.350 ;
        RECT 45.190 33.010 45.440 33.395 ;
        RECT 46.140 33.010 46.390 33.695 ;
        RECT 46.570 33.275 46.900 34.055 ;
        RECT 17.750 32.670 26.390 32.840 ;
        RECT 28.050 32.810 36.690 32.980 ;
        RECT 38.360 32.840 47.000 33.010 ;
        RECT 46.060 32.010 46.230 32.140 ;
        RECT 49.390 32.035 49.560 32.140 ;
        RECT 46.060 31.760 47.275 32.010 ;
        RECT 46.060 31.070 46.230 31.760 ;
        RECT 47.445 31.705 47.925 32.035 ;
        RECT 48.095 31.705 49.560 32.035 ;
        RECT 46.495 31.535 47.275 31.580 ;
        RECT 46.495 31.250 49.125 31.535 ;
        RECT 46.060 30.820 47.275 31.070 ;
        RECT 49.390 31.055 49.560 31.705 ;
        RECT 46.060 30.700 46.230 30.820 ;
        RECT 47.965 30.805 49.560 31.055 ;
        RECT 49.390 30.700 49.560 30.805 ;
        RECT 84.590 30.485 88.910 30.655 ;
        RECT 7.260 30.230 15.900 30.400 ;
        RECT 17.580 30.310 26.220 30.480 ;
        RECT 7.360 29.185 7.690 29.965 ;
        RECT 7.870 29.545 8.120 30.230 ;
        RECT 8.820 29.845 9.070 30.230 ;
        RECT 9.240 29.890 10.345 30.060 ;
        RECT 8.310 29.675 8.640 29.835 ;
        RECT 9.240 29.675 9.410 29.890 ;
        RECT 10.525 29.720 10.855 29.880 ;
        RECT 8.310 29.505 9.410 29.675 ;
        RECT 9.580 29.550 10.855 29.720 ;
        RECT 11.345 29.605 11.820 30.230 ;
        RECT 12.500 29.905 12.830 30.230 ;
        RECT 11.990 29.735 12.320 29.895 ;
        RECT 13.010 29.735 13.420 29.895 ;
        RECT 11.990 29.565 13.420 29.735 ;
        RECT 13.630 29.735 13.960 29.960 ;
        RECT 14.920 29.905 15.275 30.230 ;
        RECT 13.630 29.565 15.365 29.735 ;
        RECT 9.580 29.335 9.750 29.550 ;
        RECT 11.190 29.380 14.855 29.395 ;
        RECT 7.360 27.335 7.615 29.185 ;
        RECT 7.860 29.165 9.750 29.335 ;
        RECT 9.920 29.225 14.855 29.380 ;
        RECT 9.920 29.210 11.520 29.225 ;
        RECT 7.860 28.765 8.190 29.165 ;
        RECT 8.430 28.535 9.100 28.995 ;
        RECT 9.350 28.570 9.520 29.165 ;
        RECT 9.920 28.995 10.090 29.210 ;
        RECT 9.690 28.740 10.090 28.995 ;
        RECT 10.260 28.740 10.975 29.040 ;
        RECT 11.190 28.860 11.520 29.210 ;
        RECT 7.815 27.070 8.145 28.495 ;
        RECT 9.350 28.400 10.575 28.570 ;
        RECT 10.745 28.535 10.975 28.740 ;
        RECT 11.705 28.535 12.060 29.055 ;
        RECT 12.270 28.860 12.600 29.225 ;
        RECT 14.685 29.095 14.855 29.225 ;
        RECT 13.150 28.740 13.575 29.055 ;
        RECT 13.785 28.740 14.335 29.055 ;
        RECT 14.685 28.775 15.015 29.095 ;
        RECT 15.195 29.015 15.365 29.565 ;
        RECT 15.535 29.185 15.815 29.965 ;
        RECT 13.150 28.690 13.320 28.740 ;
        RECT 10.405 28.365 10.575 28.400 ;
        RECT 12.700 28.520 13.320 28.690 ;
        RECT 12.700 28.365 12.870 28.520 ;
        RECT 8.580 28.230 8.910 28.365 ;
        RECT 8.580 28.060 10.235 28.230 ;
        RECT 8.580 27.485 8.900 28.060 ;
        RECT 9.075 27.070 9.780 27.815 ;
        RECT 9.950 27.560 10.235 28.060 ;
        RECT 10.405 28.195 12.870 28.365 ;
        RECT 13.490 28.365 13.820 28.570 ;
        RECT 14.105 28.535 14.335 28.740 ;
        RECT 15.195 28.685 15.475 29.015 ;
        RECT 15.195 28.605 15.365 28.685 ;
        RECT 14.675 28.435 15.365 28.605 ;
        RECT 15.645 28.495 15.815 29.185 ;
        RECT 14.675 28.365 14.845 28.435 ;
        RECT 10.405 27.560 10.830 28.195 ;
        RECT 13.040 28.025 13.290 28.350 ;
        RECT 11.465 27.070 11.795 28.010 ;
        RECT 11.970 27.855 13.290 28.025 ;
        RECT 11.970 27.560 12.300 27.855 ;
        RECT 12.490 27.070 12.820 27.685 ;
        RECT 13.040 27.560 13.290 27.855 ;
        RECT 13.490 28.195 14.845 28.365 ;
        RECT 13.490 27.560 13.820 28.195 ;
        RECT 15.015 27.070 15.345 28.265 ;
        RECT 15.545 27.335 15.815 28.495 ;
        RECT 17.680 29.265 18.010 30.045 ;
        RECT 18.190 29.625 18.440 30.310 ;
        RECT 19.140 29.925 19.390 30.310 ;
        RECT 19.560 29.970 20.665 30.140 ;
        RECT 18.630 29.755 18.960 29.915 ;
        RECT 19.560 29.755 19.730 29.970 ;
        RECT 20.845 29.800 21.175 29.960 ;
        RECT 18.630 29.585 19.730 29.755 ;
        RECT 19.900 29.630 21.175 29.800 ;
        RECT 21.665 29.685 22.140 30.310 ;
        RECT 22.820 29.985 23.150 30.310 ;
        RECT 22.310 29.815 22.640 29.975 ;
        RECT 23.330 29.815 23.740 29.975 ;
        RECT 22.310 29.645 23.740 29.815 ;
        RECT 23.950 29.815 24.280 30.040 ;
        RECT 25.240 29.985 25.595 30.310 ;
        RECT 27.890 30.150 36.530 30.320 ;
        RECT 23.950 29.645 25.685 29.815 ;
        RECT 19.900 29.415 20.070 29.630 ;
        RECT 21.510 29.460 25.175 29.475 ;
        RECT 17.680 27.415 17.935 29.265 ;
        RECT 18.180 29.245 20.070 29.415 ;
        RECT 20.240 29.305 25.175 29.460 ;
        RECT 20.240 29.290 21.840 29.305 ;
        RECT 18.180 28.845 18.510 29.245 ;
        RECT 18.750 28.615 19.420 29.075 ;
        RECT 19.670 28.650 19.840 29.245 ;
        RECT 20.240 29.075 20.410 29.290 ;
        RECT 20.010 28.820 20.410 29.075 ;
        RECT 20.580 28.820 21.295 29.120 ;
        RECT 21.510 28.940 21.840 29.290 ;
        RECT 18.135 27.150 18.465 28.575 ;
        RECT 19.670 28.480 20.895 28.650 ;
        RECT 21.065 28.615 21.295 28.820 ;
        RECT 22.025 28.615 22.380 29.135 ;
        RECT 22.590 28.940 22.920 29.305 ;
        RECT 25.005 29.175 25.175 29.305 ;
        RECT 23.470 28.820 23.895 29.135 ;
        RECT 24.105 28.820 24.655 29.135 ;
        RECT 25.005 28.855 25.335 29.175 ;
        RECT 25.515 29.095 25.685 29.645 ;
        RECT 25.855 29.265 26.135 30.045 ;
        RECT 23.470 28.770 23.640 28.820 ;
        RECT 20.725 28.445 20.895 28.480 ;
        RECT 23.020 28.600 23.640 28.770 ;
        RECT 23.020 28.445 23.190 28.600 ;
        RECT 18.900 28.310 19.230 28.445 ;
        RECT 18.900 28.140 20.555 28.310 ;
        RECT 18.900 27.565 19.220 28.140 ;
        RECT 19.395 27.150 20.100 27.895 ;
        RECT 20.270 27.640 20.555 28.140 ;
        RECT 20.725 28.275 23.190 28.445 ;
        RECT 23.810 28.445 24.140 28.650 ;
        RECT 24.425 28.615 24.655 28.820 ;
        RECT 25.515 28.765 25.795 29.095 ;
        RECT 25.515 28.685 25.685 28.765 ;
        RECT 24.995 28.515 25.685 28.685 ;
        RECT 25.965 28.575 26.135 29.265 ;
        RECT 24.995 28.445 25.165 28.515 ;
        RECT 20.725 27.640 21.150 28.275 ;
        RECT 23.360 28.105 23.610 28.430 ;
        RECT 21.785 27.150 22.115 28.090 ;
        RECT 22.290 27.935 23.610 28.105 ;
        RECT 22.290 27.640 22.620 27.935 ;
        RECT 22.810 27.150 23.140 27.765 ;
        RECT 23.360 27.640 23.610 27.935 ;
        RECT 23.810 28.275 25.165 28.445 ;
        RECT 23.810 27.640 24.140 28.275 ;
        RECT 25.335 27.150 25.665 28.345 ;
        RECT 25.865 27.415 26.135 28.575 ;
        RECT 27.990 29.105 28.320 29.885 ;
        RECT 28.500 29.465 28.750 30.150 ;
        RECT 29.450 29.765 29.700 30.150 ;
        RECT 29.870 29.810 30.975 29.980 ;
        RECT 28.940 29.595 29.270 29.755 ;
        RECT 29.870 29.595 30.040 29.810 ;
        RECT 31.155 29.640 31.485 29.800 ;
        RECT 28.940 29.425 30.040 29.595 ;
        RECT 30.210 29.470 31.485 29.640 ;
        RECT 31.975 29.525 32.450 30.150 ;
        RECT 33.130 29.825 33.460 30.150 ;
        RECT 32.620 29.655 32.950 29.815 ;
        RECT 33.640 29.655 34.050 29.815 ;
        RECT 32.620 29.485 34.050 29.655 ;
        RECT 34.260 29.655 34.590 29.880 ;
        RECT 35.550 29.825 35.905 30.150 ;
        RECT 38.260 30.120 46.900 30.290 ;
        RECT 34.260 29.485 35.995 29.655 ;
        RECT 30.210 29.255 30.380 29.470 ;
        RECT 31.820 29.300 35.485 29.315 ;
        RECT 27.990 27.255 28.245 29.105 ;
        RECT 28.490 29.085 30.380 29.255 ;
        RECT 30.550 29.145 35.485 29.300 ;
        RECT 30.550 29.130 32.150 29.145 ;
        RECT 28.490 28.685 28.820 29.085 ;
        RECT 29.060 28.455 29.730 28.915 ;
        RECT 29.980 28.490 30.150 29.085 ;
        RECT 30.550 28.915 30.720 29.130 ;
        RECT 30.320 28.660 30.720 28.915 ;
        RECT 30.890 28.660 31.605 28.960 ;
        RECT 31.820 28.780 32.150 29.130 ;
        RECT 7.260 26.900 15.900 27.070 ;
        RECT 17.580 26.980 26.220 27.150 ;
        RECT 28.445 26.990 28.775 28.415 ;
        RECT 29.980 28.320 31.205 28.490 ;
        RECT 31.375 28.455 31.605 28.660 ;
        RECT 32.335 28.455 32.690 28.975 ;
        RECT 32.900 28.780 33.230 29.145 ;
        RECT 35.315 29.015 35.485 29.145 ;
        RECT 33.780 28.660 34.205 28.975 ;
        RECT 34.415 28.660 34.965 28.975 ;
        RECT 35.315 28.695 35.645 29.015 ;
        RECT 35.825 28.935 35.995 29.485 ;
        RECT 36.165 29.105 36.445 29.885 ;
        RECT 33.780 28.610 33.950 28.660 ;
        RECT 31.035 28.285 31.205 28.320 ;
        RECT 33.330 28.440 33.950 28.610 ;
        RECT 33.330 28.285 33.500 28.440 ;
        RECT 29.210 28.150 29.540 28.285 ;
        RECT 29.210 27.980 30.865 28.150 ;
        RECT 29.210 27.405 29.530 27.980 ;
        RECT 29.705 26.990 30.410 27.735 ;
        RECT 30.580 27.480 30.865 27.980 ;
        RECT 31.035 28.115 33.500 28.285 ;
        RECT 34.120 28.285 34.450 28.490 ;
        RECT 34.735 28.455 34.965 28.660 ;
        RECT 35.825 28.605 36.105 28.935 ;
        RECT 35.825 28.525 35.995 28.605 ;
        RECT 35.305 28.355 35.995 28.525 ;
        RECT 36.275 28.415 36.445 29.105 ;
        RECT 35.305 28.285 35.475 28.355 ;
        RECT 31.035 27.480 31.460 28.115 ;
        RECT 33.670 27.945 33.920 28.270 ;
        RECT 32.095 26.990 32.425 27.930 ;
        RECT 32.600 27.775 33.920 27.945 ;
        RECT 32.600 27.480 32.930 27.775 ;
        RECT 33.120 26.990 33.450 27.605 ;
        RECT 33.670 27.480 33.920 27.775 ;
        RECT 34.120 28.115 35.475 28.285 ;
        RECT 34.120 27.480 34.450 28.115 ;
        RECT 35.645 26.990 35.975 28.185 ;
        RECT 36.175 27.255 36.445 28.415 ;
        RECT 38.360 29.075 38.690 29.855 ;
        RECT 38.870 29.435 39.120 30.120 ;
        RECT 39.820 29.735 40.070 30.120 ;
        RECT 40.240 29.780 41.345 29.950 ;
        RECT 39.310 29.565 39.640 29.725 ;
        RECT 40.240 29.565 40.410 29.780 ;
        RECT 41.525 29.610 41.855 29.770 ;
        RECT 39.310 29.395 40.410 29.565 ;
        RECT 40.580 29.440 41.855 29.610 ;
        RECT 42.345 29.495 42.820 30.120 ;
        RECT 43.500 29.795 43.830 30.120 ;
        RECT 42.990 29.625 43.320 29.785 ;
        RECT 44.010 29.625 44.420 29.785 ;
        RECT 42.990 29.455 44.420 29.625 ;
        RECT 44.630 29.625 44.960 29.850 ;
        RECT 45.920 29.795 46.275 30.120 ;
        RECT 44.630 29.455 46.365 29.625 ;
        RECT 40.580 29.225 40.750 29.440 ;
        RECT 42.190 29.270 45.855 29.285 ;
        RECT 38.360 27.225 38.615 29.075 ;
        RECT 38.860 29.055 40.750 29.225 ;
        RECT 40.920 29.115 45.855 29.270 ;
        RECT 40.920 29.100 42.520 29.115 ;
        RECT 38.860 28.655 39.190 29.055 ;
        RECT 39.430 28.425 40.100 28.885 ;
        RECT 40.350 28.460 40.520 29.055 ;
        RECT 40.920 28.885 41.090 29.100 ;
        RECT 40.690 28.630 41.090 28.885 ;
        RECT 41.260 28.630 41.975 28.930 ;
        RECT 42.190 28.750 42.520 29.100 ;
        RECT 27.890 26.820 36.530 26.990 ;
        RECT 38.815 26.960 39.145 28.385 ;
        RECT 40.350 28.290 41.575 28.460 ;
        RECT 41.745 28.425 41.975 28.630 ;
        RECT 42.705 28.425 43.060 28.945 ;
        RECT 43.270 28.750 43.600 29.115 ;
        RECT 45.685 28.985 45.855 29.115 ;
        RECT 44.150 28.630 44.575 28.945 ;
        RECT 44.785 28.630 45.335 28.945 ;
        RECT 45.685 28.665 46.015 28.985 ;
        RECT 46.195 28.905 46.365 29.455 ;
        RECT 46.535 29.075 46.815 29.855 ;
        RECT 44.150 28.580 44.320 28.630 ;
        RECT 41.405 28.255 41.575 28.290 ;
        RECT 43.700 28.410 44.320 28.580 ;
        RECT 43.700 28.255 43.870 28.410 ;
        RECT 39.580 28.120 39.910 28.255 ;
        RECT 39.580 27.950 41.235 28.120 ;
        RECT 39.580 27.375 39.900 27.950 ;
        RECT 40.075 26.960 40.780 27.705 ;
        RECT 40.950 27.450 41.235 27.950 ;
        RECT 41.405 28.085 43.870 28.255 ;
        RECT 44.490 28.255 44.820 28.460 ;
        RECT 45.105 28.425 45.335 28.630 ;
        RECT 46.195 28.575 46.475 28.905 ;
        RECT 46.195 28.495 46.365 28.575 ;
        RECT 45.675 28.325 46.365 28.495 ;
        RECT 46.645 28.385 46.815 29.075 ;
        RECT 45.675 28.255 45.845 28.325 ;
        RECT 41.405 27.450 41.830 28.085 ;
        RECT 44.040 27.915 44.290 28.240 ;
        RECT 42.465 26.960 42.795 27.900 ;
        RECT 42.970 27.745 44.290 27.915 ;
        RECT 42.970 27.450 43.300 27.745 ;
        RECT 43.490 26.960 43.820 27.575 ;
        RECT 44.040 27.450 44.290 27.745 ;
        RECT 44.490 28.085 45.845 28.255 ;
        RECT 44.490 27.450 44.820 28.085 ;
        RECT 46.015 26.960 46.345 28.155 ;
        RECT 46.545 27.225 46.815 28.385 ;
        RECT 84.705 29.470 85.035 29.940 ;
        RECT 85.240 29.640 85.570 30.485 ;
        RECT 85.740 30.145 87.715 30.315 ;
        RECT 85.740 29.470 85.910 30.145 ;
        RECT 84.705 29.300 85.910 29.470 ;
        RECT 84.705 29.190 85.035 29.300 ;
        RECT 84.705 28.370 84.875 29.190 ;
        RECT 86.655 29.130 86.985 29.975 ;
        RECT 85.095 28.590 85.425 29.020 ;
        RECT 85.595 28.960 86.985 29.130 ;
        RECT 84.705 27.780 85.035 28.370 ;
        RECT 85.215 27.920 85.425 28.370 ;
        RECT 85.595 28.260 85.765 28.960 ;
        RECT 87.545 28.890 87.715 30.145 ;
        RECT 87.885 29.060 88.215 30.485 ;
        RECT 88.385 29.060 88.825 30.220 ;
        RECT 85.935 28.460 86.275 28.790 ;
        RECT 85.595 28.090 85.935 28.260 ;
        RECT 85.215 27.325 85.595 27.920 ;
        RECT 85.765 27.880 85.935 28.090 ;
        RECT 86.105 28.220 86.275 28.460 ;
        RECT 86.475 28.420 86.865 28.790 ;
        RECT 87.045 28.220 87.375 28.790 ;
        RECT 87.545 28.560 87.945 28.890 ;
        RECT 88.115 28.540 88.485 28.870 ;
        RECT 88.115 28.390 88.285 28.540 ;
        RECT 86.105 28.050 87.375 28.220 ;
        RECT 87.545 28.220 88.285 28.390 ;
        RECT 88.655 28.370 88.825 29.060 ;
        RECT 87.545 27.880 87.715 28.220 ;
        RECT 85.765 27.630 87.715 27.880 ;
        RECT 87.885 27.325 88.215 28.050 ;
        RECT 88.455 27.590 88.825 28.370 ;
        RECT 84.590 27.155 88.910 27.325 ;
        RECT 38.260 26.790 46.900 26.960 ;
        RECT 40.490 22.175 41.930 22.345 ;
        RECT 40.610 21.130 40.860 22.175 ;
        RECT 41.040 21.130 41.370 21.910 ;
        RECT 41.550 21.130 41.800 22.175 ;
        RECT 40.595 19.015 40.845 20.440 ;
        RECT 41.040 19.280 41.325 21.130 ;
        RECT 41.495 20.480 41.825 20.960 ;
        RECT 41.495 19.015 41.825 20.310 ;
        RECT 40.490 18.845 41.930 19.015 ;
        RECT 7.490 16.345 16.130 16.515 ;
        RECT 7.575 14.920 7.845 16.080 ;
        RECT 8.045 15.150 8.375 16.345 ;
        RECT 9.570 15.220 9.900 15.855 ;
        RECT 8.545 15.050 9.900 15.220 ;
        RECT 10.100 15.560 10.350 15.855 ;
        RECT 10.570 15.730 10.900 16.345 ;
        RECT 11.090 15.560 11.420 15.855 ;
        RECT 10.100 15.390 11.420 15.560 ;
        RECT 11.595 15.405 11.925 16.345 ;
        RECT 10.100 15.065 10.350 15.390 ;
        RECT 12.560 15.220 12.985 15.855 ;
        RECT 8.545 14.980 8.715 15.050 ;
        RECT 7.575 14.230 7.745 14.920 ;
        RECT 8.025 14.810 8.715 14.980 ;
        RECT 8.025 14.730 8.195 14.810 ;
        RECT 7.915 14.400 8.195 14.730 ;
        RECT 9.055 14.675 9.285 14.880 ;
        RECT 9.570 14.845 9.900 15.050 ;
        RECT 10.520 15.050 12.985 15.220 ;
        RECT 13.155 15.355 13.440 15.855 ;
        RECT 13.610 15.600 14.315 16.345 ;
        RECT 14.490 15.355 14.810 15.930 ;
        RECT 13.155 15.185 14.810 15.355 ;
        RECT 14.480 15.050 14.810 15.185 ;
        RECT 10.520 14.895 10.690 15.050 ;
        RECT 10.070 14.725 10.690 14.895 ;
        RECT 12.815 15.015 12.985 15.050 ;
        RECT 10.070 14.675 10.240 14.725 ;
        RECT 7.575 14.110 7.855 14.230 ;
        RECT 7.575 13.940 7.645 14.110 ;
        RECT 7.815 13.940 7.855 14.110 ;
        RECT 7.575 13.740 7.855 13.940 ;
        RECT 7.575 13.570 7.645 13.740 ;
        RECT 7.815 13.570 7.855 13.740 ;
        RECT 8.025 13.850 8.195 14.400 ;
        RECT 8.375 14.320 8.705 14.640 ;
        RECT 9.055 14.360 9.605 14.675 ;
        RECT 9.815 14.360 10.240 14.675 ;
        RECT 8.535 14.190 8.705 14.320 ;
        RECT 10.790 14.190 11.120 14.555 ;
        RECT 11.330 14.360 11.685 14.880 ;
        RECT 12.415 14.675 12.645 14.880 ;
        RECT 12.815 14.845 14.040 15.015 ;
        RECT 15.245 14.920 15.575 16.345 ;
        RECT 17.800 16.325 26.440 16.495 ;
        RECT 11.870 14.480 12.200 14.555 ;
        RECT 11.870 14.310 11.965 14.480 ;
        RECT 12.135 14.310 12.200 14.480 ;
        RECT 12.415 14.375 13.130 14.675 ;
        RECT 13.300 14.420 13.700 14.675 ;
        RECT 11.870 14.205 12.200 14.310 ;
        RECT 13.300 14.205 13.470 14.420 ;
        RECT 13.870 14.250 14.040 14.845 ;
        RECT 14.290 14.850 14.960 14.880 ;
        RECT 14.290 14.680 14.365 14.850 ;
        RECT 14.535 14.680 14.960 14.850 ;
        RECT 14.290 14.420 14.960 14.680 ;
        RECT 15.775 14.800 16.030 16.080 ;
        RECT 17.885 14.900 18.155 16.060 ;
        RECT 18.355 15.130 18.685 16.325 ;
        RECT 19.880 15.200 20.210 15.835 ;
        RECT 18.855 15.030 20.210 15.200 ;
        RECT 20.410 15.540 20.660 15.835 ;
        RECT 20.880 15.710 21.210 16.325 ;
        RECT 21.400 15.540 21.730 15.835 ;
        RECT 20.410 15.370 21.730 15.540 ;
        RECT 21.905 15.385 22.235 16.325 ;
        RECT 20.410 15.045 20.660 15.370 ;
        RECT 22.870 15.200 23.295 15.835 ;
        RECT 18.855 14.960 19.025 15.030 ;
        RECT 15.200 14.250 15.530 14.650 ;
        RECT 11.870 14.190 13.470 14.205 ;
        RECT 8.535 14.035 13.470 14.190 ;
        RECT 13.640 14.080 15.530 14.250 ;
        RECT 15.775 14.630 16.040 14.800 ;
        RECT 15.775 14.230 16.030 14.630 ;
        RECT 8.535 14.020 12.200 14.035 ;
        RECT 13.640 13.865 13.810 14.080 ;
        RECT 8.025 13.680 9.760 13.850 ;
        RECT 7.575 13.450 7.855 13.570 ;
        RECT 8.115 13.185 8.470 13.510 ;
        RECT 9.430 13.455 9.760 13.680 ;
        RECT 9.970 13.680 11.400 13.850 ;
        RECT 9.970 13.520 10.380 13.680 ;
        RECT 11.070 13.520 11.400 13.680 ;
        RECT 10.560 13.185 10.890 13.510 ;
        RECT 11.570 13.185 12.045 13.810 ;
        RECT 12.535 13.695 13.810 13.865 ;
        RECT 13.980 13.740 15.080 13.910 ;
        RECT 12.535 13.535 12.865 13.695 ;
        RECT 13.980 13.525 14.150 13.740 ;
        RECT 14.750 13.580 15.080 13.740 ;
        RECT 13.045 13.355 14.150 13.525 ;
        RECT 14.320 13.185 14.570 13.570 ;
        RECT 15.270 13.185 15.520 13.870 ;
        RECT 15.700 13.450 16.030 14.230 ;
        RECT 17.885 14.210 18.055 14.900 ;
        RECT 18.335 14.790 19.025 14.960 ;
        RECT 18.335 14.710 18.505 14.790 ;
        RECT 18.225 14.380 18.505 14.710 ;
        RECT 19.365 14.655 19.595 14.860 ;
        RECT 19.880 14.825 20.210 15.030 ;
        RECT 20.830 15.030 23.295 15.200 ;
        RECT 23.465 15.335 23.750 15.835 ;
        RECT 23.920 15.580 24.625 16.325 ;
        RECT 24.800 15.335 25.120 15.910 ;
        RECT 23.465 15.165 25.120 15.335 ;
        RECT 24.790 15.030 25.120 15.165 ;
        RECT 20.830 14.875 21.000 15.030 ;
        RECT 20.380 14.705 21.000 14.875 ;
        RECT 23.125 14.995 23.295 15.030 ;
        RECT 20.380 14.655 20.550 14.705 ;
        RECT 17.885 14.090 18.165 14.210 ;
        RECT 17.885 13.920 17.955 14.090 ;
        RECT 18.125 13.920 18.165 14.090 ;
        RECT 17.885 13.720 18.165 13.920 ;
        RECT 17.885 13.550 17.955 13.720 ;
        RECT 18.125 13.550 18.165 13.720 ;
        RECT 18.335 13.830 18.505 14.380 ;
        RECT 18.685 14.300 19.015 14.620 ;
        RECT 19.365 14.340 19.915 14.655 ;
        RECT 20.125 14.340 20.550 14.655 ;
        RECT 18.845 14.170 19.015 14.300 ;
        RECT 21.100 14.170 21.430 14.535 ;
        RECT 21.640 14.340 21.995 14.860 ;
        RECT 22.725 14.655 22.955 14.860 ;
        RECT 23.125 14.825 24.350 14.995 ;
        RECT 25.555 14.900 25.885 16.325 ;
        RECT 28.170 16.315 36.810 16.485 ;
        RECT 22.180 14.460 22.510 14.535 ;
        RECT 22.180 14.290 22.275 14.460 ;
        RECT 22.445 14.290 22.510 14.460 ;
        RECT 22.725 14.355 23.440 14.655 ;
        RECT 23.610 14.400 24.010 14.655 ;
        RECT 22.180 14.185 22.510 14.290 ;
        RECT 23.610 14.185 23.780 14.400 ;
        RECT 24.180 14.230 24.350 14.825 ;
        RECT 24.600 14.830 25.270 14.860 ;
        RECT 24.600 14.660 24.675 14.830 ;
        RECT 24.845 14.660 25.270 14.830 ;
        RECT 24.600 14.400 25.270 14.660 ;
        RECT 25.510 14.230 25.840 14.630 ;
        RECT 22.180 14.170 23.780 14.185 ;
        RECT 18.845 14.015 23.780 14.170 ;
        RECT 23.950 14.060 25.840 14.230 ;
        RECT 26.085 14.210 26.340 16.060 ;
        RECT 18.845 14.000 22.510 14.015 ;
        RECT 23.950 13.845 24.120 14.060 ;
        RECT 18.335 13.660 20.070 13.830 ;
        RECT 17.885 13.430 18.165 13.550 ;
        RECT 7.490 13.015 16.130 13.185 ;
        RECT 18.425 13.165 18.780 13.490 ;
        RECT 19.740 13.435 20.070 13.660 ;
        RECT 20.280 13.660 21.710 13.830 ;
        RECT 20.280 13.500 20.690 13.660 ;
        RECT 21.380 13.500 21.710 13.660 ;
        RECT 20.870 13.165 21.200 13.490 ;
        RECT 21.880 13.165 22.355 13.790 ;
        RECT 22.845 13.675 24.120 13.845 ;
        RECT 24.290 13.720 25.390 13.890 ;
        RECT 22.845 13.515 23.175 13.675 ;
        RECT 24.290 13.505 24.460 13.720 ;
        RECT 25.060 13.560 25.390 13.720 ;
        RECT 23.355 13.335 24.460 13.505 ;
        RECT 24.630 13.165 24.880 13.550 ;
        RECT 25.580 13.165 25.830 13.850 ;
        RECT 26.010 13.430 26.340 14.210 ;
        RECT 28.255 14.890 28.525 16.050 ;
        RECT 28.725 15.120 29.055 16.315 ;
        RECT 30.250 15.190 30.580 15.825 ;
        RECT 29.225 15.020 30.580 15.190 ;
        RECT 30.780 15.530 31.030 15.825 ;
        RECT 31.250 15.700 31.580 16.315 ;
        RECT 31.770 15.530 32.100 15.825 ;
        RECT 30.780 15.360 32.100 15.530 ;
        RECT 32.275 15.375 32.605 16.315 ;
        RECT 30.780 15.035 31.030 15.360 ;
        RECT 33.240 15.190 33.665 15.825 ;
        RECT 29.225 14.950 29.395 15.020 ;
        RECT 28.255 14.200 28.425 14.890 ;
        RECT 28.705 14.780 29.395 14.950 ;
        RECT 28.705 14.700 28.875 14.780 ;
        RECT 28.595 14.370 28.875 14.700 ;
        RECT 29.735 14.645 29.965 14.850 ;
        RECT 30.250 14.815 30.580 15.020 ;
        RECT 31.200 15.020 33.665 15.190 ;
        RECT 33.835 15.325 34.120 15.825 ;
        RECT 34.290 15.570 34.995 16.315 ;
        RECT 35.170 15.325 35.490 15.900 ;
        RECT 33.835 15.155 35.490 15.325 ;
        RECT 35.160 15.020 35.490 15.155 ;
        RECT 31.200 14.865 31.370 15.020 ;
        RECT 30.750 14.695 31.370 14.865 ;
        RECT 33.495 14.985 33.665 15.020 ;
        RECT 30.750 14.645 30.920 14.695 ;
        RECT 28.255 14.080 28.535 14.200 ;
        RECT 28.255 13.910 28.325 14.080 ;
        RECT 28.495 13.910 28.535 14.080 ;
        RECT 28.255 13.710 28.535 13.910 ;
        RECT 28.255 13.540 28.325 13.710 ;
        RECT 28.495 13.540 28.535 13.710 ;
        RECT 28.705 13.820 28.875 14.370 ;
        RECT 29.055 14.290 29.385 14.610 ;
        RECT 29.735 14.330 30.285 14.645 ;
        RECT 30.495 14.330 30.920 14.645 ;
        RECT 29.215 14.160 29.385 14.290 ;
        RECT 31.470 14.160 31.800 14.525 ;
        RECT 32.010 14.330 32.365 14.850 ;
        RECT 33.095 14.645 33.325 14.850 ;
        RECT 33.495 14.815 34.720 14.985 ;
        RECT 35.925 14.890 36.255 16.315 ;
        RECT 38.480 16.295 47.120 16.465 ;
        RECT 32.550 14.450 32.880 14.525 ;
        RECT 32.550 14.280 32.645 14.450 ;
        RECT 32.815 14.280 32.880 14.450 ;
        RECT 33.095 14.345 33.810 14.645 ;
        RECT 33.980 14.390 34.380 14.645 ;
        RECT 32.550 14.175 32.880 14.280 ;
        RECT 33.980 14.175 34.150 14.390 ;
        RECT 34.550 14.220 34.720 14.815 ;
        RECT 34.970 14.820 35.640 14.850 ;
        RECT 34.970 14.650 35.045 14.820 ;
        RECT 35.215 14.650 35.640 14.820 ;
        RECT 34.970 14.390 35.640 14.650 ;
        RECT 36.455 14.770 36.710 16.050 ;
        RECT 38.565 14.870 38.835 16.030 ;
        RECT 39.035 15.100 39.365 16.295 ;
        RECT 40.560 15.170 40.890 15.805 ;
        RECT 39.535 15.000 40.890 15.170 ;
        RECT 41.090 15.510 41.340 15.805 ;
        RECT 41.560 15.680 41.890 16.295 ;
        RECT 42.080 15.510 42.410 15.805 ;
        RECT 41.090 15.340 42.410 15.510 ;
        RECT 42.585 15.355 42.915 16.295 ;
        RECT 41.090 15.015 41.340 15.340 ;
        RECT 43.550 15.170 43.975 15.805 ;
        RECT 39.535 14.930 39.705 15.000 ;
        RECT 35.880 14.220 36.210 14.620 ;
        RECT 32.550 14.160 34.150 14.175 ;
        RECT 29.215 14.005 34.150 14.160 ;
        RECT 34.320 14.050 36.210 14.220 ;
        RECT 36.455 14.600 36.720 14.770 ;
        RECT 36.455 14.200 36.710 14.600 ;
        RECT 29.215 13.990 32.880 14.005 ;
        RECT 34.320 13.835 34.490 14.050 ;
        RECT 28.705 13.650 30.440 13.820 ;
        RECT 28.255 13.420 28.535 13.540 ;
        RECT 17.800 12.995 26.440 13.165 ;
        RECT 28.795 13.155 29.150 13.480 ;
        RECT 30.110 13.425 30.440 13.650 ;
        RECT 30.650 13.650 32.080 13.820 ;
        RECT 30.650 13.490 31.060 13.650 ;
        RECT 31.750 13.490 32.080 13.650 ;
        RECT 31.240 13.155 31.570 13.480 ;
        RECT 32.250 13.155 32.725 13.780 ;
        RECT 33.215 13.665 34.490 13.835 ;
        RECT 34.660 13.710 35.760 13.880 ;
        RECT 33.215 13.505 33.545 13.665 ;
        RECT 34.660 13.495 34.830 13.710 ;
        RECT 35.430 13.550 35.760 13.710 ;
        RECT 33.725 13.325 34.830 13.495 ;
        RECT 35.000 13.155 35.250 13.540 ;
        RECT 35.950 13.155 36.200 13.840 ;
        RECT 36.380 13.420 36.710 14.200 ;
        RECT 38.565 14.180 38.735 14.870 ;
        RECT 39.015 14.760 39.705 14.930 ;
        RECT 39.015 14.680 39.185 14.760 ;
        RECT 38.905 14.350 39.185 14.680 ;
        RECT 40.045 14.625 40.275 14.830 ;
        RECT 40.560 14.795 40.890 15.000 ;
        RECT 41.510 15.000 43.975 15.170 ;
        RECT 44.145 15.305 44.430 15.805 ;
        RECT 44.600 15.550 45.305 16.295 ;
        RECT 45.480 15.305 45.800 15.880 ;
        RECT 44.145 15.135 45.800 15.305 ;
        RECT 45.470 15.000 45.800 15.135 ;
        RECT 41.510 14.845 41.680 15.000 ;
        RECT 41.060 14.675 41.680 14.845 ;
        RECT 43.805 14.965 43.975 15.000 ;
        RECT 41.060 14.625 41.230 14.675 ;
        RECT 38.565 14.060 38.845 14.180 ;
        RECT 38.565 13.890 38.635 14.060 ;
        RECT 38.805 13.890 38.845 14.060 ;
        RECT 38.565 13.690 38.845 13.890 ;
        RECT 38.565 13.520 38.635 13.690 ;
        RECT 38.805 13.520 38.845 13.690 ;
        RECT 39.015 13.800 39.185 14.350 ;
        RECT 39.365 14.270 39.695 14.590 ;
        RECT 40.045 14.310 40.595 14.625 ;
        RECT 40.805 14.310 41.230 14.625 ;
        RECT 39.525 14.140 39.695 14.270 ;
        RECT 41.780 14.140 42.110 14.505 ;
        RECT 42.320 14.310 42.675 14.830 ;
        RECT 43.405 14.625 43.635 14.830 ;
        RECT 43.805 14.795 45.030 14.965 ;
        RECT 46.235 14.870 46.565 16.295 ;
        RECT 48.780 16.275 57.420 16.445 ;
        RECT 42.860 14.430 43.190 14.505 ;
        RECT 42.860 14.260 42.955 14.430 ;
        RECT 43.125 14.260 43.190 14.430 ;
        RECT 43.405 14.325 44.120 14.625 ;
        RECT 44.290 14.370 44.690 14.625 ;
        RECT 42.860 14.155 43.190 14.260 ;
        RECT 44.290 14.155 44.460 14.370 ;
        RECT 44.860 14.200 45.030 14.795 ;
        RECT 45.280 14.800 45.950 14.830 ;
        RECT 45.280 14.630 45.355 14.800 ;
        RECT 45.525 14.630 45.950 14.800 ;
        RECT 45.280 14.370 45.950 14.630 ;
        RECT 46.190 14.200 46.520 14.600 ;
        RECT 42.860 14.140 44.460 14.155 ;
        RECT 39.525 13.985 44.460 14.140 ;
        RECT 44.630 14.030 46.520 14.200 ;
        RECT 46.765 14.180 47.020 16.030 ;
        RECT 39.525 13.970 43.190 13.985 ;
        RECT 44.630 13.815 44.800 14.030 ;
        RECT 39.015 13.630 40.750 13.800 ;
        RECT 38.565 13.400 38.845 13.520 ;
        RECT 28.170 12.985 36.810 13.155 ;
        RECT 39.105 13.135 39.460 13.460 ;
        RECT 40.420 13.405 40.750 13.630 ;
        RECT 40.960 13.630 42.390 13.800 ;
        RECT 40.960 13.470 41.370 13.630 ;
        RECT 42.060 13.470 42.390 13.630 ;
        RECT 41.550 13.135 41.880 13.460 ;
        RECT 42.560 13.135 43.035 13.760 ;
        RECT 43.525 13.645 44.800 13.815 ;
        RECT 44.970 13.690 46.070 13.860 ;
        RECT 43.525 13.485 43.855 13.645 ;
        RECT 44.970 13.475 45.140 13.690 ;
        RECT 45.740 13.530 46.070 13.690 ;
        RECT 44.035 13.305 45.140 13.475 ;
        RECT 45.310 13.135 45.560 13.520 ;
        RECT 46.260 13.135 46.510 13.820 ;
        RECT 46.690 13.400 47.020 14.180 ;
        RECT 48.865 14.850 49.135 16.010 ;
        RECT 49.335 15.080 49.665 16.275 ;
        RECT 50.860 15.150 51.190 15.785 ;
        RECT 49.835 14.980 51.190 15.150 ;
        RECT 51.390 15.490 51.640 15.785 ;
        RECT 51.860 15.660 52.190 16.275 ;
        RECT 52.380 15.490 52.710 15.785 ;
        RECT 51.390 15.320 52.710 15.490 ;
        RECT 52.885 15.335 53.215 16.275 ;
        RECT 51.390 14.995 51.640 15.320 ;
        RECT 53.850 15.150 54.275 15.785 ;
        RECT 49.835 14.910 50.005 14.980 ;
        RECT 48.865 14.160 49.035 14.850 ;
        RECT 49.315 14.740 50.005 14.910 ;
        RECT 49.315 14.660 49.485 14.740 ;
        RECT 49.205 14.330 49.485 14.660 ;
        RECT 50.345 14.605 50.575 14.810 ;
        RECT 50.860 14.775 51.190 14.980 ;
        RECT 51.810 14.980 54.275 15.150 ;
        RECT 54.445 15.285 54.730 15.785 ;
        RECT 54.900 15.530 55.605 16.275 ;
        RECT 55.780 15.285 56.100 15.860 ;
        RECT 54.445 15.115 56.100 15.285 ;
        RECT 55.770 14.980 56.100 15.115 ;
        RECT 51.810 14.825 51.980 14.980 ;
        RECT 51.360 14.655 51.980 14.825 ;
        RECT 54.105 14.945 54.275 14.980 ;
        RECT 51.360 14.605 51.530 14.655 ;
        RECT 48.865 14.040 49.145 14.160 ;
        RECT 48.865 13.870 48.935 14.040 ;
        RECT 49.105 13.870 49.145 14.040 ;
        RECT 48.865 13.670 49.145 13.870 ;
        RECT 48.865 13.500 48.935 13.670 ;
        RECT 49.105 13.500 49.145 13.670 ;
        RECT 49.315 13.780 49.485 14.330 ;
        RECT 49.665 14.250 49.995 14.570 ;
        RECT 50.345 14.290 50.895 14.605 ;
        RECT 51.105 14.290 51.530 14.605 ;
        RECT 49.825 14.120 49.995 14.250 ;
        RECT 52.080 14.120 52.410 14.485 ;
        RECT 52.620 14.290 52.975 14.810 ;
        RECT 53.705 14.605 53.935 14.810 ;
        RECT 54.105 14.775 55.330 14.945 ;
        RECT 56.535 14.850 56.865 16.275 ;
        RECT 59.090 16.255 67.730 16.425 ;
        RECT 53.160 14.410 53.490 14.485 ;
        RECT 53.160 14.240 53.255 14.410 ;
        RECT 53.425 14.240 53.490 14.410 ;
        RECT 53.705 14.305 54.420 14.605 ;
        RECT 54.590 14.350 54.990 14.605 ;
        RECT 53.160 14.135 53.490 14.240 ;
        RECT 54.590 14.135 54.760 14.350 ;
        RECT 55.160 14.180 55.330 14.775 ;
        RECT 55.580 14.780 56.250 14.810 ;
        RECT 55.580 14.610 55.655 14.780 ;
        RECT 55.825 14.610 56.250 14.780 ;
        RECT 55.580 14.350 56.250 14.610 ;
        RECT 57.065 14.730 57.320 16.010 ;
        RECT 59.175 14.830 59.445 15.990 ;
        RECT 59.645 15.060 59.975 16.255 ;
        RECT 61.170 15.130 61.500 15.765 ;
        RECT 60.145 14.960 61.500 15.130 ;
        RECT 61.700 15.470 61.950 15.765 ;
        RECT 62.170 15.640 62.500 16.255 ;
        RECT 62.690 15.470 63.020 15.765 ;
        RECT 61.700 15.300 63.020 15.470 ;
        RECT 63.195 15.315 63.525 16.255 ;
        RECT 61.700 14.975 61.950 15.300 ;
        RECT 64.160 15.130 64.585 15.765 ;
        RECT 60.145 14.890 60.315 14.960 ;
        RECT 56.490 14.180 56.820 14.580 ;
        RECT 53.160 14.120 54.760 14.135 ;
        RECT 49.825 13.965 54.760 14.120 ;
        RECT 54.930 14.010 56.820 14.180 ;
        RECT 57.065 14.560 57.330 14.730 ;
        RECT 57.065 14.160 57.320 14.560 ;
        RECT 49.825 13.950 53.490 13.965 ;
        RECT 54.930 13.795 55.100 14.010 ;
        RECT 49.315 13.610 51.050 13.780 ;
        RECT 48.865 13.380 49.145 13.500 ;
        RECT 38.480 12.965 47.120 13.135 ;
        RECT 49.405 13.115 49.760 13.440 ;
        RECT 50.720 13.385 51.050 13.610 ;
        RECT 51.260 13.610 52.690 13.780 ;
        RECT 51.260 13.450 51.670 13.610 ;
        RECT 52.360 13.450 52.690 13.610 ;
        RECT 51.850 13.115 52.180 13.440 ;
        RECT 52.860 13.115 53.335 13.740 ;
        RECT 53.825 13.625 55.100 13.795 ;
        RECT 55.270 13.670 56.370 13.840 ;
        RECT 53.825 13.465 54.155 13.625 ;
        RECT 55.270 13.455 55.440 13.670 ;
        RECT 56.040 13.510 56.370 13.670 ;
        RECT 54.335 13.285 55.440 13.455 ;
        RECT 55.610 13.115 55.860 13.500 ;
        RECT 56.560 13.115 56.810 13.800 ;
        RECT 56.990 13.380 57.320 14.160 ;
        RECT 59.175 14.140 59.345 14.830 ;
        RECT 59.625 14.720 60.315 14.890 ;
        RECT 59.625 14.640 59.795 14.720 ;
        RECT 59.515 14.310 59.795 14.640 ;
        RECT 60.655 14.585 60.885 14.790 ;
        RECT 61.170 14.755 61.500 14.960 ;
        RECT 62.120 14.960 64.585 15.130 ;
        RECT 64.755 15.265 65.040 15.765 ;
        RECT 65.210 15.510 65.915 16.255 ;
        RECT 66.090 15.265 66.410 15.840 ;
        RECT 64.755 15.095 66.410 15.265 ;
        RECT 66.080 14.960 66.410 15.095 ;
        RECT 62.120 14.805 62.290 14.960 ;
        RECT 61.670 14.635 62.290 14.805 ;
        RECT 64.415 14.925 64.585 14.960 ;
        RECT 61.670 14.585 61.840 14.635 ;
        RECT 59.175 14.020 59.455 14.140 ;
        RECT 59.175 13.850 59.245 14.020 ;
        RECT 59.415 13.850 59.455 14.020 ;
        RECT 59.175 13.650 59.455 13.850 ;
        RECT 59.175 13.480 59.245 13.650 ;
        RECT 59.415 13.480 59.455 13.650 ;
        RECT 59.625 13.760 59.795 14.310 ;
        RECT 59.975 14.230 60.305 14.550 ;
        RECT 60.655 14.270 61.205 14.585 ;
        RECT 61.415 14.270 61.840 14.585 ;
        RECT 60.135 14.100 60.305 14.230 ;
        RECT 62.390 14.100 62.720 14.465 ;
        RECT 62.930 14.270 63.285 14.790 ;
        RECT 64.015 14.585 64.245 14.790 ;
        RECT 64.415 14.755 65.640 14.925 ;
        RECT 66.845 14.830 67.175 16.255 ;
        RECT 69.460 16.245 78.100 16.415 ;
        RECT 63.470 14.390 63.800 14.465 ;
        RECT 63.470 14.220 63.565 14.390 ;
        RECT 63.735 14.220 63.800 14.390 ;
        RECT 64.015 14.285 64.730 14.585 ;
        RECT 64.900 14.330 65.300 14.585 ;
        RECT 63.470 14.115 63.800 14.220 ;
        RECT 64.900 14.115 65.070 14.330 ;
        RECT 65.470 14.160 65.640 14.755 ;
        RECT 65.890 14.760 66.560 14.790 ;
        RECT 65.890 14.590 65.965 14.760 ;
        RECT 66.135 14.590 66.560 14.760 ;
        RECT 65.890 14.330 66.560 14.590 ;
        RECT 66.800 14.160 67.130 14.560 ;
        RECT 63.470 14.100 65.070 14.115 ;
        RECT 60.135 13.945 65.070 14.100 ;
        RECT 65.240 13.990 67.130 14.160 ;
        RECT 67.375 14.140 67.630 15.990 ;
        RECT 60.135 13.930 63.800 13.945 ;
        RECT 65.240 13.775 65.410 13.990 ;
        RECT 59.625 13.590 61.360 13.760 ;
        RECT 59.175 13.360 59.455 13.480 ;
        RECT 48.780 12.945 57.420 13.115 ;
        RECT 59.715 13.095 60.070 13.420 ;
        RECT 61.030 13.365 61.360 13.590 ;
        RECT 61.570 13.590 63.000 13.760 ;
        RECT 61.570 13.430 61.980 13.590 ;
        RECT 62.670 13.430 63.000 13.590 ;
        RECT 62.160 13.095 62.490 13.420 ;
        RECT 63.170 13.095 63.645 13.720 ;
        RECT 64.135 13.605 65.410 13.775 ;
        RECT 65.580 13.650 66.680 13.820 ;
        RECT 64.135 13.445 64.465 13.605 ;
        RECT 65.580 13.435 65.750 13.650 ;
        RECT 66.350 13.490 66.680 13.650 ;
        RECT 64.645 13.265 65.750 13.435 ;
        RECT 65.920 13.095 66.170 13.480 ;
        RECT 66.870 13.095 67.120 13.780 ;
        RECT 67.300 13.360 67.630 14.140 ;
        RECT 69.545 14.820 69.815 15.980 ;
        RECT 70.015 15.050 70.345 16.245 ;
        RECT 71.540 15.120 71.870 15.755 ;
        RECT 70.515 14.950 71.870 15.120 ;
        RECT 72.070 15.460 72.320 15.755 ;
        RECT 72.540 15.630 72.870 16.245 ;
        RECT 73.060 15.460 73.390 15.755 ;
        RECT 72.070 15.290 73.390 15.460 ;
        RECT 73.565 15.305 73.895 16.245 ;
        RECT 72.070 14.965 72.320 15.290 ;
        RECT 74.530 15.120 74.955 15.755 ;
        RECT 70.515 14.880 70.685 14.950 ;
        RECT 69.545 14.130 69.715 14.820 ;
        RECT 69.995 14.710 70.685 14.880 ;
        RECT 69.995 14.630 70.165 14.710 ;
        RECT 69.885 14.300 70.165 14.630 ;
        RECT 71.025 14.575 71.255 14.780 ;
        RECT 71.540 14.745 71.870 14.950 ;
        RECT 72.490 14.950 74.955 15.120 ;
        RECT 75.125 15.255 75.410 15.755 ;
        RECT 75.580 15.500 76.285 16.245 ;
        RECT 76.460 15.255 76.780 15.830 ;
        RECT 75.125 15.085 76.780 15.255 ;
        RECT 76.450 14.950 76.780 15.085 ;
        RECT 72.490 14.795 72.660 14.950 ;
        RECT 72.040 14.625 72.660 14.795 ;
        RECT 74.785 14.915 74.955 14.950 ;
        RECT 72.040 14.575 72.210 14.625 ;
        RECT 69.545 14.010 69.825 14.130 ;
        RECT 69.545 13.840 69.615 14.010 ;
        RECT 69.785 13.840 69.825 14.010 ;
        RECT 69.545 13.640 69.825 13.840 ;
        RECT 69.545 13.470 69.615 13.640 ;
        RECT 69.785 13.470 69.825 13.640 ;
        RECT 69.995 13.750 70.165 14.300 ;
        RECT 70.345 14.220 70.675 14.540 ;
        RECT 71.025 14.260 71.575 14.575 ;
        RECT 71.785 14.260 72.210 14.575 ;
        RECT 70.505 14.090 70.675 14.220 ;
        RECT 72.760 14.090 73.090 14.455 ;
        RECT 73.300 14.260 73.655 14.780 ;
        RECT 74.385 14.575 74.615 14.780 ;
        RECT 74.785 14.745 76.010 14.915 ;
        RECT 77.215 14.820 77.545 16.245 ;
        RECT 79.770 16.225 88.410 16.395 ;
        RECT 73.840 14.380 74.170 14.455 ;
        RECT 73.840 14.210 73.935 14.380 ;
        RECT 74.105 14.210 74.170 14.380 ;
        RECT 74.385 14.275 75.100 14.575 ;
        RECT 75.270 14.320 75.670 14.575 ;
        RECT 73.840 14.105 74.170 14.210 ;
        RECT 75.270 14.105 75.440 14.320 ;
        RECT 75.840 14.150 76.010 14.745 ;
        RECT 76.260 14.750 76.930 14.780 ;
        RECT 76.260 14.580 76.335 14.750 ;
        RECT 76.505 14.580 76.930 14.750 ;
        RECT 76.260 14.320 76.930 14.580 ;
        RECT 77.745 14.700 78.000 15.980 ;
        RECT 79.855 14.800 80.125 15.960 ;
        RECT 80.325 15.030 80.655 16.225 ;
        RECT 81.850 15.100 82.180 15.735 ;
        RECT 80.825 14.930 82.180 15.100 ;
        RECT 82.380 15.440 82.630 15.735 ;
        RECT 82.850 15.610 83.180 16.225 ;
        RECT 83.370 15.440 83.700 15.735 ;
        RECT 82.380 15.270 83.700 15.440 ;
        RECT 83.875 15.285 84.205 16.225 ;
        RECT 82.380 14.945 82.630 15.270 ;
        RECT 84.840 15.100 85.265 15.735 ;
        RECT 80.825 14.860 80.995 14.930 ;
        RECT 77.170 14.150 77.500 14.550 ;
        RECT 73.840 14.090 75.440 14.105 ;
        RECT 70.505 13.935 75.440 14.090 ;
        RECT 75.610 13.980 77.500 14.150 ;
        RECT 77.745 14.530 78.010 14.700 ;
        RECT 77.745 14.130 78.000 14.530 ;
        RECT 70.505 13.920 74.170 13.935 ;
        RECT 75.610 13.765 75.780 13.980 ;
        RECT 69.995 13.580 71.730 13.750 ;
        RECT 69.545 13.350 69.825 13.470 ;
        RECT 59.090 12.925 67.730 13.095 ;
        RECT 70.085 13.085 70.440 13.410 ;
        RECT 71.400 13.355 71.730 13.580 ;
        RECT 71.940 13.580 73.370 13.750 ;
        RECT 71.940 13.420 72.350 13.580 ;
        RECT 73.040 13.420 73.370 13.580 ;
        RECT 72.530 13.085 72.860 13.410 ;
        RECT 73.540 13.085 74.015 13.710 ;
        RECT 74.505 13.595 75.780 13.765 ;
        RECT 75.950 13.640 77.050 13.810 ;
        RECT 74.505 13.435 74.835 13.595 ;
        RECT 75.950 13.425 76.120 13.640 ;
        RECT 76.720 13.480 77.050 13.640 ;
        RECT 75.015 13.255 76.120 13.425 ;
        RECT 76.290 13.085 76.540 13.470 ;
        RECT 77.240 13.085 77.490 13.770 ;
        RECT 77.670 13.350 78.000 14.130 ;
        RECT 79.855 14.110 80.025 14.800 ;
        RECT 80.305 14.690 80.995 14.860 ;
        RECT 80.305 14.610 80.475 14.690 ;
        RECT 80.195 14.280 80.475 14.610 ;
        RECT 81.335 14.555 81.565 14.760 ;
        RECT 81.850 14.725 82.180 14.930 ;
        RECT 82.800 14.930 85.265 15.100 ;
        RECT 85.435 15.235 85.720 15.735 ;
        RECT 85.890 15.480 86.595 16.225 ;
        RECT 86.770 15.235 87.090 15.810 ;
        RECT 85.435 15.065 87.090 15.235 ;
        RECT 86.760 14.930 87.090 15.065 ;
        RECT 82.800 14.775 82.970 14.930 ;
        RECT 82.350 14.605 82.970 14.775 ;
        RECT 85.095 14.895 85.265 14.930 ;
        RECT 82.350 14.555 82.520 14.605 ;
        RECT 79.855 13.990 80.135 14.110 ;
        RECT 79.855 13.820 79.925 13.990 ;
        RECT 80.095 13.820 80.135 13.990 ;
        RECT 79.855 13.620 80.135 13.820 ;
        RECT 79.855 13.450 79.925 13.620 ;
        RECT 80.095 13.450 80.135 13.620 ;
        RECT 80.305 13.730 80.475 14.280 ;
        RECT 80.655 14.200 80.985 14.520 ;
        RECT 81.335 14.240 81.885 14.555 ;
        RECT 82.095 14.240 82.520 14.555 ;
        RECT 80.815 14.070 80.985 14.200 ;
        RECT 83.070 14.070 83.400 14.435 ;
        RECT 83.610 14.240 83.965 14.760 ;
        RECT 84.695 14.555 84.925 14.760 ;
        RECT 85.095 14.725 86.320 14.895 ;
        RECT 87.525 14.800 87.855 16.225 ;
        RECT 88.055 15.840 88.310 15.960 ;
        RECT 88.055 15.670 88.085 15.840 ;
        RECT 88.255 15.670 88.310 15.840 ;
        RECT 88.055 15.470 88.310 15.670 ;
        RECT 88.055 15.300 88.085 15.470 ;
        RECT 88.255 15.300 88.310 15.470 ;
        RECT 88.055 15.100 88.310 15.300 ;
        RECT 88.055 14.930 88.085 15.100 ;
        RECT 88.255 14.930 88.310 15.100 ;
        RECT 84.150 14.360 84.480 14.435 ;
        RECT 84.150 14.190 84.245 14.360 ;
        RECT 84.415 14.190 84.480 14.360 ;
        RECT 84.695 14.255 85.410 14.555 ;
        RECT 85.580 14.300 85.980 14.555 ;
        RECT 84.150 14.085 84.480 14.190 ;
        RECT 85.580 14.085 85.750 14.300 ;
        RECT 86.150 14.130 86.320 14.725 ;
        RECT 86.570 14.730 87.240 14.760 ;
        RECT 86.570 14.560 86.645 14.730 ;
        RECT 86.815 14.560 87.240 14.730 ;
        RECT 86.570 14.300 87.240 14.560 ;
        RECT 88.055 14.730 88.310 14.930 ;
        RECT 88.055 14.560 88.085 14.730 ;
        RECT 88.255 14.560 88.310 14.730 ;
        RECT 87.480 14.130 87.810 14.530 ;
        RECT 84.150 14.070 85.750 14.085 ;
        RECT 80.815 13.915 85.750 14.070 ;
        RECT 85.920 13.960 87.810 14.130 ;
        RECT 88.055 14.360 88.310 14.560 ;
        RECT 88.055 14.190 88.085 14.360 ;
        RECT 88.255 14.190 88.310 14.360 ;
        RECT 88.055 14.110 88.310 14.190 ;
        RECT 87.980 13.990 88.310 14.110 ;
        RECT 80.815 13.900 84.480 13.915 ;
        RECT 85.920 13.745 86.090 13.960 ;
        RECT 87.980 13.820 88.085 13.990 ;
        RECT 88.255 13.820 88.310 13.990 ;
        RECT 80.305 13.560 82.040 13.730 ;
        RECT 79.855 13.330 80.135 13.450 ;
        RECT 69.460 12.915 78.100 13.085 ;
        RECT 80.395 13.065 80.750 13.390 ;
        RECT 81.710 13.335 82.040 13.560 ;
        RECT 82.250 13.560 83.680 13.730 ;
        RECT 82.250 13.400 82.660 13.560 ;
        RECT 83.350 13.400 83.680 13.560 ;
        RECT 82.840 13.065 83.170 13.390 ;
        RECT 83.850 13.065 84.325 13.690 ;
        RECT 84.815 13.575 86.090 13.745 ;
        RECT 86.260 13.620 87.360 13.790 ;
        RECT 84.815 13.415 85.145 13.575 ;
        RECT 86.260 13.405 86.430 13.620 ;
        RECT 87.030 13.460 87.360 13.620 ;
        RECT 85.325 13.235 86.430 13.405 ;
        RECT 86.600 13.065 86.850 13.450 ;
        RECT 87.550 13.065 87.800 13.750 ;
        RECT 87.980 13.620 88.310 13.820 ;
        RECT 87.980 13.450 88.085 13.620 ;
        RECT 88.255 13.450 88.310 13.620 ;
        RECT 87.980 13.330 88.310 13.450 ;
        RECT 79.770 12.895 88.410 13.065 ;
      LAYER met1 ;
        RECT 138.120 224.730 138.760 225.210 ;
        RECT 138.120 47.375 138.310 224.730 ;
        RECT 82.325 47.185 138.310 47.375 ;
        RECT 7.340 36.000 15.980 36.490 ;
        RECT 6.750 34.650 9.430 34.755 ;
        RECT 11.275 34.650 11.565 34.695 ;
        RECT 12.235 34.650 12.525 34.695 ;
        RECT 6.750 34.510 12.525 34.650 ;
        RECT 6.750 34.425 9.430 34.510 ;
        RECT 11.275 34.465 11.565 34.510 ;
        RECT 12.235 34.465 12.525 34.510 ;
        RECT 6.750 29.005 7.040 34.425 ;
        RECT 11.740 33.160 12.070 34.365 ;
        RECT 14.310 34.345 14.640 36.000 ;
        RECT 17.750 35.840 26.390 36.330 ;
        RECT 28.050 35.980 36.690 36.470 ;
        RECT 38.360 36.010 47.000 36.500 ;
        RECT 15.630 34.535 19.550 34.695 ;
        RECT 15.630 34.490 19.575 34.535 ;
        RECT 21.685 34.490 21.975 34.535 ;
        RECT 22.645 34.490 22.935 34.535 ;
        RECT 15.630 34.350 22.935 34.490 ;
        RECT 15.630 34.305 19.575 34.350 ;
        RECT 21.685 34.305 21.975 34.350 ;
        RECT 22.645 34.305 22.935 34.350 ;
        RECT 15.630 34.215 19.550 34.305 ;
        RECT 24.640 34.225 24.900 35.840 ;
        RECT 25.940 34.675 29.860 34.845 ;
        RECT 25.940 34.630 29.875 34.675 ;
        RECT 31.985 34.630 32.275 34.675 ;
        RECT 32.945 34.630 33.235 34.675 ;
        RECT 25.940 34.490 33.235 34.630 ;
        RECT 25.940 34.445 29.875 34.490 ;
        RECT 31.985 34.445 32.275 34.490 ;
        RECT 32.945 34.445 33.235 34.490 ;
        RECT 25.940 34.365 29.860 34.445 ;
        RECT 7.340 32.670 15.980 33.160 ;
        RECT 22.090 33.000 22.440 34.205 ;
        RECT 32.420 33.140 32.780 34.295 ;
        RECT 34.910 34.225 35.230 35.980 ;
        RECT 36.330 34.660 40.250 34.775 ;
        RECT 42.295 34.660 42.585 34.705 ;
        RECT 43.255 34.660 43.545 34.705 ;
        RECT 45.240 34.665 45.760 36.010 ;
        RECT 36.330 34.520 43.545 34.660 ;
        RECT 36.330 34.295 40.250 34.520 ;
        RECT 42.295 34.475 42.585 34.520 ;
        RECT 43.255 34.475 43.545 34.520 ;
        RECT 42.760 33.170 43.050 34.365 ;
        RECT 45.190 34.345 45.780 34.665 ;
        RECT 46.680 34.065 47.790 34.375 ;
        RECT 17.750 32.510 26.390 33.000 ;
        RECT 28.050 32.650 36.690 33.140 ;
        RECT 38.360 32.680 47.000 33.170 ;
        RECT 45.900 30.700 46.390 32.140 ;
        RECT 47.440 31.715 47.790 34.065 ;
        RECT 7.260 30.070 15.900 30.560 ;
        RECT 17.580 30.150 26.220 30.640 ;
        RECT 7.350 29.005 7.630 29.045 ;
        RECT 6.740 28.725 7.630 29.005 ;
        RECT 8.630 27.230 9.020 28.925 ;
        RECT 11.170 28.875 11.570 30.070 ;
        RECT 10.715 28.720 11.005 28.765 ;
        RECT 11.675 28.720 11.965 28.765 ;
        RECT 14.020 28.720 17.940 28.915 ;
        RECT 10.715 28.580 17.940 28.720 ;
        RECT 10.715 28.535 11.005 28.580 ;
        RECT 11.675 28.535 11.965 28.580 ;
        RECT 14.020 28.435 17.940 28.580 ;
        RECT 18.950 27.310 19.330 28.955 ;
        RECT 21.520 28.945 21.850 30.150 ;
        RECT 27.890 29.990 36.530 30.480 ;
        RECT 21.035 28.800 21.325 28.845 ;
        RECT 21.995 28.800 22.285 28.845 ;
        RECT 24.360 28.800 28.280 28.995 ;
        RECT 21.035 28.660 28.280 28.800 ;
        RECT 21.035 28.615 21.325 28.660 ;
        RECT 21.995 28.615 22.285 28.660 ;
        RECT 24.360 28.515 28.280 28.660 ;
        RECT 7.260 26.740 15.900 27.230 ;
        RECT 17.580 26.820 26.220 27.310 ;
        RECT 29.140 27.150 29.580 28.865 ;
        RECT 31.830 28.805 32.190 29.990 ;
        RECT 38.260 29.960 46.900 30.450 ;
        RECT 31.345 28.640 31.635 28.685 ;
        RECT 32.305 28.640 32.595 28.685 ;
        RECT 34.540 28.640 38.670 28.885 ;
        RECT 31.345 28.500 38.670 28.640 ;
        RECT 31.345 28.455 31.635 28.500 ;
        RECT 32.305 28.455 32.595 28.500 ;
        RECT 34.540 28.495 38.670 28.500 ;
        RECT 34.705 28.455 34.995 28.495 ;
        RECT 27.890 26.660 36.530 27.150 ;
        RECT 39.510 27.120 39.950 28.835 ;
        RECT 42.200 28.775 42.560 29.960 ;
        RECT 47.400 28.715 47.750 31.515 ;
        RECT 49.230 30.700 49.720 32.140 ;
        RECT 41.715 28.610 42.005 28.655 ;
        RECT 42.675 28.610 42.965 28.655 ;
        RECT 44.720 28.610 47.750 28.715 ;
        RECT 82.325 28.815 82.515 47.185 ;
        RECT 84.590 30.325 88.910 30.815 ;
        RECT 88.385 29.080 152.475 29.450 ;
        RECT 85.095 28.815 85.440 29.000 ;
        RECT 88.385 28.970 152.530 29.080 ;
        RECT 88.385 28.860 152.540 28.970 ;
        RECT 82.325 28.650 85.440 28.815 ;
        RECT 82.325 28.625 85.425 28.650 ;
        RECT 41.715 28.495 47.750 28.610 ;
        RECT 41.715 28.470 47.740 28.495 ;
        RECT 41.715 28.425 42.005 28.470 ;
        RECT 42.675 28.425 42.965 28.470 ;
        RECT 44.720 28.375 47.740 28.470 ;
        RECT 86.460 28.430 86.870 28.820 ;
        RECT 87.030 28.350 87.560 28.800 ;
        RECT 149.000 28.690 152.540 28.860 ;
        RECT 38.260 26.630 46.900 27.120 ;
        RECT 84.590 26.995 88.910 27.485 ;
        RECT 4.450 22.450 4.860 22.580 ;
        RECT 40.490 22.450 41.930 22.505 ;
        RECT 4.450 22.205 41.930 22.450 ;
        RECT 4.450 21.930 4.860 22.205 ;
        RECT 40.490 22.015 41.930 22.205 ;
        RECT 40.910 20.300 41.330 20.870 ;
        RECT 41.520 20.790 41.920 21.020 ;
        RECT 41.535 20.430 41.840 20.790 ;
        RECT 41.100 20.220 41.325 20.300 ;
        RECT 1.470 19.035 2.420 19.400 ;
        RECT 40.490 19.035 41.930 19.175 ;
        RECT 1.470 18.665 42.465 19.035 ;
        RECT 1.470 18.420 2.420 18.665 ;
        RECT 7.490 16.540 16.130 16.675 ;
        RECT 17.800 16.540 26.440 16.655 ;
        RECT 7.490 16.430 16.160 16.540 ;
        RECT 16.130 16.300 16.160 16.430 ;
        RECT 17.780 16.490 26.440 16.540 ;
        RECT 28.170 16.490 36.810 16.645 ;
        RECT 38.480 16.490 47.120 16.625 ;
        RECT 48.780 16.500 57.420 16.605 ;
        RECT 17.780 16.410 26.460 16.490 ;
        RECT 17.780 16.300 17.800 16.410 ;
        RECT 26.440 16.250 26.460 16.410 ;
        RECT 28.080 16.400 36.820 16.490 ;
        RECT 28.080 16.250 28.170 16.400 ;
        RECT 36.810 16.250 36.820 16.400 ;
        RECT 38.440 16.380 47.120 16.490 ;
        RECT 48.740 16.430 57.420 16.500 ;
        RECT 59.090 16.450 67.730 16.585 ;
        RECT 69.460 16.450 78.100 16.575 ;
        RECT 79.770 16.450 88.410 16.555 ;
        RECT 59.090 16.430 67.790 16.450 ;
        RECT 38.440 16.250 38.480 16.380 ;
        RECT 48.740 16.360 57.450 16.430 ;
        RECT 48.740 16.260 48.780 16.360 ;
        RECT 57.420 16.190 57.450 16.360 ;
        RECT 59.070 16.340 67.790 16.430 ;
        RECT 59.070 16.190 59.090 16.340 ;
        RECT 67.730 16.210 67.790 16.340 ;
        RECT 69.410 16.330 78.100 16.450 ;
        RECT 69.410 16.210 69.460 16.330 ;
        RECT 79.680 16.310 88.410 16.450 ;
        RECT 79.680 16.210 79.770 16.310 ;
        RECT 7.520 16.180 8.020 16.185 ;
        RECT 9.025 14.835 9.315 14.880 ;
        RECT 10.480 14.835 10.960 15.050 ;
        RECT 11.425 14.850 11.715 14.880 ;
        RECT 11.425 14.835 11.485 14.850 ;
        RECT 9.025 14.695 11.485 14.835 ;
        RECT 9.025 14.650 9.315 14.695 ;
        RECT 10.480 14.550 10.960 14.695 ;
        RECT 11.425 14.680 11.485 14.695 ;
        RECT 11.655 14.835 11.715 14.850 ;
        RECT 12.385 14.835 12.675 14.880 ;
        RECT 14.590 14.870 14.860 16.185 ;
        RECT 11.655 14.695 12.675 14.835 ;
        RECT 11.655 14.680 11.715 14.695 ;
        RECT 11.425 14.650 11.715 14.680 ;
        RECT 12.385 14.650 12.675 14.695 ;
        RECT 11.880 14.150 12.230 14.550 ;
        RECT 14.290 14.440 14.950 14.870 ;
        RECT 15.830 14.860 19.600 14.890 ;
        RECT 15.830 14.815 19.625 14.860 ;
        RECT 21.735 14.815 22.025 14.860 ;
        RECT 22.695 14.815 22.985 14.860 ;
        RECT 24.900 14.850 25.170 16.165 ;
        RECT 26.090 14.860 26.370 15.020 ;
        RECT 26.090 14.850 29.890 14.860 ;
        RECT 15.830 14.675 22.985 14.815 ;
        RECT 15.830 14.630 19.625 14.675 ;
        RECT 21.735 14.630 22.025 14.675 ;
        RECT 22.695 14.630 22.985 14.675 ;
        RECT 15.830 14.560 19.600 14.630 ;
        RECT 11.960 13.345 12.120 14.150 ;
        RECT 22.190 14.130 22.540 14.530 ;
        RECT 24.600 14.420 25.260 14.850 ;
        RECT 26.090 14.805 29.995 14.850 ;
        RECT 32.105 14.805 32.395 14.850 ;
        RECT 33.065 14.805 33.355 14.850 ;
        RECT 35.270 14.840 35.540 16.155 ;
        RECT 26.090 14.665 33.355 14.805 ;
        RECT 26.090 14.620 29.995 14.665 ;
        RECT 32.105 14.620 32.395 14.665 ;
        RECT 33.065 14.620 33.355 14.665 ;
        RECT 26.090 14.570 29.890 14.620 ;
        RECT 26.090 14.550 26.370 14.570 ;
        RECT 22.270 13.325 22.430 14.130 ;
        RECT 32.560 14.120 32.910 14.520 ;
        RECT 34.970 14.410 35.630 14.840 ;
        RECT 36.510 14.830 40.280 14.860 ;
        RECT 36.510 14.785 40.305 14.830 ;
        RECT 42.415 14.785 42.705 14.830 ;
        RECT 43.375 14.785 43.665 14.830 ;
        RECT 45.580 14.820 45.850 16.135 ;
        RECT 36.510 14.645 43.665 14.785 ;
        RECT 36.510 14.600 40.305 14.645 ;
        RECT 42.415 14.600 42.705 14.645 ;
        RECT 43.375 14.600 43.665 14.645 ;
        RECT 36.510 14.530 40.280 14.600 ;
        RECT 7.480 13.100 7.490 13.320 ;
        RECT 32.640 13.315 32.800 14.120 ;
        RECT 42.870 14.100 43.220 14.500 ;
        RECT 45.280 14.390 45.940 14.820 ;
        RECT 46.810 14.810 50.570 14.830 ;
        RECT 46.770 14.765 50.605 14.810 ;
        RECT 52.715 14.765 53.005 14.810 ;
        RECT 53.675 14.765 53.965 14.810 ;
        RECT 55.880 14.800 56.150 16.115 ;
        RECT 46.770 14.625 53.965 14.765 ;
        RECT 46.770 14.580 50.605 14.625 ;
        RECT 52.715 14.580 53.005 14.625 ;
        RECT 53.675 14.580 53.965 14.625 ;
        RECT 46.770 14.500 50.570 14.580 ;
        RECT 46.810 14.490 50.570 14.500 ;
        RECT 42.950 13.295 43.110 14.100 ;
        RECT 53.170 14.080 53.520 14.480 ;
        RECT 55.580 14.370 56.240 14.800 ;
        RECT 57.120 14.790 60.890 14.820 ;
        RECT 57.120 14.745 60.915 14.790 ;
        RECT 63.025 14.745 63.315 14.790 ;
        RECT 63.985 14.745 64.275 14.790 ;
        RECT 66.190 14.780 66.460 16.095 ;
        RECT 67.380 14.790 67.660 14.950 ;
        RECT 67.380 14.780 71.180 14.790 ;
        RECT 57.120 14.605 64.275 14.745 ;
        RECT 57.120 14.560 60.915 14.605 ;
        RECT 63.025 14.560 63.315 14.605 ;
        RECT 63.985 14.560 64.275 14.605 ;
        RECT 57.120 14.490 60.890 14.560 ;
        RECT 53.250 13.275 53.410 14.080 ;
        RECT 63.480 14.060 63.830 14.460 ;
        RECT 65.890 14.350 66.550 14.780 ;
        RECT 67.380 14.735 71.285 14.780 ;
        RECT 73.395 14.735 73.685 14.780 ;
        RECT 74.355 14.735 74.645 14.780 ;
        RECT 76.560 14.770 76.830 16.085 ;
        RECT 67.380 14.595 74.645 14.735 ;
        RECT 67.380 14.550 71.285 14.595 ;
        RECT 73.395 14.550 73.685 14.595 ;
        RECT 74.355 14.550 74.645 14.595 ;
        RECT 67.380 14.500 71.180 14.550 ;
        RECT 67.380 14.480 67.660 14.500 ;
        RECT 63.560 13.255 63.720 14.060 ;
        RECT 73.850 14.050 74.200 14.450 ;
        RECT 76.260 14.340 76.920 14.770 ;
        RECT 77.800 14.760 81.570 14.790 ;
        RECT 77.800 14.715 81.595 14.760 ;
        RECT 83.705 14.715 83.995 14.760 ;
        RECT 84.665 14.715 84.955 14.760 ;
        RECT 86.870 14.750 87.140 16.065 ;
        RECT 77.800 14.575 84.955 14.715 ;
        RECT 77.800 14.530 81.595 14.575 ;
        RECT 83.705 14.530 83.995 14.575 ;
        RECT 84.665 14.530 84.955 14.575 ;
        RECT 77.800 14.460 81.570 14.530 ;
        RECT 73.930 13.245 74.090 14.050 ;
        RECT 84.160 14.030 84.510 14.430 ;
        RECT 86.570 14.320 87.230 14.750 ;
        RECT 88.050 14.360 88.690 14.380 ;
        RECT 84.240 13.225 84.400 14.030 ;
        RECT 88.050 13.790 89.700 14.360 ;
        RECT 16.130 13.100 16.160 13.190 ;
        RECT 7.480 12.950 16.160 13.100 ;
        RECT 17.780 13.080 17.800 13.190 ;
        RECT 26.440 13.080 26.510 13.210 ;
        RECT 17.780 12.970 26.510 13.080 ;
        RECT 28.130 13.070 28.170 13.210 ;
        RECT 28.130 12.970 36.810 13.070 ;
        RECT 17.780 12.950 26.440 12.970 ;
        RECT 7.480 12.910 16.130 12.950 ;
        RECT 7.490 12.855 16.130 12.910 ;
        RECT 17.800 12.835 26.440 12.950 ;
        RECT 28.170 12.825 36.810 12.970 ;
        RECT 38.410 13.050 38.480 13.130 ;
        RECT 47.120 13.050 47.130 13.130 ;
        RECT 38.410 12.890 47.130 13.050 ;
        RECT 48.750 13.030 48.780 13.130 ;
        RECT 57.420 13.030 57.450 13.110 ;
        RECT 48.750 12.890 57.450 13.030 ;
        RECT 38.480 12.805 47.120 12.890 ;
        RECT 48.780 12.870 57.450 12.890 ;
        RECT 59.070 13.010 59.090 13.110 ;
        RECT 67.730 13.010 67.780 13.110 ;
        RECT 59.070 12.870 67.780 13.010 ;
        RECT 69.400 13.000 69.460 13.110 ;
        RECT 78.100 13.000 78.120 13.130 ;
        RECT 69.400 12.890 78.120 13.000 ;
        RECT 79.740 12.980 79.770 13.130 ;
        RECT 79.740 12.890 88.410 12.980 ;
        RECT 69.400 12.870 78.100 12.890 ;
        RECT 48.780 12.785 57.420 12.870 ;
        RECT 59.090 12.765 67.730 12.870 ;
        RECT 69.460 12.755 78.100 12.870 ;
        RECT 79.770 12.735 88.410 12.890 ;
        RECT 151.960 0.870 152.540 28.690 ;
        RECT 151.950 0.170 152.570 0.870 ;
      LAYER met2 ;
        RECT 138.120 224.730 138.760 225.210 ;
        RECT 10.620 36.030 11.590 36.490 ;
        RECT 21.630 35.870 22.600 36.330 ;
        RECT 31.760 36.020 32.730 36.480 ;
        RECT 42.130 36.060 43.100 36.520 ;
        RECT 10.750 32.690 11.610 33.130 ;
        RECT 21.720 32.490 22.550 32.990 ;
        RECT 31.990 32.630 32.820 33.130 ;
        RECT 42.370 32.650 43.200 33.150 ;
        RECT 47.340 32.530 87.020 33.340 ;
        RECT 45.910 31.160 46.330 31.920 ;
        RECT 10.760 30.080 11.590 30.580 ;
        RECT 21.730 30.200 22.560 30.700 ;
        RECT 31.990 30.110 32.820 30.610 ;
        RECT 49.240 30.590 49.750 32.230 ;
        RECT 42.370 30.000 43.200 30.500 ;
        RECT 84.570 30.300 85.010 30.830 ;
        RECT 86.460 29.300 87.000 32.530 ;
        RECT 86.460 28.430 86.870 29.300 ;
        RECT 11.240 26.760 12.210 27.220 ;
        RECT 21.330 26.850 22.300 27.310 ;
        RECT 31.630 26.680 32.600 27.140 ;
        RECT 42.230 26.610 43.200 27.070 ;
        RECT 85.900 26.980 86.650 27.480 ;
        RECT 4.450 21.930 4.860 22.580 ;
        RECT 87.030 21.310 87.550 28.800 ;
        RECT 10.630 20.350 41.270 20.870 ;
        RECT 41.485 20.640 89.610 21.310 ;
        RECT 10.630 20.220 11.220 20.350 ;
        RECT 1.470 18.420 2.420 19.400 ;
        RECT 10.640 14.970 10.940 20.220 ;
        RECT 11.950 16.310 13.240 16.680 ;
        RECT 22.220 16.270 23.510 16.640 ;
        RECT 31.960 16.320 33.250 16.690 ;
        RECT 42.490 16.230 43.780 16.600 ;
        RECT 53.050 16.270 54.340 16.640 ;
        RECT 63.260 16.210 64.550 16.580 ;
        RECT 73.510 16.180 74.800 16.550 ;
        RECT 83.850 16.200 85.140 16.570 ;
        RECT 10.520 14.610 10.970 14.970 ;
        RECT 88.940 13.870 89.610 20.640 ;
        RECT 11.740 12.880 13.030 13.250 ;
        RECT 21.820 12.840 23.110 13.210 ;
        RECT 32.080 12.940 33.370 13.310 ;
        RECT 42.320 12.860 43.610 13.230 ;
        RECT 53.180 12.860 54.470 13.230 ;
        RECT 63.240 12.820 64.530 13.190 ;
        RECT 73.680 12.840 74.970 13.210 ;
        RECT 83.960 12.830 85.250 13.200 ;
        RECT 151.950 0.170 152.570 0.870 ;
      LAYER met3 ;
        RECT 138.120 224.730 138.760 225.210 ;
        RECT 1.950 36.700 49.825 37.710 ;
        RECT 10.615 36.075 11.625 36.700 ;
        RECT 21.615 35.895 22.625 36.700 ;
        RECT 31.725 36.045 32.735 36.700 ;
        RECT 42.145 36.045 43.155 36.700 ;
        RECT 10.750 31.980 11.630 33.190 ;
        RECT 21.710 31.980 22.590 32.950 ;
        RECT 31.970 31.980 32.850 33.130 ;
        RECT 42.350 31.980 43.230 33.170 ;
        RECT 5.100 31.100 46.450 31.980 ;
        RECT 10.750 30.080 11.630 31.100 ;
        RECT 21.710 30.180 22.590 31.100 ;
        RECT 31.970 30.060 32.850 31.100 ;
        RECT 42.350 29.990 43.230 31.100 ;
        RECT 48.705 30.625 49.715 36.700 ;
        RECT 83.985 33.040 84.995 33.085 ;
        RECT 83.895 32.030 89.960 33.040 ;
        RECT 11.215 25.770 12.225 27.245 ;
        RECT 21.325 25.770 22.335 27.295 ;
        RECT 31.625 25.770 32.635 27.125 ;
        RECT 42.235 25.770 43.245 27.185 ;
        RECT 1.890 24.760 46.960 25.770 ;
        RECT 4.450 21.930 4.860 22.580 ;
        RECT 1.470 18.420 2.420 19.400 ;
        RECT 83.985 18.040 84.995 32.030 ;
        RECT 85.895 26.690 87.745 27.695 ;
        RECT 85.895 24.840 89.960 26.690 ;
        RECT 2.320 17.250 85.050 18.040 ;
        RECT 2.620 17.140 85.050 17.250 ;
        RECT 7.520 17.030 85.050 17.140 ;
        RECT 12.005 16.045 13.015 17.030 ;
        RECT 22.245 16.215 23.255 17.030 ;
        RECT 32.085 16.215 33.095 17.030 ;
        RECT 42.545 16.215 43.555 17.030 ;
        RECT 53.225 16.115 54.235 17.030 ;
        RECT 63.435 16.215 64.445 17.030 ;
        RECT 73.655 16.055 74.665 17.030 ;
        RECT 83.985 16.115 84.995 17.030 ;
        RECT 11.760 11.330 13.060 13.460 ;
        RECT 21.780 11.330 23.080 13.460 ;
        RECT 32.090 11.330 33.390 13.460 ;
        RECT 42.330 11.330 43.630 13.300 ;
        RECT 53.140 11.330 54.440 13.240 ;
        RECT 63.230 11.330 64.530 13.210 ;
        RECT 73.660 11.330 74.960 13.210 ;
        RECT 83.900 11.330 85.200 13.180 ;
        RECT 86.115 11.330 87.605 24.840 ;
        RECT 5.030 9.840 87.790 11.330 ;
        RECT 151.950 0.170 152.570 0.870 ;
      LAYER met4 ;
        RECT 138.610 224.780 138.670 225.130 ;
  END
END tt_um_ohmy90_ringOscillator
END LIBRARY

