* SPICE3 file created from tt_um_ohmy90_adders.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
C0 Y A 0.0476f
C1 Y VPWR 0.12758f
C2 A VPWR 0.03703f
C3 VGND VPB 0.00948f
C4 Y VPB 0.01774f
C5 Y VGND 0.09984f
C6 VPB A 0.04506f
C7 VPB VPWR 0.05448f
C8 VGND A 0.04004f
C9 VGND VPWR 0.03382f
C10 VGND VNB 0.25113f
C11 Y VNB 0.0961f
C12 VPWR VNB 0.21892f
C13 A VNB 0.16664f
C14 VPB VNB 0.33898f
.ends

.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X a_1290_413#
+ a_757_363# a_1478_413# a_277_47# a_750_97# a_27_413# a_923_363# a_193_47# a_834_97#
+ a_247_21# a_668_97# a_193_413# a_27_47#
X0 a_277_47# a_247_21# a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X1 VGND S0 a_247_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08138 pd=0.96719 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X2 a_834_97# a_247_21# a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=0.10858 pd=1.36 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=4318,272
X3 VGND A3 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0.08138 pd=0.96719 as=0.10855 ps=1.36 w=0.42 l=0.15
**devattr s=4316,272 d=2268,138
X4 a_1290_413# S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.08399 ps=0.95455 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X5 a_834_97# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10858 pd=1.36 as=0.08138 ps=0.96719 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X6 a_750_97# S0 a_757_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1274 pd=1.16667 as=0.10855 ps=1.36 w=0.42 l=0.15
**devattr s=4316,272 d=2268,138
X7 a_27_47# S0 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.09322 ps=1.07 w=0.42 l=0.15
**devattr s=3409,185 d=4368,272
X8 X a_1478_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12594 ps=1.49685 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X9 VPWR A1 a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.08399 pd=0.95455 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X10 VPWR S0 a_247_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.08399 pd=0.95455 as=0.1083 ps=1.36 w=0.42 l=0.15
**devattr s=4332,272 d=4316,272
X11 X a_1478_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.19997 ps=2.27273 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X12 a_193_47# A0 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.08138 ps=0.96719 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X13 a_750_97# a_1290_413# a_1478_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1274 pd=1.16667 as=0.09209 ps=0.99 w=0.42 l=0.15
**devattr s=3683,198 d=10752,424
X14 a_1478_413# S1 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09209 pd=0.99 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=3683,198
X15 a_1290_413# S1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.08138 ps=0.96719 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X16 a_277_47# a_247_21# a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.09322 pd=1.07 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3409,185
X17 a_750_97# S0 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.10855 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X18 a_923_363# a_247_21# a_750_97# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09013 pd=0.995 as=0.1274 ps=1.16667 w=0.42 l=0.15
**devattr s=2268,138 d=3605,199
X19 a_757_363# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.36 as=0.08399 ps=0.95455 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X20 VPWR A3 a_923_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.08399 pd=0.95455 as=0.09013 ps=0.995 w=0.42 l=0.15
**devattr s=3605,199 d=2268,138
X21 a_277_47# a_1290_413# a_1478_413# VNB sky130_fd_pr__nfet_01v8 ad=0.09322 pd=1.07 as=0.15102 ps=1.285 w=0.42 l=0.15
**devattr s=6041,257 d=4368,272
X22 a_193_413# A0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.36 as=0.08399 ps=0.95455 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X23 a_193_413# S0 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.36 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=4316,272
X24 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08138 pd=0.96719 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X25 a_1478_413# S1 a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=0.15102 pd=1.285 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=6041,257
C0 VPB A0 0.08019f
C1 a_668_97# S0 0.03f
C2 a_1290_413# a_247_21# 0.00705f
C3 S0 a_27_47# 0.01792f
C4 a_750_97# VPWR 0.22609f
C5 S1 a_247_21# 0
C6 a_1290_413# a_277_47# 0.33858f
C7 a_193_413# a_750_97# 0
C8 VGND VPWR 0.05896f
C9 S1 a_277_47# 0.06116f
C10 a_193_413# VGND 0
C11 A0 S0 0.00186f
C12 a_27_413# VPWR 0.08385f
C13 VPB A3 0.07252f
C14 a_27_413# a_193_413# 0.05551f
C15 a_757_363# A3 0.03224f
C16 X a_1290_413# 0.00208f
C17 a_668_97# a_750_97# 0.04662f
C18 A3 a_834_97# 0.03609f
C19 a_668_97# VGND 0.22352f
C20 X S1 0
C21 a_27_47# VGND 0.22952f
C22 a_193_413# VPWR 0.18442f
C23 S0 A3 0.00317f
C24 a_1478_413# a_247_21# 0
C25 VPB a_1290_413# 0.14223f
C26 a_193_47# VGND 0.00175f
C27 VPB S1 0.21534f
C28 a_1478_413# a_277_47# 0.09435f
C29 A2 A3 0.15492f
C30 A0 a_750_97# 0
C31 a_757_363# a_1290_413# 0.0098f
C32 a_27_413# a_27_47# 0.00987f
C33 a_1290_413# a_834_97# 0.01242f
C34 A0 VGND 0.01709f
C35 a_757_363# S1 0.00151f
C36 S1 a_834_97# 0.00189f
C37 a_668_97# VPWR 0.00181f
C38 a_247_21# a_277_47# 0.35203f
C39 a_27_47# VPWR 0.0018f
C40 A0 a_27_413# 0.04892f
C41 A2 a_1290_413# 0.00165f
C42 a_923_363# a_757_363# 0.00988f
C43 a_923_363# a_834_97# 0
C44 A2 S1 0.06853f
C45 a_1478_413# X 0.12698f
C46 a_193_47# VPWR 0
C47 a_750_97# A3 0.03406f
C48 A1 a_247_21# 0
C49 A3 VGND 0.01161f
C50 A1 a_277_47# 0.00101f
C51 A0 VPWR 0.01747f
C52 A0 a_193_413# 0.00145f
C53 VPB a_1478_413# 0.07712f
C54 X a_247_21# 0
C55 a_1290_413# a_750_97# 0.17579f
C56 X a_277_47# 0
C57 a_1290_413# VGND 0.06373f
C58 S1 a_750_97# 0.06323f
C59 S1 VGND 0.04087f
C60 VPB a_247_21# 0.22297f
C61 a_193_47# a_27_47# 0.00648f
C62 A3 VPWR 0.012f
C63 VPB a_277_47# 0.03677f
C64 a_757_363# a_247_21# 0.02645f
C65 A0 a_27_47# 0.04574f
C66 a_834_97# a_247_21# 0.02707f
C67 a_923_363# a_750_97# 0.00222f
C68 a_757_363# a_277_47# 0
C69 a_834_97# a_277_47# 0.04391f
C70 VPB A1 0.0741f
C71 A0 a_193_47# 0
C72 S0 a_247_21# 0.39319f
C73 a_1290_413# VPWR 0.0823f
C74 S0 a_277_47# 0.03381f
C75 A2 a_247_21# 0.00145f
C76 S1 VPWR 0.0409f
C77 A2 a_277_47# 0.01375f
C78 VPB X 0.01181f
C79 a_668_97# A3 0.0033f
C80 a_1478_413# a_750_97# 0.1456f
C81 a_27_47# A3 0
C82 a_1478_413# VGND 0.18885f
C83 a_923_363# VPWR 0.00225f
C84 VPB a_757_363# 0.0237f
C85 a_668_97# a_1290_413# 0
C86 VPB a_834_97# 0.00426f
C87 a_750_97# a_247_21# 0.12371f
C88 VGND a_247_21# 0.09412f
C89 a_750_97# a_277_47# 0.26678f
C90 VGND a_277_47# 0.41112f
C91 a_757_363# a_834_97# 0.01352f
C92 VPB S0 0.31074f
C93 A1 a_750_97# 0
C94 a_1478_413# VPWR 0.21151f
C95 VPB A2 0.07872f
C96 A1 VGND 0.01705f
C97 a_27_413# a_247_21# 0.00549f
C98 S0 a_757_363# 0.03305f
C99 S0 a_834_97# 0
C100 a_27_413# a_277_47# 0.05408f
C101 A2 a_757_363# 0.03541f
C102 A2 a_834_97# 0.04394f
C103 X a_750_97# 0
C104 A1 a_27_413# 0.0413f
C105 a_247_21# VPWR 0.15063f
C106 X VGND 0.05939f
C107 a_193_413# a_247_21# 0.09132f
C108 VPWR a_277_47# 0.05706f
C109 a_193_413# a_277_47# 0.0594f
C110 a_1290_413# A3 0
C111 VPB a_750_97# 0.05933f
C112 VPB VGND 0.01387f
C113 S1 A3 0
C114 A1 VPWR 0.01712f
C115 A1 a_193_413# 0
C116 a_757_363# a_750_97# 0.13413f
C117 a_750_97# a_834_97# 0.0296f
C118 VGND a_834_97# 0.09477f
C119 VPB a_27_413# 0.02285f
C120 a_668_97# a_247_21# 0.01881f
C121 a_923_363# A3 0
C122 a_27_47# a_247_21# 0.0457f
C123 S0 a_750_97# 0.09449f
C124 X VPWR 0.05937f
C125 a_668_97# a_277_47# 0.02235f
C126 S0 VGND 0.06675f
C127 S1 a_1290_413# 0.15612f
C128 a_27_47# a_277_47# 0.08551f
C129 A2 a_750_97# 0.01619f
C130 A2 VGND 0.0122f
C131 a_193_47# a_277_47# 0
C132 VPB VPWR 0.22689f
C133 A1 a_27_47# 0.03909f
C134 VPB a_193_413# 0.01733f
C135 A0 a_247_21# 0.07359f
C136 S0 a_27_413# 0
C137 a_923_363# a_1290_413# 0
C138 A0 a_277_47# 0.05427f
C139 a_757_363# VPWR 0.24812f
C140 a_834_97# VPWR 0
C141 A0 A1 0.14123f
C142 S0 VPWR 0.0687f
C143 a_750_97# VGND 0.05676f
C144 S0 a_193_413# 0.01772f
C145 A2 VPWR 0.0129f
C146 A3 a_247_21# 0.07395f
C147 VPB a_668_97# 0.00146f
C148 VPB a_27_47# 0.00324f
C149 a_1478_413# a_1290_413# 0.10432f
C150 A3 a_277_47# 0.0121f
C151 a_1478_413# S1 0.00517f
C152 a_27_413# a_750_97# 0
C153 a_668_97# a_834_97# 0.05583f
C154 a_27_413# VGND 0.00189f
C155 VGND VNB 1.07507f
C156 X VNB 0.09236f
C157 S1 VNB 0.32062f
C158 A2 VNB 0.11249f
C159 A3 VNB 0.11926f
C160 S0 VNB 0.46486f
C161 VPWR VNB 0.86887f
C162 A0 VNB 0.10257f
C163 A1 VNB 0.17585f
C164 VPB VNB 1.9337f
C165 a_834_97# VNB 0.02499f
C166 a_668_97# VNB 0.02039f
C167 a_27_47# VNB 0.04207f
C168 a_1478_413# VNB 0.16413f
C169 a_1290_413# VNB 0.2199f
C170 a_750_97# VNB 0.04192f
C171 a_757_363# VNB 0.00666f
C172 a_277_47# VNB 0.07984f
C173 a_247_21# VNB 0.34344f
C174 a_193_413# VNB 0.00373f
C175 a_27_413# VNB 0.02865f
.ends

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X a_117_297# a_285_297# a_285_47#
+ a_35_297#
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13813 ps=1.4 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.13813 pd=1.4 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.13813 pd=1.4 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13813 ps=1.4 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
C0 A a_285_297# 0.00749f
C1 B a_35_297# 0.203f
C2 VPWR B 0.07031f
C3 VPB a_285_297# 0.01327f
C4 VGND X 0.1729f
C5 VGND A 0.03254f
C6 VPWR a_35_297# 0.09604f
C7 VGND VPB 0.00696f
C8 A X 0.00166f
C9 a_285_297# B 0.05532f
C10 VGND a_117_297# 0.00177f
C11 VGND a_285_47# 0.00552f
C12 VPB X 0.01541f
C13 A VPB 0.05101f
C14 a_285_297# a_35_297# 0.02504f
C15 VPWR a_285_297# 0.24631f
C16 VGND B 0.03045f
C17 a_117_297# X 0
C18 a_285_47# X 0.00206f
C19 VGND a_35_297# 0.17666f
C20 VGND VPWR 0.06426f
C21 B X 0.01488f
C22 A B 0.22134f
C23 X a_35_297# 0.166f
C24 VPB B 0.06969f
C25 VPWR X 0.05365f
C26 A a_35_297# 0.06334f
C27 A VPWR 0.03484f
C28 VGND a_285_297# 0.00394f
C29 VPB a_35_297# 0.06993f
C30 VPB VPWR 0.06891f
C31 a_117_297# B 0.00777f
C32 a_285_47# B 0
C33 a_117_297# a_35_297# 0.00641f
C34 a_117_297# VPWR 0.00852f
C35 a_285_47# a_35_297# 0.00723f
C36 a_285_47# VPWR 0
C37 a_285_297# X 0.07125f
C38 VGND VNB 0.43488f
C39 X VNB 0.06491f
C40 VPWR VNB 0.33278f
C41 A VNB 0.16672f
C42 B VNB 0.21337f
C43 VPB VNB 0.69336f
C44 a_285_297# VNB 0.00137f
C45 a_35_297# VNB 0.25457f
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X a_145_75# a_59_75#
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.10288 pd=0.95413 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.24495 ps=2.27174 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.08777 pd=0.81645 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.10288 ps=0.95413 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.13583 ps=1.26355 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
C0 VPWR a_145_75# 0
C1 a_59_75# VPB 0.05631f
C2 VGND B 0.01146f
C3 X a_59_75# 0.10872f
C4 B VPB 0.06287f
C5 X B 0.00276f
C6 VGND VPWR 0.04608f
C7 B a_59_75# 0.14331f
C8 VPWR VPB 0.07293f
C9 A VGND 0.01472f
C10 X VPWR 0.11122f
C11 VGND a_145_75# 0.00468f
C12 VPWR a_59_75# 0.15028f
C13 A VPB 0.08057f
C14 A X 0
C15 VPWR B 0.01175f
C16 A a_59_75# 0.08088f
C17 X a_145_75# 0
C18 a_59_75# a_145_75# 0.00658f
C19 A B 0.09709f
C20 VGND VPB 0.008f
C21 VGND X 0.09933f
C22 VGND a_59_75# 0.11564f
C23 A VPWR 0.03623f
C24 X VPB 0.01265f
C25 VGND VNB 0.3114f
C26 X VNB 0.10018f
C27 B VNB 0.11287f
C28 A VNB 0.17379f
C29 VPWR VNB 0.27345f
C30 VPB VNB 0.51617f
C31 a_59_75# VNB 0.17706f
.ends

.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X a_150_297# a_68_297#
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0873 pd=0.93866 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4010,197
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0873 ps=0.93866 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1351 ps=1.45268 w=0.65 l=0.15
**devattr s=4010,197 d=6760,364
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.08622 pd=0.78972 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5830,267
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.20528 ps=1.88028 w=1 l=0.15
**devattr s=5830,267 d=13600,536
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
C0 VPB VGND 0.0112f
C1 B X 0
C2 VPWR a_150_297# 0.00193f
C3 A VPB 0.03097f
C4 VPWR VPB 0.08053f
C5 a_68_297# a_150_297# 0.00477f
C6 a_68_297# VPB 0.06114f
C7 A VGND 0.03465f
C8 VPWR VGND 0.04645f
C9 VPB B 0.0462f
C10 A VPWR 0.00846f
C11 a_150_297# X 0
C12 a_68_297# VGND 0.11796f
C13 VPB X 0.0209f
C14 A a_68_297# 0.15786f
C15 VPWR a_68_297# 0.08898f
C16 B VGND 0.04365f
C17 A B 0.07509f
C18 VGND X 0.11395f
C19 VPWR B 0.00855f
C20 A X 0.01305f
C21 VPWR X 0.12857f
C22 a_68_297# B 0.09843f
C23 a_68_297# X 0.10534f
C24 a_150_297# VGND 0
C25 VGND VNB 0.32043f
C26 X VNB 0.10095f
C27 A VNB 0.11072f
C28 B VNB 0.18272f
C29 VPWR VNB 0.26856f
C30 VPB VNB 0.51617f
C31 a_68_297# VNB 0.15387f
.ends

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X a_109_47# a_197_47# a_303_47#
+ a_27_47#
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1394 ps=0.98731 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3319 ps=2.35075 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.1394 ps=0.98731 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1394 pd=0.98731 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.15409 pd=1.04411 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1394 pd=0.98731 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.23846 ps=1.61589 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
C0 a_303_47# a_27_47# 0.00119f
C1 VPWR a_27_47# 0.32628f
C2 B a_197_47# 0.00623f
C3 B VGND 0.04527f
C4 D VPB 0.07823f
C5 a_109_47# a_27_47# 0.00578f
C6 A B 0.08391f
C7 X VPWR 0.09451f
C8 VPB VGND 0.00852f
C9 D C 0.18016f
C10 A VPB 0.09066f
C11 D a_303_47# 0.00119f
C12 D VPWR 0.02073f
C13 a_197_47# C 0.00123f
C14 VPB B 0.06433f
C15 C VGND 0.04082f
C16 X a_27_47# 0.07537f
C17 a_303_47# VGND 0.00381f
C18 VPWR a_197_47# 0
C19 VPWR VGND 0.06618f
C20 B C 0.16061f
C21 VPWR A 0.044f
C22 a_109_47# VGND 0.00223f
C23 D a_27_47# 0.10658f
C24 VPWR B 0.02308f
C25 VPB C 0.06088f
C26 a_109_47# B 0.00153f
C27 a_197_47# a_27_47# 0.00167f
C28 VGND a_27_47# 0.13176f
C29 D X 0.00746f
C30 VPWR VPB 0.07695f
C31 A a_27_47# 0.15343f
C32 X VGND 0.09025f
C33 B a_27_47# 0.12972f
C34 a_303_47# C 0.00527f
C35 VPWR C 0.02103f
C36 a_109_47# C 0
C37 VPWR a_303_47# 0
C38 VPB a_27_47# 0.08205f
C39 D VGND 0.0898f
C40 a_109_47# VPWR 0
C41 a_197_47# VGND 0.00387f
C42 X VPB 0.01107f
C43 C a_27_47# 0.05159f
C44 A VGND 0.01512f
C45 VGND VNB 0.39291f
C46 X VNB 0.09332f
C47 VPWR VNB 0.33454f
C48 D VNB 0.13027f
C49 C VNB 0.10983f
C50 B VNB 0.11212f
C51 A VNB 0.22098f
C52 VPB VNB 0.69336f
C53 a_27_47# VNB 0.17489f
.ends

.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X a_277_297# a_205_297# a_27_297#
+ a_109_297#
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.07685 ps=0.85082 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.07685 ps=0.85082 w=0.42 l=0.15
**devattr s=4368,272 d=2772,150
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0877 pd=0.79268 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=5930,268
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.11894 ps=1.31674 w=0.65 l=0.15
**devattr s=4075,198 d=7020,368
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.2088 ps=1.88732 w=1 l=0.15
**devattr s=5930,268 d=10800,508
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.07685 pd=0.85082 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2772,150 d=2268,138
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2772,150
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.07685 pd=0.85082 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2268,138 d=4075,198
C0 VPB a_27_297# 0.05168f
C1 C VPWR 0.00723f
C2 B VGND 0.01587f
C3 a_277_297# a_27_297# 0.00876f
C4 a_109_297# VGND 0
C5 VPB A 0.03298f
C6 a_277_297# A 0
C7 D VPB 0.04052f
C8 VGND C 0.0191f
C9 B a_27_297# 0.15929f
C10 a_109_297# a_27_297# 0.00695f
C11 X VPB 0.01089f
C12 B A 0.06391f
C13 X a_277_297# 0
C14 VGND VPWR 0.05464f
C15 C a_27_297# 0.15835f
C16 D B 0.00287f
C17 A C 0.02804f
C18 a_205_297# C 0.00261f
C19 X B 0
C20 a_27_297# VPWR 0.08397f
C21 D C 0.09543f
C22 A VPWR 0.00769f
C23 a_205_297# VPWR 0
C24 VPB B 0.10612f
C25 VGND a_27_297# 0.23515f
C26 D VPWR 0.00503f
C27 a_277_297# B 0
C28 A VGND 0.01596f
C29 a_205_297# VGND 0
C30 VPB C 0.03382f
C31 X VPWR 0.08784f
C32 D VGND 0.05172f
C33 a_277_297# C 0
C34 A a_27_297# 0.16258f
C35 VPB VPWR 0.07497f
C36 a_205_297# a_27_297# 0.00412f
C37 X VGND 0.03541f
C38 D a_27_297# 0.05404f
C39 a_277_297# VPWR 0
C40 B C 0.09165f
C41 a_109_297# C 0.00356f
C42 D A 0
C43 VPB VGND 0.00796f
C44 X a_27_297# 0.0991f
C45 B VPWR 0.19276f
C46 a_277_297# VGND 0
C47 a_109_297# VPWR 0
C48 X A 0.00133f
C49 VGND VNB 0.36697f
C50 X VNB 0.08835f
C51 A VNB 0.10929f
C52 C VNB 0.10488f
C53 D VNB 0.17526f
C54 B VNB 0.11467f
C55 VPWR VNB 0.28998f
C56 VPB VNB 0.60476f
C57 a_27_297# VNB 0.16291f
.ends

.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X a_181_47# a_109_47# a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07394 pd=0.75265 as=0.0805 ps=0.94333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07394 pd=0.75265 as=0.0805 ps=0.94333 w=0.42 l=0.15
**devattr s=2646,147 d=5689,267
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=1764,126
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10335 pd=0.89495 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5266,228
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0805 pd=0.94333 as=0.07394 ps=0.75265 w=0.42 l=0.15
**devattr s=2268,138 d=2646,147
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.17604 ps=1.79204 w=1 l=0.15
**devattr s=5689,267 d=10400,504
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.15995 ps=1.38505 w=0.65 l=0.15
**devattr s=5266,228 d=6760,364
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
C0 VPWR a_109_47# 0
C1 C VPB 0.0347f
C2 a_27_47# A 0.15687f
C3 B VPWR 0.12845f
C4 VGND a_181_47# 0.00261f
C5 VGND X 0.07078f
C6 a_27_47# VGND 0.13361f
C7 B VPB 0.08363f
C8 C a_181_47# 0.00151f
C9 C X 0.01492f
C10 VPB VPWR 0.07946f
C11 a_27_47# C 0.1862f
C12 VGND A 0.01538f
C13 a_27_47# a_109_47# 0.00517f
C14 X B 0.00111f
C15 a_181_47# VPWR 0
C16 a_27_47# B 0.06246f
C17 X VPWR 0.07662f
C18 a_27_47# VPWR 0.14545f
C19 a_109_47# A 0
C20 C VGND 0.07031f
C21 X VPB 0.01208f
C22 B A 0.08692f
C23 a_27_47# VPB 0.05008f
C24 VGND a_109_47# 0.00123f
C25 VPWR A 0.01846f
C26 VGND B 0.00714f
C27 VGND VPWR 0.04751f
C28 VPB A 0.0426f
C29 a_27_47# a_181_47# 0.00401f
C30 C B 0.07462f
C31 a_27_47# X 0.08704f
C32 VGND VPB 0.00604f
C33 C VPWR 0.00464f
C34 VGND VNB 0.30013f
C35 X VNB 0.09228f
C36 C VNB 0.12026f
C37 A VNB 0.17412f
C38 VPWR VNB 0.27425f
C39 B VNB 0.10179f
C40 VPB VNB 0.51617f
C41 a_27_47# VNB 0.17719f
.ends

.subckt CLA sky130_fd_sc_hd__and4_1_1/a_303_47# sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__xor2_1_0/VPB
+ sky130_fd_sc_hd__and2_1_5/VPB a_187_n2185# sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__or2_1_0/a_150_297#
+ sky130_fd_sc_hd__or4_1_0/D sky130_fd_sc_hd__and2_1_5/a_59_75# sky130_fd_sc_hd__and4_1_1/VGND
+ sky130_fd_sc_hd__and3_1_0/a_109_47# sky130_fd_sc_hd__or4_1_0/VPWR sky130_fd_sc_hd__and3_1_0/a_181_47#
+ sky130_fd_sc_hd__xor2_1_0/a_285_297# sky130_fd_sc_hd__and2_1_0/B sky130_fd_sc_hd__or4_1_0/B
+ sky130_fd_sc_hd__or4_1_0/a_109_297# sky130_fd_sc_hd__and2_1_4/VPWR sky130_fd_sc_hd__and2_1_0/A
+ VNB sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__and3_1_0/a_27_47# a_187_n2435#
+ sky130_fd_sc_hd__and3_1_0/VPWR sky130_fd_sc_hd__and4_1_1/VPB sky130_fd_sc_hd__xor2_1_0/a_285_47#
+ a_19_n2185# sky130_fd_sc_hd__xor2_1_0/a_35_297# sky130_fd_sc_hd__and2_1_4/a_145_75#
+ sky130_fd_sc_hd__and2_1_0/a_145_75# sky130_fd_sc_hd__and4_1_1/a_27_47# a_155_n4715#
+ sky130_fd_sc_hd__or4_1_0/VGND sky130_fd_sc_hd__or4_1_0/A sky130_fd_sc_hd__and2_1_4/VGND
+ sky130_fd_sc_hd__or2_1_0/a_68_297# sky130_fd_sc_hd__and2_1_0/VPB a_195_n517# a_n63_n2185#
+ a_197_n3749# sky130_fd_sc_hd__or4_1_0/X sky130_fd_sc_hd__and4_1_0/a_109_47# a_195_n767#
+ a_197_n3999# sky130_fd_sc_hd__and2_1_5/VPWR sky130_fd_sc_hd__and3_1_0/VGND sky130_fd_sc_hd__or2_1_0/VPWR
+ a_67_n1483# sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and2_1_5/a_145_75# sky130_fd_sc_hd__and2_1_0/a_59_75#
+ sky130_fd_sc_hd__and4_1_0/VPWR a_153_n1483# a_27_n517# a_69_n4715# sky130_fd_sc_hd__or2_1_0/B
+ sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__or4_1_0/a_277_297# sky130_fd_sc_hd__and4_1_0/a_197_47#
+ sky130_fd_sc_hd__and2_1_4/VPB sky130_fd_sc_hd__xor2_1_0/a_117_297# sky130_fd_sc_hd__and3_1_0/VPB
+ sky130_fd_sc_hd__and4_1_0/a_303_47# sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and4_1_1/a_109_47#
+ sky130_fd_sc_hd__or4_1_0/VPB sky130_fd_sc_hd__or4_1_0/a_27_297# a_29_n3749# sky130_fd_sc_hd__and2_1_5/VGND
+ sky130_fd_sc_hd__or4_1_0/a_205_297# sky130_fd_sc_hd__and2_1_4/a_59_75# sky130_fd_sc_hd__or2_1_0/VGND
+ a_n53_n3749# a_n55_n517# sky130_fd_sc_hd__and4_1_1/A sky130_fd_sc_hd__xor2_1_0/B
+ sky130_fd_sc_hd__and4_1_0/VGND sky130_fd_sc_hd__xor2_1_0/A sky130_fd_sc_hd__or4_1_0/C
+ sky130_fd_sc_hd__and4_1_1/VPWR a_59_n3151# sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and4_1_1/a_197_47#
+ B VPB X a_145_n3151# A
Xsky130_fd_sc_hd__xor2_1_3 A B A VNB VPB B X a_19_n2185# a_187_n2185# a_187_n2435#
+ a_n63_n2185# sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__and2_1_0 sky130_fd_sc_hd__and2_1_0/A sky130_fd_sc_hd__and2_1_0/B
+ sky130_fd_sc_hd__and2_1_0/A VNB sky130_fd_sc_hd__and2_1_0/VPB sky130_fd_sc_hd__and2_1_0/B
+ sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and2_1_0/a_145_75# sky130_fd_sc_hd__and2_1_0/a_59_75#
+ sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_1 A B A VNB VPB B X a_153_n1483# a_67_n1483# sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_3 A B A VNB VPB B X a_145_n3151# a_59_n3151# sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_2 A B A VNB VPB B X a_155_n4715# a_69_n4715# sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_4 X X sky130_fd_sc_hd__and2_1_4/VGND VNB sky130_fd_sc_hd__and2_1_4/VPB
+ sky130_fd_sc_hd__and2_1_4/VPWR sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__and2_1_4/a_145_75#
+ sky130_fd_sc_hd__and2_1_4/a_59_75# sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_5 X X sky130_fd_sc_hd__and2_1_5/VGND VNB sky130_fd_sc_hd__and2_1_5/VPB
+ sky130_fd_sc_hd__and2_1_5/VPWR sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and2_1_5/a_145_75#
+ sky130_fd_sc_hd__and2_1_5/a_59_75# sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__or2_1_0 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__or2_1_0/VGND
+ VNB sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__or2_1_0/VPWR sky130_fd_sc_hd__or4_1_0/A
+ sky130_fd_sc_hd__or2_1_0/a_150_297# sky130_fd_sc_hd__or2_1_0/a_68_297# sky130_fd_sc_hd__or2_1
Xsky130_fd_sc_hd__and4_1_0 X sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__xor2_1_0/X
+ X sky130_fd_sc_hd__and4_1_0/VGND VNB sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__and4_1_0/VPWR
+ sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__and4_1_0/a_109_47# sky130_fd_sc_hd__and4_1_0/a_197_47#
+ sky130_fd_sc_hd__and4_1_0/a_303_47# sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__and4_1
Xsky130_fd_sc_hd__and4_1_1 sky130_fd_sc_hd__and4_1_1/A X sky130_fd_sc_hd__and4_1_1/C
+ sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and4_1_1/VGND VNB sky130_fd_sc_hd__and4_1_1/VPB
+ sky130_fd_sc_hd__and4_1_1/VPWR sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__and4_1_1/a_109_47#
+ sky130_fd_sc_hd__and4_1_1/a_197_47# sky130_fd_sc_hd__and4_1_1/a_303_47# sky130_fd_sc_hd__and4_1_1/a_27_47#
+ sky130_fd_sc_hd__and4_1
Xsky130_fd_sc_hd__or4_1_0 sky130_fd_sc_hd__or4_1_0/A sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__or4_1_0/C
+ sky130_fd_sc_hd__or4_1_0/D sky130_fd_sc_hd__or4_1_0/VGND VNB sky130_fd_sc_hd__or4_1_0/VPB
+ sky130_fd_sc_hd__or4_1_0/VPWR sky130_fd_sc_hd__or4_1_0/X sky130_fd_sc_hd__or4_1_0/a_277_297#
+ sky130_fd_sc_hd__or4_1_0/a_205_297# sky130_fd_sc_hd__or4_1_0/a_27_297# sky130_fd_sc_hd__or4_1_0/a_109_297#
+ sky130_fd_sc_hd__or4_1
Xsky130_fd_sc_hd__and3_1_0 X X X sky130_fd_sc_hd__and3_1_0/VGND VNB sky130_fd_sc_hd__and3_1_0/VPB
+ sky130_fd_sc_hd__and3_1_0/VPWR sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__and3_1_0/a_181_47#
+ sky130_fd_sc_hd__and3_1_0/a_109_47# sky130_fd_sc_hd__and3_1_0/a_27_47# sky130_fd_sc_hd__and3_1
Xsky130_fd_sc_hd__xor2_1_0 sky130_fd_sc_hd__xor2_1_0/A sky130_fd_sc_hd__xor2_1_0/B
+ sky130_fd_sc_hd__xor2_1_0/A VNB sky130_fd_sc_hd__xor2_1_0/VPB sky130_fd_sc_hd__xor2_1_0/B
+ sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__xor2_1_0/a_117_297# sky130_fd_sc_hd__xor2_1_0/a_285_297#
+ sky130_fd_sc_hd__xor2_1_0/a_285_47# sky130_fd_sc_hd__xor2_1_0/a_35_297# sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_1 A B A VNB VPB B X a_27_n517# a_195_n517# a_195_n767# a_n55_n517#
+ sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_2 A B A VNB VPB B X a_29_n3749# a_197_n3749# a_197_n3999#
+ a_n53_n3749# sky130_fd_sc_hd__xor2_1
C0 a_n53_n3749# B 0.04711f
C1 sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__or4_1_0/B 0
C2 a_19_n2185# A -0
C3 sky130_fd_sc_hd__and4_1_0/VGND sky130_fd_sc_hd__and4_1_0/VPWR -0.03588f
C4 sky130_fd_sc_hd__and4_1_0/B A 0.00988f
C5 a_59_n3151# X 0.0142f
C6 sky130_fd_sc_hd__and2_1_0/B a_n55_n517# 0
C7 sky130_fd_sc_hd__or4_1_0/a_27_297# sky130_fd_sc_hd__xor2_1_0/X 0
C8 X sky130_fd_sc_hd__and4_1_1/VPB 0.00801f
C9 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__or4_1_0/A 0.34666f
C10 a_n63_n2185# a_n53_n3749# 0.00102f
C11 sky130_fd_sc_hd__and3_1_0/VPB sky130_fd_sc_hd__and3_1_0/a_27_47# -0
C12 sky130_fd_sc_hd__and3_1_0/a_109_47# A 0
C13 sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__or4_1_0/C 0
C14 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__and4_1_0/B 0
C15 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__or4_1_0/B 0
C16 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and4_1_1/VPWR 0.26064f
C17 sky130_fd_sc_hd__and2_1_5/VPWR sky130_fd_sc_hd__and4_1_1/a_303_47# 0
C18 a_27_n517# A -0
C19 sky130_fd_sc_hd__and3_1_0/a_27_47# sky130_fd_sc_hd__and4_1_0/VGND 0
C20 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__and4_1_0/VPWR 0.00502f
C21 sky130_fd_sc_hd__and4_1_1/VGND sky130_fd_sc_hd__and4_1_1/a_303_47# -0
C22 A a_197_n3749# 0
C23 sky130_fd_sc_hd__and4_1_0/a_27_47# B 0
C24 X sky130_fd_sc_hd__or4_1_0/C 0.07492f
C25 sky130_fd_sc_hd__or2_1_0/a_150_297# X 0
C26 B sky130_fd_sc_hd__and4_1_0/VPWR 0.00173f
C27 sky130_fd_sc_hd__and2_1_4/VPB sky130_fd_sc_hd__and4_1_0/VGND 0
C28 sky130_fd_sc_hd__and3_1_0/VGND sky130_fd_sc_hd__and3_1_0/a_109_47# -0
C29 sky130_fd_sc_hd__and3_1_0/VGND sky130_fd_sc_hd__and2_1_4/VPWR 0.07231f
C30 a_67_n1483# a_n55_n517# 0.00144f
C31 sky130_fd_sc_hd__or4_1_0/a_109_297# sky130_fd_sc_hd__or4_1_0/VGND -0
C32 a_195_n767# a_n55_n517# 0
C33 sky130_fd_sc_hd__and4_1_1/a_197_47# sky130_fd_sc_hd__or4_1_0/B 0
C34 sky130_fd_sc_hd__and2_1_4/a_145_75# X 0.00133f
C35 sky130_fd_sc_hd__and2_1_5/a_59_75# VPB 0
C36 VPB sky130_fd_sc_hd__and4_1_0/B 0.01097f
C37 sky130_fd_sc_hd__and2_1_0/a_59_75# sky130_fd_sc_hd__xor2_1_0/X 0
C38 sky130_fd_sc_hd__and2_1_5/VGND a_n55_n517# 0
C39 a_153_n1483# X 0.0017f
C40 sky130_fd_sc_hd__and3_1_0/a_27_47# B 0
C41 a_59_n3151# sky130_fd_sc_hd__or4_1_0/C 0
C42 sky130_fd_sc_hd__and2_1_5/VPB X 0.03446f
C43 VPB sky130_fd_sc_hd__and2_1_4/VPWR 0
C44 sky130_fd_sc_hd__and2_1_0/A sky130_fd_sc_hd__xor2_1_0/VPB 0
C45 sky130_fd_sc_hd__or4_1_0/VPB sky130_fd_sc_hd__or4_1_0/VGND -0.00395f
C46 sky130_fd_sc_hd__xor2_1_0/a_285_297# sky130_fd_sc_hd__xor2_1_0/a_35_297# 0
C47 a_69_n4715# A 0.02702f
C48 a_n63_n2185# sky130_fd_sc_hd__and3_1_0/a_27_47# 0
C49 sky130_fd_sc_hd__xor2_1_0/A sky130_fd_sc_hd__xor2_1_0/VPB -0
C50 sky130_fd_sc_hd__or2_1_0/VGND X 0.00322f
C51 sky130_fd_sc_hd__and4_1_1/A X 0.09388f
C52 B a_29_n3749# 0.00416f
C53 sky130_fd_sc_hd__and2_1_4/VGND sky130_fd_sc_hd__and2_1_4/a_59_75# -0
C54 sky130_fd_sc_hd__and3_1_0/VPB sky130_fd_sc_hd__and2_1_5/a_59_75# 0
C55 sky130_fd_sc_hd__and3_1_0/VPB sky130_fd_sc_hd__and4_1_0/B 0.00114f
C56 sky130_fd_sc_hd__xor2_1_0/X A 0
C57 sky130_fd_sc_hd__and2_1_4/VPB B 0
C58 sky130_fd_sc_hd__or4_1_0/a_27_297# sky130_fd_sc_hd__or2_1_0/A 0.00184f
C59 sky130_fd_sc_hd__and3_1_0/a_181_47# A 0
C60 sky130_fd_sc_hd__and3_1_0/VPB sky130_fd_sc_hd__and2_1_4/VPWR 0
C61 sky130_fd_sc_hd__or4_1_0/a_27_297# sky130_fd_sc_hd__or2_1_0/VPWR 0
C62 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and4_1_0/VPB 0
C63 sky130_fd_sc_hd__and2_1_5/a_59_75# sky130_fd_sc_hd__and4_1_0/VGND 0
C64 sky130_fd_sc_hd__and4_1_0/VGND sky130_fd_sc_hd__and4_1_0/B 0.04218f
C65 sky130_fd_sc_hd__and2_1_0/B sky130_fd_sc_hd__xor2_1_0/VPB 0
C66 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__xor2_1_0/X 0.00515f
C67 sky130_fd_sc_hd__xor2_1_0/B sky130_fd_sc_hd__and2_1_0/VPB 0.00406f
C68 sky130_fd_sc_hd__or2_1_0/a_150_297# sky130_fd_sc_hd__or4_1_0/C 0
C69 sky130_fd_sc_hd__or2_1_0/VPWR sky130_fd_sc_hd__xor2_1_0/X 0
C70 sky130_fd_sc_hd__or4_1_0/X sky130_fd_sc_hd__or4_1_0/A 0.00737f
C71 sky130_fd_sc_hd__and4_1_0/VGND sky130_fd_sc_hd__and2_1_4/VPWR 0
C72 a_195_n517# X 0.01091f
C73 sky130_fd_sc_hd__and2_1_0/A X 0.02789f
C74 sky130_fd_sc_hd__and4_1_1/A sky130_fd_sc_hd__and4_1_1/VPB 0
C75 sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__or2_1_0/A 0.12539f
C76 sky130_fd_sc_hd__and3_1_0/VGND sky130_fd_sc_hd__xor2_1_0/X 0
C77 sky130_fd_sc_hd__and4_1_1/C X 0.19117f
C78 sky130_fd_sc_hd__and2_1_5/a_59_75# sky130_fd_sc_hd__or4_1_0/B 0
C79 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__or4_1_0/B 0
C80 sky130_fd_sc_hd__and2_1_0/a_59_75# A 0
C81 sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__or2_1_0/VPWR -0.00376f
C82 sky130_fd_sc_hd__and4_1_1/a_27_47# X 0.04852f
C83 sky130_fd_sc_hd__or4_1_0/VPB X 0
C84 B a_155_n4715# 0
C85 a_69_n4715# VPB 0
C86 sky130_fd_sc_hd__or4_1_0/a_205_297# sky130_fd_sc_hd__or4_1_0/VGND -0
C87 a_19_n2185# B 0.00416f
C88 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__and4_1_0/a_109_47# 0
C89 sky130_fd_sc_hd__and2_1_5/a_59_75# B 0
C90 VPB sky130_fd_sc_hd__xor2_1_0/X 0
C91 B sky130_fd_sc_hd__and4_1_0/B 0.01591f
C92 sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__and3_1_0/VGND 0.00866f
C93 sky130_fd_sc_hd__and2_1_0/B X 0.00148f
C94 sky130_fd_sc_hd__or2_1_0/VGND sky130_fd_sc_hd__or4_1_0/C 0.00393f
C95 sky130_fd_sc_hd__or2_1_0/VGND sky130_fd_sc_hd__or2_1_0/a_150_297# -0
C96 a_195_n517# sky130_fd_sc_hd__xor2_1_0/B 0
C97 a_n63_n2185# a_19_n2185# -0
C98 sky130_fd_sc_hd__and2_1_5/VPWR X 0.25442f
C99 B sky130_fd_sc_hd__and2_1_4/VPWR 0
C100 sky130_fd_sc_hd__and2_1_0/A sky130_fd_sc_hd__xor2_1_0/B 0
C101 sky130_fd_sc_hd__and4_1_1/VGND X -0.0125f
C102 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and4_1_1/VPB 0.00112f
C103 sky130_fd_sc_hd__or2_1_0/a_68_297# sky130_fd_sc_hd__and3_1_0/VPWR 0
C104 sky130_fd_sc_hd__or4_1_0/VPWR sky130_fd_sc_hd__or4_1_0/VGND -0.0364f
C105 sky130_fd_sc_hd__or4_1_0/VPWR sky130_fd_sc_hd__or4_1_0/D -0.00384f
C106 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__and2_1_5/a_145_75# 0
C107 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__and3_1_0/VPWR 0
C108 a_27_n517# B 0.00416f
C109 sky130_fd_sc_hd__xor2_1_0/A sky130_fd_sc_hd__xor2_1_0/B 0.06504f
C110 B a_197_n3749# 0.00778f
C111 sky130_fd_sc_hd__and4_1_0/VPB a_67_n1483# 0
C112 sky130_fd_sc_hd__and3_1_0/VPB sky130_fd_sc_hd__xor2_1_0/X 0
C113 sky130_fd_sc_hd__and2_1_0/VPB sky130_fd_sc_hd__and4_1_1/A 0
C114 sky130_fd_sc_hd__or4_1_0/a_109_297# sky130_fd_sc_hd__or4_1_0/C 0
C115 sky130_fd_sc_hd__and2_1_0/a_145_75# X 0
C116 a_197_n3999# A 0.0022f
C117 sky130_fd_sc_hd__xor2_1_0/a_117_297# sky130_fd_sc_hd__xor2_1_0/B 0.00416f
C118 sky130_fd_sc_hd__and2_1_5/VPB sky130_fd_sc_hd__and4_1_1/A 0
C119 a_n63_n2185# a_197_n3749# 0
C120 sky130_fd_sc_hd__and2_1_5/VGND sky130_fd_sc_hd__and4_1_0/VPB 0.00281f
C121 sky130_fd_sc_hd__and4_1_0/VGND sky130_fd_sc_hd__xor2_1_0/X 0.03811f
C122 sky130_fd_sc_hd__and2_1_0/a_59_75# VPB 0.0016f
C123 sky130_fd_sc_hd__and2_1_0/B sky130_fd_sc_hd__xor2_1_0/B 0.00243f
C124 sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__or4_1_0/VGND 0.00146f
C125 sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__or4_1_0/D 0.00282f
C126 sky130_fd_sc_hd__and2_1_4/VGND X 0.06329f
C127 sky130_fd_sc_hd__and3_1_0/VGND A 0.00212f
C128 sky130_fd_sc_hd__and3_1_0/VPB sky130_fd_sc_hd__or2_1_0/B 0.01095f
C129 sky130_fd_sc_hd__and3_1_0/a_27_47# sky130_fd_sc_hd__and2_1_4/a_59_75# 0
C130 sky130_fd_sc_hd__or4_1_0/VPWR sky130_fd_sc_hd__and4_1_0/VPB 0
C131 sky130_fd_sc_hd__or2_1_0/VPWR sky130_fd_sc_hd__or2_1_0/A 0.15486f
C132 sky130_fd_sc_hd__and4_1_1/VGND sky130_fd_sc_hd__and4_1_1/VPB -0.0052f
C133 a_67_n1483# X 0.01753f
C134 sky130_fd_sc_hd__and3_1_0/a_27_47# sky130_fd_sc_hd__and3_1_0/VPWR -0.00561f
C135 sky130_fd_sc_hd__or4_1_0/VGND sky130_fd_sc_hd__or4_1_0/A 0.05672f
C136 sky130_fd_sc_hd__or4_1_0/D sky130_fd_sc_hd__or4_1_0/A 0.01787f
C137 a_195_n767# X 0
C138 sky130_fd_sc_hd__or4_1_0/a_27_297# sky130_fd_sc_hd__or4_1_0/B 0.00778f
C139 sky130_fd_sc_hd__or4_1_0/VPB sky130_fd_sc_hd__or4_1_0/C 0.00393f
C140 sky130_fd_sc_hd__or4_1_0/VGND sky130_fd_sc_hd__or2_1_0/a_68_297# 0
C141 sky130_fd_sc_hd__or2_1_0/a_68_297# sky130_fd_sc_hd__or4_1_0/D 0
C142 sky130_fd_sc_hd__or4_1_0/VGND sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C143 sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__and4_1_0/VGND 0.00665f
C144 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__or4_1_0/D 0.00126f
C145 sky130_fd_sc_hd__and2_1_5/VGND X 0.08784f
C146 sky130_fd_sc_hd__and2_1_0/A sky130_fd_sc_hd__and2_1_0/VPB 0.00109f
C147 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__or4_1_0/B 0.04167f
C148 VPB A 0.05774f
C149 sky130_fd_sc_hd__or4_1_0/D sky130_fd_sc_hd__and4_1_0/VPWR 0
C150 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__and4_1_1/VPWR 0.00963f
C151 sky130_fd_sc_hd__and4_1_1/a_109_47# X 0
C152 sky130_fd_sc_hd__xor2_1_0/A sky130_fd_sc_hd__and2_1_0/VPB 0.01565f
C153 a_69_n4715# B 0.06183f
C154 sky130_fd_sc_hd__xor2_1_0/a_35_297# sky130_fd_sc_hd__and4_1_0/B 0.00153f
C155 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and2_1_5/VPB 0.00946f
C156 sky130_fd_sc_hd__or4_1_0/a_277_297# sky130_fd_sc_hd__or4_1_0/VGND -0
C157 a_n53_n3749# X 0.00394f
C158 a_59_n3151# a_67_n1483# 0
C159 sky130_fd_sc_hd__and2_1_5/a_59_75# a_n55_n517# 0
C160 a_n55_n517# sky130_fd_sc_hd__and4_1_0/B 0.0065f
C161 B sky130_fd_sc_hd__xor2_1_0/X 0
C162 sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__or4_1_0/A 0
C163 sky130_fd_sc_hd__and2_1_5/VPB sky130_fd_sc_hd__and4_1_1/a_27_47# 0
C164 sky130_fd_sc_hd__and2_1_0/A sky130_fd_sc_hd__and4_1_1/A 0
C165 sky130_fd_sc_hd__and4_1_0/VPWR sky130_fd_sc_hd__and4_1_0/a_197_47# -0
C166 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and4_1_1/A 0.04301f
C167 sky130_fd_sc_hd__and2_1_0/B sky130_fd_sc_hd__and2_1_0/VPB 0.01331f
C168 sky130_fd_sc_hd__and4_1_1/a_27_47# sky130_fd_sc_hd__and4_1_1/A 0.00637f
C169 sky130_fd_sc_hd__or2_1_0/VPB X 0.00576f
C170 sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__and4_1_0/VPWR -0
C171 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and4_1_0/a_109_47# 0.00197f
C172 sky130_fd_sc_hd__and2_1_5/VPB sky130_fd_sc_hd__and2_1_5/VPWR -0.00635f
C173 sky130_fd_sc_hd__and2_1_4/VGND sky130_fd_sc_hd__or4_1_0/C 0.01004f
C174 sky130_fd_sc_hd__and4_1_0/VGND A 0.00151f
C175 sky130_fd_sc_hd__or4_1_0/A X 0.00572f
C176 sky130_fd_sc_hd__and2_1_5/VPB sky130_fd_sc_hd__and4_1_1/VGND 0
C177 a_n53_n3749# a_59_n3151# 0
C178 a_145_n3151# A 0.00152f
C179 sky130_fd_sc_hd__or2_1_0/a_68_297# X 0.0035f
C180 a_n63_n2185# sky130_fd_sc_hd__or2_1_0/B 0
C181 sky130_fd_sc_hd__or4_1_0/a_205_297# sky130_fd_sc_hd__or4_1_0/C 0
C182 sky130_fd_sc_hd__and4_1_0/a_27_47# X 0.06054f
C183 sky130_fd_sc_hd__xor2_1_0/a_285_297# sky130_fd_sc_hd__xor2_1_0/B 0.00746f
C184 sky130_fd_sc_hd__and2_1_5/VPWR sky130_fd_sc_hd__and4_1_1/A 0
C185 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__and4_1_0/VGND 0.06679f
C186 sky130_fd_sc_hd__and2_1_0/a_59_75# B 0
C187 sky130_fd_sc_hd__and4_1_1/VGND sky130_fd_sc_hd__and4_1_1/A -0.007f
C188 sky130_fd_sc_hd__and2_1_5/a_59_75# sky130_fd_sc_hd__and3_1_0/VPWR 0
C189 sky130_fd_sc_hd__and3_1_0/a_27_47# sky130_fd_sc_hd__and4_1_0/VPB 0
C190 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and3_1_0/VPWR 0
C191 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and2_1_0/A 0
C192 sky130_fd_sc_hd__and4_1_0/VPWR X 0.05837f
C193 sky130_fd_sc_hd__and2_1_0/A sky130_fd_sc_hd__xor2_1_0/A 0.00306f
C194 sky130_fd_sc_hd__and3_1_0/VPB sky130_fd_sc_hd__and3_1_0/VGND -0.00287f
C195 sky130_fd_sc_hd__and4_1_0/a_303_47# sky130_fd_sc_hd__and4_1_0/VPWR -0
C196 sky130_fd_sc_hd__or2_1_0/VPWR sky130_fd_sc_hd__and4_1_0/VGND 0.00285f
C197 sky130_fd_sc_hd__and3_1_0/a_109_47# sky130_fd_sc_hd__and3_1_0/VPWR -0
C198 sky130_fd_sc_hd__and2_1_4/a_59_75# sky130_fd_sc_hd__and2_1_4/VPWR -0.00137f
C199 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and4_1_1/a_27_47# 0.03795f
C200 sky130_fd_sc_hd__or4_1_0/VPWR sky130_fd_sc_hd__or4_1_0/C -0.00292f
C201 a_187_n2185# A 0
C202 sky130_fd_sc_hd__and2_1_0/B a_195_n517# 0
C203 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__or4_1_0/B 0.00147f
C204 sky130_fd_sc_hd__and2_1_0/B sky130_fd_sc_hd__and2_1_0/A 0.03965f
C205 sky130_fd_sc_hd__or2_1_0/a_68_297# sky130_fd_sc_hd__and4_1_1/VPB 0
C206 sky130_fd_sc_hd__and3_1_0/a_27_47# X 0.17069f
C207 B A 1.17029f
C208 sky130_fd_sc_hd__xor2_1_0/a_117_297# sky130_fd_sc_hd__xor2_1_0/A -0
C209 sky130_fd_sc_hd__and4_1_1/a_197_47# X 0
C210 sky130_fd_sc_hd__and2_1_0/B sky130_fd_sc_hd__xor2_1_0/A 0.19937f
C211 sky130_fd_sc_hd__or2_1_0/VPWR sky130_fd_sc_hd__or4_1_0/B 0
C212 sky130_fd_sc_hd__xor2_1_0/a_35_297# sky130_fd_sc_hd__xor2_1_0/X 0.0029f
C213 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and2_1_5/VPWR 0.072f
C214 sky130_fd_sc_hd__and2_1_5/VGND sky130_fd_sc_hd__and2_1_5/VPB -0.0046f
C215 a_n63_n2185# A 0.03465f
C216 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and4_1_1/VGND 0.19171f
C217 sky130_fd_sc_hd__or2_1_0/A B 0
C218 sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__or4_1_0/C 0.00412f
C219 a_n55_n517# sky130_fd_sc_hd__xor2_1_0/X 0
C220 X a_29_n3749# 0
C221 sky130_fd_sc_hd__and2_1_5/VPWR sky130_fd_sc_hd__and4_1_1/a_27_47# 0
C222 sky130_fd_sc_hd__and2_1_4/VPB X 0.03834f
C223 sky130_fd_sc_hd__and4_1_1/a_27_47# sky130_fd_sc_hd__and4_1_1/VGND -0.014f
C224 sky130_fd_sc_hd__or4_1_0/A sky130_fd_sc_hd__or4_1_0/C 0.18125f
C225 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and4_1_1/a_303_47# 0.00135f
C226 sky130_fd_sc_hd__xor2_1_0/VPB sky130_fd_sc_hd__and4_1_0/B 0
C227 sky130_fd_sc_hd__and2_1_0/A sky130_fd_sc_hd__and2_1_0/a_145_75# 0.00152f
C228 sky130_fd_sc_hd__or2_1_0/a_68_297# sky130_fd_sc_hd__or4_1_0/C 0.00324f
C229 sky130_fd_sc_hd__and4_1_1/VPWR sky130_fd_sc_hd__and4_1_1/a_303_47# -0
C230 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__or4_1_0/C 0
C231 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and4_1_0/a_197_47# 0.00195f
C232 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and4_1_0/a_109_47# 0
C233 a_195_n517# a_67_n1483# 0
C234 sky130_fd_sc_hd__and3_1_0/VPB sky130_fd_sc_hd__and4_1_0/VGND 0.00717f
C235 sky130_fd_sc_hd__and2_1_5/VPWR sky130_fd_sc_hd__and4_1_1/VGND 0.0025f
C236 sky130_fd_sc_hd__and2_1_0/A a_67_n1483# 0
C237 a_187_n2185# VPB -0
C238 sky130_fd_sc_hd__and2_1_5/a_59_75# sky130_fd_sc_hd__and4_1_0/VPB 0
C239 a_n63_n2185# sky130_fd_sc_hd__and3_1_0/VGND 0
C240 sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__and4_1_0/B 0.0108f
C241 sky130_fd_sc_hd__and2_1_0/a_59_75# sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.00144f
C242 sky130_fd_sc_hd__and2_1_4/VPB a_59_n3151# 0
C243 sky130_fd_sc_hd__xor2_1_0/a_285_47# sky130_fd_sc_hd__xor2_1_0/B -0
C244 sky130_fd_sc_hd__and2_1_4/a_59_75# sky130_fd_sc_hd__xor2_1_0/X 0
C245 VPB B 0.08228f
C246 sky130_fd_sc_hd__and2_1_0/a_59_75# a_n55_n517# 0
C247 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and3_1_0/VPWR 0
C248 sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__or2_1_0/VGND -0.00683f
C249 sky130_fd_sc_hd__or4_1_0/a_109_297# sky130_fd_sc_hd__or4_1_0/VPWR -0
C250 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and2_1_5/VGND 0.01061f
C251 sky130_fd_sc_hd__and3_1_0/a_27_47# sky130_fd_sc_hd__or4_1_0/C 0
C252 sky130_fd_sc_hd__and3_1_0/a_181_47# sky130_fd_sc_hd__and3_1_0/VPWR -0
C253 a_n63_n2185# VPB 0.00419f
C254 sky130_fd_sc_hd__or2_1_0/VGND sky130_fd_sc_hd__or4_1_0/A 0.01452f
C255 a_19_n2185# X 0
C256 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and4_1_1/a_109_47# 0.0023f
C257 sky130_fd_sc_hd__and2_1_5/VPB sky130_fd_sc_hd__and4_1_0/VPWR 0
C258 sky130_fd_sc_hd__and2_1_5/a_59_75# X 0.10648f
C259 sky130_fd_sc_hd__or2_1_0/VGND sky130_fd_sc_hd__or2_1_0/a_68_297# -0.00129f
C260 sky130_fd_sc_hd__and2_1_0/B a_67_n1483# 0
C261 sky130_fd_sc_hd__and4_1_0/B X 0.65102f
C262 sky130_fd_sc_hd__xor2_1_0/a_35_297# A 0
C263 sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__and3_1_0/VPWR 0.04682f
C264 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and4_1_0/a_303_47# 0
C265 sky130_fd_sc_hd__and3_1_0/a_109_47# X 0.0025f
C266 sky130_fd_sc_hd__and3_1_0/VPB B 0
C267 sky130_fd_sc_hd__or4_1_0/VPB sky130_fd_sc_hd__or4_1_0/VPWR -0.00543f
C268 a_n55_n517# A 0.03423f
C269 sky130_fd_sc_hd__xor2_1_0/a_285_297# sky130_fd_sc_hd__xor2_1_0/A -0
C270 sky130_fd_sc_hd__and2_1_4/VPB sky130_fd_sc_hd__or4_1_0/C 0.00887f
C271 X sky130_fd_sc_hd__and2_1_4/VPWR 0.13242f
C272 sky130_fd_sc_hd__or4_1_0/VGND sky130_fd_sc_hd__or4_1_0/a_27_297# -0.00274f
C273 sky130_fd_sc_hd__and2_1_5/VGND sky130_fd_sc_hd__and2_1_5/VPWR -0.03541f
C274 a_27_n517# X 0
C275 sky130_fd_sc_hd__and3_1_0/VPB a_n63_n2185# 0
C276 sky130_fd_sc_hd__or4_1_0/a_109_297# sky130_fd_sc_hd__or4_1_0/A 0.00223f
C277 sky130_fd_sc_hd__and4_1_0/VGND B 0
C278 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__or2_1_0/VPB 0
C279 X a_197_n3749# 0.01127f
C280 sky130_fd_sc_hd__and2_1_5/VPWR sky130_fd_sc_hd__and4_1_1/a_109_47# 0
C281 A sky130_fd_sc_hd__and4_1_0/a_109_47# 0
C282 sky130_fd_sc_hd__and2_1_0/B sky130_fd_sc_hd__xor2_1_0/a_285_297# 0
C283 sky130_fd_sc_hd__and4_1_1/a_109_47# sky130_fd_sc_hd__and4_1_1/VGND -0
C284 sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__and4_1_1/a_27_47# 0
C285 sky130_fd_sc_hd__and3_1_0/a_27_47# sky130_fd_sc_hd__or2_1_0/VGND 0
C286 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and4_1_1/VPB 0
C287 X sky130_fd_sc_hd__and2_1_5/a_145_75# 0.00203f
C288 sky130_fd_sc_hd__xor2_1_0/B sky130_fd_sc_hd__and4_1_0/B 0
C289 sky130_fd_sc_hd__xor2_1_0/VPB sky130_fd_sc_hd__xor2_1_0/X 0.00903f
C290 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__or2_1_0/a_68_297# 0
C291 a_59_n3151# sky130_fd_sc_hd__and2_1_4/VPWR 0
C292 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__and4_1_0/a_109_47# 0
C293 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C294 sky130_fd_sc_hd__and4_1_1/a_27_47# sky130_fd_sc_hd__or4_1_0/A 0
C295 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and4_1_0/a_197_47# 0.00123f
C296 sky130_fd_sc_hd__or4_1_0/VPB sky130_fd_sc_hd__or4_1_0/A 0.01474f
C297 sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__or4_1_0/a_27_297# 0
C298 sky130_fd_sc_hd__and4_1_1/a_27_47# sky130_fd_sc_hd__or2_1_0/a_68_297# 0
C299 sky130_fd_sc_hd__and2_1_4/a_59_75# A 0
C300 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and4_1_0/VPWR 0.01347f
C301 sky130_fd_sc_hd__or4_1_0/VPB sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C302 a_59_n3151# a_197_n3749# 0
C303 a_187_n2185# B 0.00766f
C304 sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__xor2_1_0/X 0.00937f
C305 sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__and4_1_1/VGND 0
C306 sky130_fd_sc_hd__xor2_1_0/a_35_297# VPB 0
C307 sky130_fd_sc_hd__or4_1_0/VPB sky130_fd_sc_hd__and4_1_0/VPWR 0
C308 a_n55_n517# VPB 0.00367f
C309 sky130_fd_sc_hd__or4_1_0/a_205_297# sky130_fd_sc_hd__or4_1_0/VPWR -0
C310 sky130_fd_sc_hd__or4_1_0/a_27_297# X 0
C311 sky130_fd_sc_hd__and4_1_1/VGND sky130_fd_sc_hd__or2_1_0/a_68_297# 0
C312 a_69_n4715# X 0
C313 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__and2_1_4/VPWR 0.01674f
C314 a_n63_n2185# B 0.04714f
C315 sky130_fd_sc_hd__and2_1_0/a_59_75# sky130_fd_sc_hd__xor2_1_0/VPB 0
C316 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and4_1_1/a_197_47# 0.00243f
C317 sky130_fd_sc_hd__xor2_1_0/X X 0.79943f
C318 sky130_fd_sc_hd__and3_1_0/VGND sky130_fd_sc_hd__and2_1_4/a_59_75# 0
C319 sky130_fd_sc_hd__and4_1_1/VPWR X -0.00415f
C320 sky130_fd_sc_hd__and3_1_0/VGND sky130_fd_sc_hd__and3_1_0/VPWR -0.03312f
C321 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and4_1_0/a_303_47# 0.00175f
C322 sky130_fd_sc_hd__and2_1_0/VPB sky130_fd_sc_hd__and4_1_0/B 0.00562f
C323 sky130_fd_sc_hd__and3_1_0/a_181_47# X 0.00275f
C324 sky130_fd_sc_hd__xor2_1_0/a_285_47# sky130_fd_sc_hd__xor2_1_0/A 0.0022f
C325 sky130_fd_sc_hd__and2_1_4/a_145_75# sky130_fd_sc_hd__and2_1_4/VPWR -0
C326 sky130_fd_sc_hd__and2_1_5/VPB sky130_fd_sc_hd__and4_1_0/B 0.00629f
C327 sky130_fd_sc_hd__or2_1_0/B X 0.09665f
C328 sky130_fd_sc_hd__xor2_1_0/VPB A 0
C329 sky130_fd_sc_hd__and2_1_4/a_59_75# VPB 0
C330 sky130_fd_sc_hd__or4_1_0/a_205_297# sky130_fd_sc_hd__or4_1_0/A 0.00121f
C331 a_69_n4715# a_59_n3151# 0
C332 VPB sky130_fd_sc_hd__and3_1_0/VPWR 0
C333 sky130_fd_sc_hd__or4_1_0/VGND sky130_fd_sc_hd__or2_1_0/A 0.00352f
C334 sky130_fd_sc_hd__and2_1_5/a_59_75# sky130_fd_sc_hd__and4_1_1/A 0
C335 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__or4_1_0/D 0.00173f
C336 sky130_fd_sc_hd__and4_1_1/A sky130_fd_sc_hd__and4_1_0/B 0
C337 sky130_fd_sc_hd__and2_1_5/VPWR sky130_fd_sc_hd__and4_1_1/a_197_47# 0
C338 A sky130_fd_sc_hd__and4_1_0/a_197_47# 0
C339 a_67_n1483# sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C340 sky130_fd_sc_hd__and4_1_1/a_197_47# sky130_fd_sc_hd__and4_1_1/VGND -0
C341 sky130_fd_sc_hd__or4_1_0/VGND sky130_fd_sc_hd__or2_1_0/VPWR 0
C342 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and4_1_1/VPB 0.02121f
C343 sky130_fd_sc_hd__or2_1_0/VPWR sky130_fd_sc_hd__or4_1_0/D 0.0035f
C344 sky130_fd_sc_hd__xor2_1_0/B sky130_fd_sc_hd__xor2_1_0/X 0.03047f
C345 a_67_n1483# sky130_fd_sc_hd__and4_1_0/VPWR 0
C346 sky130_fd_sc_hd__and4_1_1/VPWR sky130_fd_sc_hd__and4_1_1/VPB -0.0058f
C347 sky130_fd_sc_hd__and2_1_0/a_59_75# X 0.00215f
C348 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__and4_1_0/a_197_47# 0
C349 sky130_fd_sc_hd__or4_1_0/VPWR sky130_fd_sc_hd__or4_1_0/A 0.01499f
C350 sky130_fd_sc_hd__and3_1_0/VPB sky130_fd_sc_hd__and2_1_4/a_59_75# 0
C351 sky130_fd_sc_hd__or4_1_0/X sky130_fd_sc_hd__or4_1_0/B 0.00161f
C352 sky130_fd_sc_hd__and2_1_5/VGND sky130_fd_sc_hd__and4_1_0/VPWR 0.06986f
C353 sky130_fd_sc_hd__and3_1_0/VPB sky130_fd_sc_hd__and3_1_0/VPWR -0.00263f
C354 a_187_n2435# A 0.0022f
C355 sky130_fd_sc_hd__or4_1_0/a_27_297# sky130_fd_sc_hd__or4_1_0/C 0.03414f
C356 sky130_fd_sc_hd__or4_1_0/VPWR sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C357 sky130_fd_sc_hd__and3_1_0/a_27_47# sky130_fd_sc_hd__and2_1_4/VGND 0
C358 a_187_n2185# a_n55_n517# 0
C359 a_195_n517# sky130_fd_sc_hd__and4_1_0/B 0.00425f
C360 sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__or2_1_0/A 0.00385f
C361 sky130_fd_sc_hd__xor2_1_0/a_35_297# B 0
C362 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__and4_1_1/a_303_47# 0
C363 sky130_fd_sc_hd__or4_1_0/VPWR sky130_fd_sc_hd__and4_1_0/VPWR 0
C364 sky130_fd_sc_hd__and2_1_0/A sky130_fd_sc_hd__and4_1_0/B 0.03609f
C365 sky130_fd_sc_hd__and4_1_0/VGND sky130_fd_sc_hd__and2_1_4/a_59_75# 0
C366 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and2_1_5/a_59_75# 0.00218f
C367 a_n55_n517# B 0.04704f
C368 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and4_1_0/B 0
C369 sky130_fd_sc_hd__and4_1_0/VGND sky130_fd_sc_hd__and3_1_0/VPWR 0.123f
C370 A X 0.25089f
C371 sky130_fd_sc_hd__xor2_1_0/A sky130_fd_sc_hd__and4_1_0/B 0.00331f
C372 sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__or4_1_0/A 0.01132f
C373 sky130_fd_sc_hd__or4_1_0/a_277_297# sky130_fd_sc_hd__or4_1_0/VPWR -0
C374 sky130_fd_sc_hd__and4_1_0/a_303_47# A 0
C375 sky130_fd_sc_hd__and4_1_1/a_27_47# sky130_fd_sc_hd__and4_1_0/B 0
C376 sky130_fd_sc_hd__and2_1_4/VPB sky130_fd_sc_hd__and2_1_4/VGND -0.00451f
C377 a_n63_n2185# a_n55_n517# 0
C378 sky130_fd_sc_hd__and2_1_0/a_59_75# sky130_fd_sc_hd__xor2_1_0/B 0
C379 sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__and4_1_0/a_27_47# 0.00132f
C380 sky130_fd_sc_hd__or2_1_0/A X 0.04432f
C381 sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__or4_1_0/C 0.00406f
C382 sky130_fd_sc_hd__or2_1_0/a_68_297# sky130_fd_sc_hd__or4_1_0/A 0.00411f
C383 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__and4_1_0/a_303_47# 0
C384 sky130_fd_sc_hd__and2_1_0/B sky130_fd_sc_hd__and4_1_0/B 0.02591f
C385 sky130_fd_sc_hd__and2_1_0/VPB sky130_fd_sc_hd__xor2_1_0/X 0.00261f
C386 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__or4_1_0/A 0
C387 sky130_fd_sc_hd__or2_1_0/VPWR X 0.00738f
C388 sky130_fd_sc_hd__and2_1_0/VPB sky130_fd_sc_hd__and4_1_1/VPWR 0
C389 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__or2_1_0/a_68_297# 0
C390 sky130_fd_sc_hd__and2_1_5/VPWR sky130_fd_sc_hd__and2_1_5/a_59_75# -0.00969f
C391 sky130_fd_sc_hd__and2_1_5/VPWR sky130_fd_sc_hd__and4_1_0/B 0.00455f
C392 sky130_fd_sc_hd__and2_1_5/VPB sky130_fd_sc_hd__xor2_1_0/X 0.0094f
C393 sky130_fd_sc_hd__and4_1_0/VPWR sky130_fd_sc_hd__or4_1_0/A 0
C394 a_59_n3151# A 0.02803f
C395 sky130_fd_sc_hd__and2_1_5/a_59_75# sky130_fd_sc_hd__and4_1_1/VGND 0
C396 a_187_n2185# sky130_fd_sc_hd__and3_1_0/VPWR 0
C397 sky130_fd_sc_hd__and3_1_0/VGND X 0.1323f
C398 sky130_fd_sc_hd__xor2_1_0/B A 0
C399 sky130_fd_sc_hd__and2_1_4/a_59_75# B 0
C400 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__and4_1_0/VPWR -0
C401 sky130_fd_sc_hd__or4_1_0/a_277_297# sky130_fd_sc_hd__or4_1_0/A 0.00182f
C402 B sky130_fd_sc_hd__and3_1_0/VPWR 0.00199f
C403 sky130_fd_sc_hd__and4_1_0/VGND sky130_fd_sc_hd__or4_1_0/D 0
C404 sky130_fd_sc_hd__and4_1_1/A sky130_fd_sc_hd__xor2_1_0/X 0.03531f
C405 sky130_fd_sc_hd__and4_1_1/A sky130_fd_sc_hd__and4_1_1/VPWR -0.00839f
C406 sky130_fd_sc_hd__and2_1_0/a_145_75# sky130_fd_sc_hd__and4_1_0/B 0
C407 sky130_fd_sc_hd__and3_1_0/a_27_47# sky130_fd_sc_hd__or4_1_0/A 0
C408 a_n63_n2185# sky130_fd_sc_hd__and3_1_0/VPWR 0
C409 VPB X 0.07236f
C410 sky130_fd_sc_hd__and3_1_0/a_27_47# sky130_fd_sc_hd__or2_1_0/a_68_297# 0
C411 sky130_fd_sc_hd__and4_1_0/VGND sky130_fd_sc_hd__and4_1_0/a_197_47# -0
C412 sky130_fd_sc_hd__or2_1_0/VPWR sky130_fd_sc_hd__and4_1_1/VPB 0
C413 sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__or2_1_0/VGND 0.05365f
C414 sky130_fd_sc_hd__and3_1_0/a_27_47# sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C415 sky130_fd_sc_hd__or4_1_0/VGND sky130_fd_sc_hd__or4_1_0/B -0.00228f
C416 sky130_fd_sc_hd__and2_1_5/VPWR sky130_fd_sc_hd__and2_1_5/a_145_75# -0
C417 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__or4_1_0/D 0
C418 a_67_n1483# sky130_fd_sc_hd__and4_1_0/B 0.00159f
C419 sky130_fd_sc_hd__and3_1_0/a_27_47# sky130_fd_sc_hd__and4_1_0/VPWR 0
C420 a_195_n767# sky130_fd_sc_hd__and4_1_0/B 0
C421 sky130_fd_sc_hd__and2_1_4/VGND sky130_fd_sc_hd__and2_1_4/VPWR -0.02765f
C422 sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__and4_1_0/VGND -0.00404f
C423 sky130_fd_sc_hd__xor2_1_0/a_35_297# a_n55_n517# 0.00102f
C424 sky130_fd_sc_hd__and2_1_0/A sky130_fd_sc_hd__xor2_1_0/X 0
C425 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__or4_1_0/C 0.00317f
C426 sky130_fd_sc_hd__and2_1_5/VGND sky130_fd_sc_hd__and2_1_5/a_59_75# -0.00121f
C427 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__or2_1_0/a_150_297# 0.00183f
C428 sky130_fd_sc_hd__and2_1_5/VGND sky130_fd_sc_hd__and4_1_0/B 0.00461f
C429 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__xor2_1_0/X 0.1163f
C430 sky130_fd_sc_hd__and3_1_0/VPB X 0.0389f
C431 sky130_fd_sc_hd__and2_1_4/VPB sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C432 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and4_1_1/VPWR -0.00444f
C433 sky130_fd_sc_hd__xor2_1_0/A sky130_fd_sc_hd__xor2_1_0/X 0.03369f
C434 a_59_n3151# VPB 0.00186f
C435 sky130_fd_sc_hd__or2_1_0/VPWR sky130_fd_sc_hd__or4_1_0/C 0.00157f
C436 sky130_fd_sc_hd__and2_1_0/VPB A 0
C437 sky130_fd_sc_hd__or2_1_0/VPWR sky130_fd_sc_hd__or2_1_0/a_150_297# -0
C438 sky130_fd_sc_hd__and4_1_1/a_27_47# sky130_fd_sc_hd__xor2_1_0/X 0.12778f
C439 sky130_fd_sc_hd__or4_1_0/VPB sky130_fd_sc_hd__xor2_1_0/X 0
C440 a_153_n1483# A 0.00151f
C441 sky130_fd_sc_hd__xor2_1_0/VPB B 0
C442 sky130_fd_sc_hd__xor2_1_0/B VPB 0
C443 sky130_fd_sc_hd__and4_1_1/a_27_47# sky130_fd_sc_hd__and4_1_1/VPWR -0.01767f
C444 sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__or4_1_0/B 0
C445 sky130_fd_sc_hd__and4_1_0/VGND X 0.26798f
C446 sky130_fd_sc_hd__xor2_1_0/a_285_297# sky130_fd_sc_hd__and4_1_0/B 0
C447 sky130_fd_sc_hd__xor2_1_0/a_117_297# sky130_fd_sc_hd__xor2_1_0/X 0
C448 sky130_fd_sc_hd__and3_1_0/VGND sky130_fd_sc_hd__or4_1_0/C 0
C449 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__or2_1_0/B 0
C450 a_145_n3151# X 0
C451 sky130_fd_sc_hd__and4_1_0/VGND sky130_fd_sc_hd__and4_1_0/a_303_47# -0
C452 sky130_fd_sc_hd__and2_1_0/B sky130_fd_sc_hd__xor2_1_0/X 0.01218f
C453 sky130_fd_sc_hd__and2_1_5/VPWR sky130_fd_sc_hd__xor2_1_0/X 0.1083f
C454 sky130_fd_sc_hd__and2_1_0/a_59_75# a_195_n517# 0
C455 sky130_fd_sc_hd__and2_1_4/VPB sky130_fd_sc_hd__and3_1_0/a_27_47# 0
C456 sky130_fd_sc_hd__and4_1_0/VPB B 0
C457 sky130_fd_sc_hd__and4_1_1/VGND sky130_fd_sc_hd__xor2_1_0/X 0.04307f
C458 sky130_fd_sc_hd__and2_1_0/a_59_75# sky130_fd_sc_hd__and2_1_0/A 0.0274f
C459 sky130_fd_sc_hd__and4_1_1/VGND sky130_fd_sc_hd__and4_1_1/VPWR -0.04789f
C460 sky130_fd_sc_hd__or4_1_0/B X 0.00752f
C461 sky130_fd_sc_hd__or2_1_0/VGND sky130_fd_sc_hd__or2_1_0/A 0.0375f
C462 B a_187_n2435# 0
C463 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__and4_1_1/A 0
C464 sky130_fd_sc_hd__and2_1_0/a_59_75# sky130_fd_sc_hd__xor2_1_0/A 0
C465 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__or4_1_0/A 0
C466 a_187_n2185# X 0.01155f
C467 sky130_fd_sc_hd__or2_1_0/a_68_297# sky130_fd_sc_hd__and4_1_0/B 0
C468 sky130_fd_sc_hd__or2_1_0/VPWR sky130_fd_sc_hd__or2_1_0/VGND -0.03781f
C469 sky130_fd_sc_hd__and2_1_5/a_59_75# sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C470 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__and4_1_0/B 0.03791f
C471 sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__and4_1_1/VGND 0
C472 B X 0.38254f
C473 a_195_n517# A 0
C474 sky130_fd_sc_hd__and2_1_5/a_59_75# sky130_fd_sc_hd__and4_1_0/VPWR 0
C475 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and4_1_0/VPWR 0.0319f
C476 sky130_fd_sc_hd__and2_1_0/A A 0.00268f
C477 sky130_fd_sc_hd__and2_1_0/B sky130_fd_sc_hd__and2_1_0/a_59_75# 0.05693f
C478 sky130_fd_sc_hd__and3_1_0/VPB sky130_fd_sc_hd__or4_1_0/C 0
C479 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__and2_1_4/VPWR 0
C480 a_67_n1483# sky130_fd_sc_hd__xor2_1_0/X 0
C481 a_n63_n2185# X 0.01073f
C482 sky130_fd_sc_hd__or4_1_0/a_109_297# sky130_fd_sc_hd__or2_1_0/A 0
C483 sky130_fd_sc_hd__xor2_1_0/A A 0
C484 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__and4_1_1/VPB 0.00459f
C485 a_187_n2185# a_59_n3151# 0
C486 sky130_fd_sc_hd__and4_1_0/VGND sky130_fd_sc_hd__or4_1_0/C 0
C487 sky130_fd_sc_hd__or4_1_0/VPWR sky130_fd_sc_hd__or4_1_0/a_27_297# -0.01391f
C488 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__or2_1_0/A 0.00427f
C489 sky130_fd_sc_hd__and2_1_4/a_59_75# sky130_fd_sc_hd__and3_1_0/VPWR 0
C490 sky130_fd_sc_hd__and4_1_0/VGND sky130_fd_sc_hd__or2_1_0/a_150_297# 0
C491 sky130_fd_sc_hd__and2_1_5/VGND sky130_fd_sc_hd__xor2_1_0/X 0.11264f
C492 sky130_fd_sc_hd__and3_1_0/a_27_47# sky130_fd_sc_hd__and2_1_5/a_59_75# 0
C493 sky130_fd_sc_hd__and3_1_0/a_27_47# sky130_fd_sc_hd__and4_1_0/B 0
C494 a_59_n3151# B 0.05725f
C495 sky130_fd_sc_hd__and2_1_0/B A 0
C496 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__or2_1_0/VPWR 0
C497 sky130_fd_sc_hd__or4_1_0/VPB sky130_fd_sc_hd__or2_1_0/A 0
C498 sky130_fd_sc_hd__and4_1_1/a_109_47# sky130_fd_sc_hd__xor2_1_0/X 0
C499 a_69_n4715# a_n53_n3749# 0.00144f
C500 sky130_fd_sc_hd__or4_1_0/VPWR sky130_fd_sc_hd__xor2_1_0/X 0
C501 sky130_fd_sc_hd__xor2_1_0/B B 0
C502 sky130_fd_sc_hd__xor2_1_0/VPB a_n55_n517# 0
C503 sky130_fd_sc_hd__and4_1_1/a_109_47# sky130_fd_sc_hd__and4_1_1/VPWR -0
C504 sky130_fd_sc_hd__and3_1_0/a_27_47# sky130_fd_sc_hd__and2_1_4/VPWR 0
C505 sky130_fd_sc_hd__and4_1_1/a_27_47# sky130_fd_sc_hd__or2_1_0/VPWR 0
C506 sky130_fd_sc_hd__xor2_1_0/a_285_297# sky130_fd_sc_hd__xor2_1_0/X 0.0032f
C507 a_n63_n2185# a_59_n3151# 0.00144f
C508 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__or4_1_0/C 0.00801f
C509 sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__or4_1_0/a_27_297# 0
C510 sky130_fd_sc_hd__and3_1_0/VPB sky130_fd_sc_hd__or2_1_0/VGND 0.00189f
C511 sky130_fd_sc_hd__and2_1_0/a_59_75# a_67_n1483# 0
C512 sky130_fd_sc_hd__and4_1_1/VGND sky130_fd_sc_hd__or2_1_0/A 0.00602f
C513 sky130_fd_sc_hd__or4_1_0/a_27_297# sky130_fd_sc_hd__or4_1_0/A 0.11867f
C514 sky130_fd_sc_hd__and2_1_4/VPB sky130_fd_sc_hd__and2_1_4/VPWR -0
C515 sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__xor2_1_0/X 0
C516 sky130_fd_sc_hd__and2_1_0/A VPB 0.00317f
C517 sky130_fd_sc_hd__or4_1_0/a_27_297# sky130_fd_sc_hd__or2_1_0/a_68_297# 0
C518 B sky130_fd_sc_hd__or4_1_0/C 0
C519 sky130_fd_sc_hd__and4_1_1/VGND sky130_fd_sc_hd__or2_1_0/VPWR 0.02529f
C520 sky130_fd_sc_hd__or4_1_0/a_27_297# sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C521 sky130_fd_sc_hd__xor2_1_0/A VPB 0
C522 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__or4_1_0/A 0
C523 sky130_fd_sc_hd__xor2_1_0/a_35_297# X 0
C524 sky130_fd_sc_hd__or2_1_0/a_68_297# sky130_fd_sc_hd__xor2_1_0/X 0
C525 sky130_fd_sc_hd__and2_1_5/VPB sky130_fd_sc_hd__or4_1_0/B 0
C526 a_67_n1483# A 0.02856f
C527 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__xor2_1_0/X 0.03227f
C528 sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__or2_1_0/B 0.00342f
C529 a_n55_n517# X 0.00926f
C530 a_195_n767# A 0.0022f
C531 sky130_fd_sc_hd__xor2_1_0/a_285_297# sky130_fd_sc_hd__and2_1_0/a_59_75# 0
C532 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and4_1_0/VPWR 0.13704f
C533 sky130_fd_sc_hd__and2_1_0/VPB B 0.00364f
C534 sky130_fd_sc_hd__and2_1_0/B VPB 0.00134f
C535 sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__or4_1_0/A 0
C536 sky130_fd_sc_hd__and2_1_5/VGND A 0
C537 sky130_fd_sc_hd__and4_1_1/A sky130_fd_sc_hd__or4_1_0/B 0
C538 sky130_fd_sc_hd__and2_1_5/VPB B 0
C539 sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__or2_1_0/a_68_297# 0.00803f
C540 sky130_fd_sc_hd__and2_1_5/a_59_75# sky130_fd_sc_hd__and4_1_0/B 0.00451f
C541 sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C542 X sky130_fd_sc_hd__and4_1_0/a_109_47# 0.00198f
C543 a_n53_n3749# A 0.03479f
C544 sky130_fd_sc_hd__or4_1_0/VGND sky130_fd_sc_hd__or4_1_0/D -0
C545 sky130_fd_sc_hd__and3_1_0/a_27_47# sky130_fd_sc_hd__xor2_1_0/X 0
C546 sky130_fd_sc_hd__xor2_1_0/a_285_297# A 0
C547 sky130_fd_sc_hd__xor2_1_0/B sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.04603f
C548 sky130_fd_sc_hd__and4_1_1/a_197_47# sky130_fd_sc_hd__xor2_1_0/X 0
C549 sky130_fd_sc_hd__or4_1_0/VPWR sky130_fd_sc_hd__or2_1_0/A 0
C550 sky130_fd_sc_hd__xor2_1_0/B a_n55_n517# 0
C551 sky130_fd_sc_hd__and4_1_1/a_197_47# sky130_fd_sc_hd__and4_1_1/VPWR -0
C552 sky130_fd_sc_hd__and2_1_4/a_59_75# X 0.06657f
C553 a_27_n517# sky130_fd_sc_hd__and4_1_0/B 0
C554 X sky130_fd_sc_hd__and3_1_0/VPWR 0.34434f
C555 sky130_fd_sc_hd__xor2_1_0/a_285_47# sky130_fd_sc_hd__xor2_1_0/X 0
C556 sky130_fd_sc_hd__and2_1_4/VPB sky130_fd_sc_hd__xor2_1_0/X 0
C557 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__or4_1_0/B 0.00425f
C558 sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__and3_1_0/a_27_47# 0.00879f
C559 a_67_n1483# VPB 0.00126f
C560 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and2_1_5/a_145_75# 0
C561 a_195_n517# B 0.00754f
C562 sky130_fd_sc_hd__and4_1_1/a_27_47# sky130_fd_sc_hd__or4_1_0/B 0.00909f
C563 sky130_fd_sc_hd__or4_1_0/VPB sky130_fd_sc_hd__or4_1_0/B 0.01215f
C564 sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__or2_1_0/A 0.03627f
C565 sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__or4_1_0/D 0
C566 sky130_fd_sc_hd__and2_1_0/A B 0.13596f
C567 sky130_fd_sc_hd__and4_1_0/a_27_47# A 0
C568 sky130_fd_sc_hd__or4_1_0/X sky130_fd_sc_hd__or4_1_0/C 0.00286f
C569 sky130_fd_sc_hd__and2_1_5/VGND VPB 0
C570 sky130_fd_sc_hd__xor2_1_0/A B 0.01159f
C571 sky130_fd_sc_hd__and2_1_4/VPB sky130_fd_sc_hd__or2_1_0/B 0
C572 sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__or2_1_0/VPWR -0.00808f
C573 a_59_n3151# sky130_fd_sc_hd__and2_1_4/a_59_75# 0
C574 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__or4_1_0/A 0.04857f
C575 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__or2_1_0/a_68_297# 0.08751f
C576 sky130_fd_sc_hd__and2_1_5/VPWR sky130_fd_sc_hd__or4_1_0/B 0
C577 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__or2_1_0/A 0.00364f
C578 sky130_fd_sc_hd__or2_1_0/VPWR sky130_fd_sc_hd__or4_1_0/A 0.06282f
C579 sky130_fd_sc_hd__xor2_1_0/a_35_297# sky130_fd_sc_hd__and2_1_0/VPB 0.0035f
C580 a_n53_n3749# VPB 0.00422f
C581 sky130_fd_sc_hd__or4_1_0/VGND X 0
C582 sky130_fd_sc_hd__and4_1_1/VGND sky130_fd_sc_hd__or4_1_0/B 0.04642f
C583 sky130_fd_sc_hd__or4_1_0/D X 0
C584 sky130_fd_sc_hd__or2_1_0/VPWR sky130_fd_sc_hd__or2_1_0/a_68_297# -0.00741f
C585 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__and4_1_0/VPWR 0.00913f
C586 sky130_fd_sc_hd__or2_1_0/VPWR sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C587 sky130_fd_sc_hd__and2_1_0/B B 0.00168f
C588 a_n55_n517# sky130_fd_sc_hd__and2_1_0/VPB 0
C589 a_67_n1483# sky130_fd_sc_hd__and4_1_0/VGND 0
C590 sky130_fd_sc_hd__xor2_1_0/VPB X 0
C591 sky130_fd_sc_hd__and3_1_0/a_27_47# A 0.00153f
C592 sky130_fd_sc_hd__and2_1_5/VPB a_n55_n517# 0
C593 sky130_fd_sc_hd__and2_1_5/a_59_75# sky130_fd_sc_hd__xor2_1_0/X 0.03095f
C594 sky130_fd_sc_hd__and3_1_0/VGND sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C595 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__xor2_1_0/X 0.3542f
C596 X sky130_fd_sc_hd__and4_1_0/a_197_47# 0.00174f
C597 sky130_fd_sc_hd__and2_1_4/a_59_75# sky130_fd_sc_hd__or4_1_0/C 0.00834f
C598 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and4_1_1/VPWR 0
C599 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__and3_1_0/VPWR 0
C600 A a_29_n3749# -0
C601 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and2_1_4/VPWR 0
C602 sky130_fd_sc_hd__and4_1_0/VPB X 0.02141f
C603 a_69_n4715# a_197_n3749# 0
C604 sky130_fd_sc_hd__and4_1_0/a_27_47# VPB 0
C605 a_187_n2435# X 0
C606 a_187_n2185# a_67_n1483# 0
C607 VPB sky130_fd_sc_hd__and4_1_0/VPWR 0
C608 sky130_fd_sc_hd__and2_1_5/VGND sky130_fd_sc_hd__or4_1_0/B 0.00369f
C609 sky130_fd_sc_hd__and3_1_0/VGND sky130_fd_sc_hd__and3_1_0/a_27_47# -0.00436f
C610 sky130_fd_sc_hd__xor2_1_0/VPB sky130_fd_sc_hd__xor2_1_0/B 0.00802f
C611 a_195_n517# sky130_fd_sc_hd__xor2_1_0/a_35_297# 0
C612 a_67_n1483# B 0.05542f
C613 sky130_fd_sc_hd__and2_1_0/A sky130_fd_sc_hd__xor2_1_0/a_35_297# 0
C614 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and2_1_5/a_145_75# 0
C615 a_195_n517# a_n55_n517# 0
C616 sky130_fd_sc_hd__and4_1_1/a_109_47# sky130_fd_sc_hd__or4_1_0/B 0
C617 sky130_fd_sc_hd__or4_1_0/VPWR sky130_fd_sc_hd__or4_1_0/B 0.18661f
C618 sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__and4_1_0/VGND 0.00246f
C619 sky130_fd_sc_hd__and2_1_0/a_59_75# sky130_fd_sc_hd__and4_1_0/B 0.01295f
C620 sky130_fd_sc_hd__and2_1_0/A a_n55_n517# 0
C621 sky130_fd_sc_hd__xor2_1_0/A sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.03404f
C622 sky130_fd_sc_hd__and4_1_0/a_303_47# X 0.00226f
C623 a_n63_n2185# a_67_n1483# 0.00115f
C624 sky130_fd_sc_hd__and3_1_0/VPB sky130_fd_sc_hd__and4_1_0/a_27_47# 0.00142f
C625 sky130_fd_sc_hd__or4_1_0/VGND sky130_fd_sc_hd__or4_1_0/C 0.17252f
C626 sky130_fd_sc_hd__and4_1_1/C a_n55_n517# 0
C627 sky130_fd_sc_hd__or4_1_0/D sky130_fd_sc_hd__or4_1_0/C 0.02304f
C628 sky130_fd_sc_hd__or2_1_0/VGND sky130_fd_sc_hd__and3_1_0/VPWR 0.00385f
C629 sky130_fd_sc_hd__and3_1_0/a_27_47# VPB 0
C630 sky130_fd_sc_hd__and2_1_4/VPB sky130_fd_sc_hd__and3_1_0/VGND 0.00107f
C631 sky130_fd_sc_hd__xor2_1_0/A a_n55_n517# 0
C632 sky130_fd_sc_hd__and4_1_0/VGND sky130_fd_sc_hd__or2_1_0/a_68_297# 0.00157f
C633 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and4_1_1/a_303_47# 0.00124f
C634 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__and4_1_0/VGND -0.00307f
C635 A a_155_n4715# 0.00154f
C636 sky130_fd_sc_hd__and2_1_0/B sky130_fd_sc_hd__xor2_1_0/a_35_297# 0
C637 a_69_n4715# VNB 0.1752f
C638 a_n53_n3749# VNB 0.24712f
C639 a_59_n3151# VNB 0.17114f
C640 a_n63_n2185# VNB 0.24424f
C641 a_67_n1483# VNB 0.17003f
C642 a_n55_n517# VNB 0.24496f
C643 a_197_n3749# VNB 0.00137f
C644 a_195_n517# VNB 0.00137f
C645 sky130_fd_sc_hd__xor2_1_0/A VNB 0.45606f
C646 sky130_fd_sc_hd__xor2_1_0/B VNB 0.59565f
C647 sky130_fd_sc_hd__xor2_1_0/VPB VNB 0.69336f
C648 sky130_fd_sc_hd__xor2_1_0/a_285_297# VNB 0.00137f
C649 sky130_fd_sc_hd__xor2_1_0/a_35_297# VNB 0.25457f
C650 sky130_fd_sc_hd__and3_1_0/VGND VNB 0.30013f
C651 sky130_fd_sc_hd__or2_1_0/B VNB 0.46058f
C652 sky130_fd_sc_hd__and3_1_0/VPWR VNB 0.27425f
C653 sky130_fd_sc_hd__and3_1_0/VPB VNB 0.51617f
C654 sky130_fd_sc_hd__and3_1_0/a_27_47# VNB 0.17719f
C655 sky130_fd_sc_hd__or4_1_0/VGND VNB 0.36697f
C656 sky130_fd_sc_hd__or4_1_0/X VNB 0.08835f
C657 sky130_fd_sc_hd__or4_1_0/D VNB 0.17526f
C658 sky130_fd_sc_hd__or4_1_0/B VNB 0.82103f
C659 sky130_fd_sc_hd__or4_1_0/VPWR VNB 0.28998f
C660 sky130_fd_sc_hd__or4_1_0/VPB VNB 0.60476f
C661 sky130_fd_sc_hd__or4_1_0/a_27_297# VNB 0.16291f
C662 sky130_fd_sc_hd__and4_1_1/VGND VNB 0.39291f
C663 sky130_fd_sc_hd__and4_1_1/VPWR VNB 0.33454f
C664 sky130_fd_sc_hd__and4_1_1/A VNB 0.23645f
C665 sky130_fd_sc_hd__and4_1_1/VPB VNB 0.69336f
C666 sky130_fd_sc_hd__and4_1_1/a_27_47# VNB 0.17489f
C667 sky130_fd_sc_hd__and4_1_0/VGND VNB 0.39291f
C668 sky130_fd_sc_hd__or2_1_0/A VNB 0.322f
C669 sky130_fd_sc_hd__and4_1_0/VPWR VNB 0.33454f
C670 sky130_fd_sc_hd__xor2_1_0/X VNB 1.89172f
C671 sky130_fd_sc_hd__and4_1_0/B VNB 0.74819f
C672 sky130_fd_sc_hd__and4_1_0/VPB VNB 0.69336f
C673 sky130_fd_sc_hd__and4_1_0/a_27_47# VNB 0.17489f
C674 sky130_fd_sc_hd__or2_1_0/VGND VNB 0.32043f
C675 sky130_fd_sc_hd__or4_1_0/A VNB 0.45644f
C676 sky130_fd_sc_hd__or2_1_0/VPWR VNB 0.26856f
C677 sky130_fd_sc_hd__or2_1_0/VPB VNB 0.51617f
C678 sky130_fd_sc_hd__or2_1_0/a_68_297# VNB 0.15387f
C679 sky130_fd_sc_hd__and2_1_5/VGND VNB 0.3114f
C680 sky130_fd_sc_hd__and4_1_1/C VNB 0.33836f
C681 sky130_fd_sc_hd__and2_1_5/VPWR VNB 0.27345f
C682 sky130_fd_sc_hd__and2_1_5/VPB VNB 0.51617f
C683 sky130_fd_sc_hd__and2_1_5/a_59_75# VNB 0.17706f
C684 sky130_fd_sc_hd__and2_1_4/VGND VNB 0.3114f
C685 sky130_fd_sc_hd__or4_1_0/C VNB 1.46406f
C686 sky130_fd_sc_hd__and2_1_4/VPWR VNB 0.27345f
C687 sky130_fd_sc_hd__and2_1_4/VPB VNB 0.51617f
C688 sky130_fd_sc_hd__and2_1_4/a_59_75# VNB 0.17706f
C689 X VNB 5.38837f
C690 A VNB 2.72305f
C691 B VNB 2.14424f
C692 VPB VNB 3.62859f
C693 sky130_fd_sc_hd__and2_1_0/B VNB 0.2887f
C694 sky130_fd_sc_hd__and2_1_0/A VNB 0.39407f
C695 sky130_fd_sc_hd__and2_1_0/VPB VNB 0.51617f
C696 sky130_fd_sc_hd__and2_1_0/a_59_75# VNB 0.17706f
C697 a_187_n2185# VNB 0.00137f
.ends

.subckt sky130_fd_sc_hd__fa_1 A B CIN VGND VNB VPB VPWR COUT SUM a_1163_413# a_738_413#
+ a_1163_47# a_208_47# a_382_413# a_738_47# a_995_47# a_1091_47# a_76_199# a_1091_413#
+ a_382_47# a_208_413#
X0 a_76_199# B a_208_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=2268,138
X1 VGND A a_382_47# VNB sky130_fd_pr__nfet_01v8 ad=0.07384 pd=0.80236 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X2 a_738_413# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.07885 ps=0.80769 w=0.42 l=0.15
**devattr s=2268,138 d=2478,143
X3 a_1091_47# CIN a_995_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X4 VPWR CIN a_738_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07885 pd=0.80769 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X5 a_382_413# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.07885 ps=0.80769 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X6 a_1163_47# B a_1091_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X7 VPWR A a_382_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07885 pd=0.80769 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X8 a_995_47# a_76_199# a_738_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2772,150
X9 a_382_413# CIN a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X10 SUM a_995_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11427 ps=1.24175 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X11 a_208_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.07384 ps=0.80236 w=0.42 l=0.15
**devattr s=4094,199 d=2520,144
X12 VGND CIN a_738_47# VNB sky130_fd_pr__nfet_01v8 ad=0.07384 pd=0.80236 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X13 a_76_199# B a_208_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=2268,138
X14 a_208_413# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.07885 ps=0.80769 w=0.42 l=0.15
**devattr s=5914,269 d=2520,144
X15 a_738_413# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.07885 ps=0.80769 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X16 VGND A a_1163_47# VNB sky130_fd_pr__nfet_01v8 ad=0.07384 pd=0.80236 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=4094,199
X17 a_738_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.07384 ps=0.80236 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X18 a_738_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.07384 ps=0.80236 w=0.42 l=0.15
**devattr s=2268,138 d=2478,143
X19 a_1163_413# B a_1091_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X20 VPWR A a_1163_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07885 pd=0.80769 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=5914,269
X21 a_382_47# CIN a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X22 a_382_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.07384 ps=0.80236 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X23 SUM a_995_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.18773 ps=1.92308 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X24 a_995_47# a_76_199# a_738_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2772,150
X25 VPWR a_76_199# COUT VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18773 pd=1.92308 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X26 a_1091_413# CIN a_995_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X27 VGND a_76_199# COUT VNB sky130_fd_pr__nfet_01v8 ad=0.11427 pd=1.24175 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
C0 VGND SUM 0.07127f
C1 a_1163_47# SUM 0
C2 a_382_413# B 0.03303f
C3 VPB a_382_47# 0.00139f
C4 VPWR COUT 0.06663f
C5 A COUT 0.00345f
C6 VGND a_382_47# 0.14174f
C7 a_738_413# a_76_199# 0.00386f
C8 a_1163_413# a_738_413# 0
C9 a_738_413# a_995_47# 0.02283f
C10 B a_76_199# 0.13093f
C11 a_1163_413# B 0
C12 VPB CIN 0.23153f
C13 B a_995_47# 0.08206f
C14 VGND CIN 0.06042f
C15 A a_738_47# 0.04461f
C16 a_76_199# COUT 0.12975f
C17 a_1091_47# B 0
C18 B SUM 0.00111f
C19 VPWR a_1091_413# 0
C20 A VPWR 0.0705f
C21 B a_382_47# 0.01781f
C22 a_208_47# COUT 0
C23 a_738_413# CIN 0.07973f
C24 a_738_47# a_76_199# 0.03622f
C25 a_382_413# VPWR 0.15069f
C26 A a_382_413# 0.01121f
C27 B CIN 0.61202f
C28 a_738_47# a_995_47# 0.02301f
C29 VPB VGND 0.00519f
C30 a_1163_47# VGND 0.00175f
C31 a_76_199# VPWR 0.19016f
C32 a_76_199# a_1091_413# 0
C33 A a_76_199# 0.73176f
C34 a_738_47# a_1091_47# 0
C35 a_1163_413# VPWR 0
C36 a_995_47# VPWR 0.21287f
C37 a_1163_413# A 0
C38 a_995_47# a_1091_413# 0.00487f
C39 a_208_413# VPWR 0
C40 A a_995_47# 0.16271f
C41 A a_208_413# 0
C42 a_738_47# a_382_47# 0.00847f
C43 a_382_413# a_76_199# 0.03016f
C44 A a_1091_47# 0
C45 A a_208_47# 0
C46 VPWR SUM 0.07457f
C47 a_738_413# VPB 0.01092f
C48 A SUM 0.0054f
C49 VPB B 0.33717f
C50 A a_382_47# 0.04028f
C51 a_738_47# CIN 0.04534f
C52 B VGND 0.0456f
C53 a_995_47# a_76_199# 0.04882f
C54 a_1163_47# B 0
C55 a_208_413# a_76_199# 0.00682f
C56 a_1163_413# a_995_47# 0.00758f
C57 VPB COUT 0.01094f
C58 CIN VPWR 0.0577f
C59 a_1091_47# a_76_199# 0
C60 A CIN 0.45517f
C61 a_76_199# a_208_47# 0.00696f
C62 VGND COUT 0.05567f
C63 a_76_199# SUM 0
C64 a_1091_47# a_995_47# 0.00559f
C65 a_995_47# SUM 0.1439f
C66 a_76_199# a_382_47# 0.06611f
C67 a_382_413# CIN 0.08907f
C68 a_738_413# B 0.0177f
C69 VPB a_738_47# 0
C70 a_738_47# VGND 0.14671f
C71 CIN a_76_199# 0.21032f
C72 a_1163_47# a_738_47# 0
C73 CIN a_995_47# 0.05108f
C74 VPB VPWR 0.15613f
C75 A VPB 0.27513f
C76 B COUT 0
C77 VGND VPWR 0.04263f
C78 A VGND 0.10267f
C79 a_1163_47# A 0
C80 a_382_413# VPB 0.01154f
C81 CIN a_382_47# 0.03325f
C82 a_738_47# B 0.00556f
C83 VPB a_76_199# 0.10454f
C84 VGND a_76_199# 0.41492f
C85 VPB a_995_47# 0.05213f
C86 a_738_413# VPWR 0.14479f
C87 a_738_413# a_1091_413# 0
C88 A a_738_413# 0.01182f
C89 VGND a_995_47# 0.19875f
C90 a_1163_47# a_995_47# 0.00792f
C91 B VPWR 0.25287f
C92 B a_1091_413# 0
C93 A B 0.77269f
C94 a_1091_47# VGND 0
C95 VPB SUM 0.01793f
C96 a_382_413# a_738_413# 0.00985f
C97 VGND a_208_47# 0.00161f
C98 SUM VNB 0.10031f
C99 VGND VNB 0.81236f
C100 VPWR VNB 0.66922f
C101 COUT VNB 0.09411f
C102 CIN VNB 0.32537f
C103 B VNB 0.47131f
C104 A VNB 0.49582f
C105 VPB VNB 1.49072f
C106 a_738_47# VNB 0.01584f
C107 a_382_47# VNB 0.01578f
C108 a_738_413# VNB 0.00484f
C109 a_382_413# VNB 0.00345f
C110 a_995_47# VNB 0.1359f
C111 a_76_199# VNB 0.2795f
.ends

.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X a_505_21# a_535_374# a_439_47#
+ a_218_47# a_76_199# a_218_374#
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.08461 pd=0.79726 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.08461 ps=0.79726 w=0.42 l=0.15
**devattr s=2772,150 d=4704,280
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.08461 ps=0.79726 w=0.42 l=0.15
**devattr s=6334,279 d=3066,157
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.11336 pd=0.94775 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=5796,222
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=7728,268
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.11336 ps=0.94775 w=0.42 l=0.15
**devattr s=5796,222 d=4368,272
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
**devattr s=3990,179 d=2772,150
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
**devattr s=7728,268 d=1764,126
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=3990,179
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11336 ps=0.94775 w=0.42 l=0.15
**devattr s=4514,209 d=2772,150
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.20146 pd=1.89823 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=6334,279
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.17543 pd=1.46675 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4514,209
C0 A0 a_505_21# 0.03829f
C1 X a_76_199# 0.07764f
C2 a_76_199# A1 0.18667f
C3 X VPB 0.01205f
C4 A1 VPB 0.07208f
C5 VPWR a_76_199# 0.05421f
C6 a_439_47# A0 0.00369f
C7 a_535_374# a_76_199# 0
C8 VPWR VPB 0.10994f
C9 VGND a_218_47# 0.00328f
C10 VPWR X 0.12783f
C11 VPWR A1 0.01137f
C12 a_76_199# S 0.31816f
C13 a_76_199# VGND 0.16013f
C14 S VPB 0.16849f
C15 VGND VPB 0.01345f
C16 VPWR a_535_374# 0
C17 X S 0.00823f
C18 X VGND 0.05864f
C19 A1 S 0.08722f
C20 A1 VGND 0.07521f
C21 a_505_21# VPB 0.07806f
C22 VPWR S 0.39244f
C23 VPWR VGND 0.08036f
C24 a_535_374# S 0.00526f
C25 a_535_374# VGND 0
C26 A1 a_505_21# 0.09927f
C27 a_76_199# a_218_374# 0.00557f
C28 VPWR a_505_21# 0.08183f
C29 a_76_199# A0 0.05444f
C30 VGND S 0.03296f
C31 A0 VPB 0.1066f
C32 a_439_47# A1 0.00498f
C33 VPWR a_439_47# 0
C34 S a_505_21# 0.19751f
C35 A0 A1 0.2668f
C36 VGND a_505_21# 0.12387f
C37 VPWR a_218_374# 0.00177f
C38 VPWR A0 0.00732f
C39 a_439_47# VGND 0.00354f
C40 a_76_199# a_218_47# 0.00783f
C41 a_218_374# S 0.00688f
C42 VGND a_218_374# 0
C43 A0 S 0.03411f
C44 A0 VGND 0.04323f
C45 X a_218_47# 0
C46 a_76_199# VPB 0.04809f
C47 VPWR a_218_47# 0
C48 VGND VNB 0.49866f
C49 A1 VNB 0.14042f
C50 A0 VNB 0.13429f
C51 S VNB 0.26814f
C52 VPWR VNB 0.41925f
C53 X VNB 0.09236f
C54 VPB VNB 0.87055f
C55 a_505_21# VNB 0.24676f
C56 a_76_199# VNB 0.13947f
.ends

.subckt tt_um_ohmy90_adders clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5] ua[6]
+ ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0]
+ uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0]
+ uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0]
+ uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0]
+ uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7] VDPWR
Xsky130_fd_sc_hd__inv_1_4 sky130_fd_sc_hd__inv_1_4/A VDPWR VDPWR VDPWR VDPWR sky130_fd_sc_hd__inv_1_5/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_5 sky130_fd_sc_hd__inv_1_5/A VDPWR VDPWR VDPWR VDPWR sky130_fd_sc_hd__inv_1_6/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_6 sky130_fd_sc_hd__inv_1_6/A VDPWR VDPWR VDPWR VDPWR sky130_fd_sc_hd__inv_1_7/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_7 sky130_fd_sc_hd__inv_1_7/A VDPWR VDPWR VDPWR VDPWR sky130_fd_sc_hd__inv_1_8/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_8 sky130_fd_sc_hd__inv_1_8/A VDPWR VDPWR VDPWR VDPWR sky130_fd_sc_hd__inv_1_9/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_9 sky130_fd_sc_hd__inv_1_9/A VDPWR VDPWR VDPWR VDPWR sky130_fd_sc_hd__inv_1_9/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__mux4_1_0 VDPWR sky130_fd_sc_hd__inv_1_2/A sky130_fd_sc_hd__inv_1_0/A
+ sky130_fd_sc_hd__inv_1_1/A ui_in[0] ui_in[1] VDPWR VDPWR VDPWR VDPWR ua[0] sky130_fd_sc_hd__mux4_1_0/a_1290_413#
+ sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__mux4_1_0/a_1478_413# ui_in[1]
+ sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__mux4_1_0/a_923_363#
+ sky130_fd_sc_hd__mux4_1_0/a_193_47# sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__mux4_1_0/a_247_21#
+ sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__mux4_1_0/a_27_47#
+ sky130_fd_sc_hd__mux4_1
XCLA_0 CLA_0/sky130_fd_sc_hd__and4_1_1/a_303_47# VDPWR VDPWR VDPWR CLA_0/a_187_n2185#
+ CLA_0/sky130_fd_sc_hd__and4_1_0/a_27_47# CLA_0/sky130_fd_sc_hd__or2_1_0/a_150_297#
+ VDPWR CLA_0/sky130_fd_sc_hd__and2_1_5/a_59_75# VDPWR CLA_0/sky130_fd_sc_hd__and3_1_0/a_109_47#
+ VDPWR CLA_0/sky130_fd_sc_hd__and3_1_0/a_181_47# CLA_0/sky130_fd_sc_hd__xor2_1_0/a_285_297#
+ VDPWR CLA_0/sky130_fd_sc_hd__or4_1_0/B CLA_0/sky130_fd_sc_hd__or4_1_0/a_109_297#
+ VDPWR VDPWR VDPWR VDPWR CLA_0/sky130_fd_sc_hd__and3_1_0/a_27_47# CLA_0/a_187_n2435#
+ VDPWR VDPWR CLA_0/sky130_fd_sc_hd__xor2_1_0/a_285_47# CLA_0/a_19_n2185# CLA_0/sky130_fd_sc_hd__xor2_1_0/a_35_297#
+ CLA_0/sky130_fd_sc_hd__and2_1_4/a_145_75# CLA_0/sky130_fd_sc_hd__and2_1_0/a_145_75#
+ CLA_0/sky130_fd_sc_hd__and4_1_1/a_27_47# CLA_0/a_155_n4715# VDPWR CLA_0/sky130_fd_sc_hd__or4_1_0/A
+ VDPWR CLA_0/sky130_fd_sc_hd__or2_1_0/a_68_297# VDPWR CLA_0/a_195_n517# CLA_0/a_n63_n2185#
+ CLA_0/a_197_n3749# CLA_0/sky130_fd_sc_hd__or4_1_0/X CLA_0/sky130_fd_sc_hd__and4_1_0/a_109_47#
+ CLA_0/a_195_n767# CLA_0/a_197_n3999# VDPWR VDPWR VDPWR CLA_0/a_67_n1483# CLA_0/sky130_fd_sc_hd__and4_1_0/B
+ CLA_0/sky130_fd_sc_hd__and2_1_5/a_145_75# CLA_0/sky130_fd_sc_hd__and2_1_0/a_59_75#
+ VDPWR CLA_0/a_153_n1483# CLA_0/a_27_n517# CLA_0/a_69_n4715# CLA_0/sky130_fd_sc_hd__or2_1_0/B
+ CLA_0/sky130_fd_sc_hd__or2_1_0/A CLA_0/sky130_fd_sc_hd__or4_1_0/a_277_297# CLA_0/sky130_fd_sc_hd__and4_1_0/a_197_47#
+ VDPWR CLA_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# VDPWR CLA_0/sky130_fd_sc_hd__and4_1_0/a_303_47#
+ CLA_0/sky130_fd_sc_hd__and4_1_1/C CLA_0/sky130_fd_sc_hd__and4_1_1/a_109_47# VDPWR
+ CLA_0/sky130_fd_sc_hd__or4_1_0/a_27_297# CLA_0/a_29_n3749# VDPWR CLA_0/sky130_fd_sc_hd__or4_1_0/a_205_297#
+ CLA_0/sky130_fd_sc_hd__and2_1_4/a_59_75# VDPWR CLA_0/a_n53_n3749# CLA_0/a_n55_n517#
+ sky130_fd_sc_hd__inv_1_2/Y VDPWR VDPWR VDPWR CLA_0/sky130_fd_sc_hd__or4_1_0/C VDPWR
+ CLA_0/a_59_n3151# CLA_0/sky130_fd_sc_hd__xor2_1_0/X CLA_0/sky130_fd_sc_hd__and4_1_1/a_197_47#
+ VDPWR VDPWR VDPWR CLA_0/a_145_n3151# VDPWR CLA
XCLA_1 a_11777_15239# VDPWR VDPWR VDPWR a_9621_13111# a_11225_14223# a_11810_13649#
+ VDPWR a_10923_15189# VDPWR a_10923_12931# VDPWR a_10995_12931# a_9619_16343# VDPWR
+ CLA_1/sky130_fd_sc_hd__or4_1_0/B a_12697_14007# VDPWR VDPWR VDPWR VDPWR a_11165_13381#
+ a_9621_12861# VDPWR VDPWR a_9619_16093# a_9453_13111# a_9861_16543# a_10955_11939#
+ a_9577_15377# a_12009_15689# a_9589_10581# VDPWR CLA_1/sky130_fd_sc_hd__or4_1_0/A
+ VDPWR a_11949_13849# VDPWR a_9629_14779# a_9863_13311# a_9631_11547# sky130_fd_sc_hd__inv_1_2/A
+ a_10799_13773# a_9629_14529# a_9631_11297# VDPWR VDPWR VDPWR a_9749_14235# CLA_1/sky130_fd_sc_hd__and4_1_0/B
+ a_10761_14767# a_9739_15799# VDPWR a_9587_13813# a_9461_14779# a_9751_11003# CLA_1/sky130_fd_sc_hd__or2_1_0/B
+ CLA_1/sky130_fd_sc_hd__or2_1_0/A a_12865_14007# a_10887_13773# VDPWR a_9451_16343#
+ VDPWR a_10993_13773# CLA_1/sky130_fd_sc_hd__and4_1_1/C a_11583_15239# VDPWR a_13029_14207#
+ a_9463_11547# VDPWR a_12793_14007# a_11117_12361# VDPWR a_9873_11747# a_9871_14979#
+ CLA_0/sky130_fd_sc_hd__or4_1_0/X VDPWR VDPWR VDPWR CLA_1/sky130_fd_sc_hd__or4_1_0/C
+ VDPWR a_9741_12567# CLA_1/sky130_fd_sc_hd__xor2_1_0/X a_11671_15239# VDPWR VDPWR
+ VDPWR a_9579_12145# VDPWR CLA
Xsky130_fd_sc_hd__fa_1_0 VDPWR VDPWR sky130_fd_sc_hd__inv_1_0/Y VDPWR VDPWR VDPWR
+ VDPWR sky130_fd_sc_hd__fa_1_1/CIN sky130_fd_sc_hd__fa_1_0/SUM a_2049_1791# a_2313_1791#
+ a_2049_2157# a_3010_2157# a_2676_1791# a_2313_2157# a_1920_2241# a_2145_2157# a_3169_2241#
+ a_2145_1791# a_2676_2157# a_3010_1791# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_10 VDPWR VDPWR sky130_fd_sc_hd__inv_1_1/Y VDPWR VDPWR VDPWR
+ VDPWR sky130_fd_sc_hd__fa_1_8/CIN sky130_fd_sc_hd__fa_1_10/SUM a_2079_5051# a_2343_5051#
+ a_2079_5417# a_3040_5417# a_2706_5051# a_2343_5417# a_1950_5501# a_2175_5417# a_3199_5501#
+ a_2175_5051# a_2706_5417# a_3040_5051# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_1 VDPWR VDPWR sky130_fd_sc_hd__fa_1_1/CIN VDPWR VDPWR VDPWR
+ VDPWR sky130_fd_sc_hd__fa_1_2/CIN sky130_fd_sc_hd__fa_1_1/SUM a_4119_1787# a_4383_1787#
+ a_4119_2153# a_5080_2153# a_4746_1787# a_4383_2153# a_3990_2237# a_4215_2153# a_5239_2237#
+ a_4215_1787# a_4746_2153# a_5080_1787# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_11 VDPWR VDPWR sky130_fd_sc_hd__fa_1_9/COUT VDPWR VDPWR VDPWR
+ VDPWR sky130_fd_sc_hd__mux2_1_0/S sky130_fd_sc_hd__fa_1_11/SUM a_8167_5049# a_8431_5049#
+ a_8167_5415# a_9128_5415# a_8794_5049# a_8431_5415# a_8038_5499# a_8263_5415# a_9287_5499#
+ a_8263_5049# a_8794_5415# a_9128_5049# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_2 VDPWR VDPWR sky130_fd_sc_hd__fa_1_2/CIN VDPWR VDPWR VDPWR
+ VDPWR sky130_fd_sc_hd__fa_1_3/CIN sky130_fd_sc_hd__fa_1_2/SUM a_6071_1787# a_6335_1787#
+ a_6071_2153# a_7032_2153# a_6698_1787# a_6335_2153# a_5942_2237# a_6167_2153# a_7191_2237#
+ a_6167_1787# a_6698_2153# a_7032_1787# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_12 VDPWR VDPWR sky130_fd_sc_hd__fa_1_12/CIN VDPWR VDPWR VDPWR
+ VDPWR sky130_fd_sc_hd__fa_1_12/COUT sky130_fd_sc_hd__fa_1_12/SUM a_12323_5459# a_12587_5459#
+ a_12323_5825# a_13284_5825# a_12950_5459# a_12587_5825# a_12194_5909# a_12419_5825#
+ a_13443_5909# a_12419_5459# a_12950_5825# a_13284_5459# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_3 VDPWR VDPWR sky130_fd_sc_hd__fa_1_3/CIN VDPWR VDPWR VDPWR
+ VDPWR sky130_fd_sc_hd__fa_1_4/CIN sky130_fd_sc_hd__fa_1_3/SUM a_8073_1793# a_8337_1793#
+ a_8073_2159# a_9034_2159# a_8700_1793# a_8337_2159# a_7944_2243# a_8169_2159# a_9193_2243#
+ a_8169_1793# a_8700_2159# a_9034_1793# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_13 VDPWR VDPWR VDPWR VDPWR VDPWR VDPWR VDPWR sky130_fd_sc_hd__fa_1_12/CIN
+ sky130_fd_sc_hd__fa_1_13/SUM a_10261_5471# a_10525_5471# a_10261_5837# a_11222_5837#
+ a_10888_5471# a_10525_5837# a_10132_5921# a_10357_5837# a_11381_5921# a_10357_5471#
+ a_10888_5837# a_11222_5471# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_4 VDPWR VDPWR sky130_fd_sc_hd__fa_1_4/CIN VDPWR VDPWR VDPWR
+ VDPWR sky130_fd_sc_hd__fa_1_5/CIN sky130_fd_sc_hd__fa_1_4/SUM a_10025_1793# a_10289_1793#
+ a_10025_2159# a_10986_2159# a_10652_1793# a_10289_2159# a_9896_2243# a_10121_2159#
+ a_11145_2243# a_10121_1793# a_10652_2159# a_10986_1793# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_14 VDPWR VDPWR sky130_fd_sc_hd__fa_1_14/CIN VDPWR VDPWR VDPWR
+ VDPWR sky130_fd_sc_hd__fa_1_15/CIN sky130_fd_sc_hd__fa_1_14/SUM a_14281_5467# a_14545_5467#
+ a_14281_5833# a_15242_5833# a_14908_5467# a_14545_5833# a_14152_5917# a_14377_5833#
+ a_15401_5917# a_14377_5467# a_14908_5833# a_15242_5467# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_5 VDPWR VDPWR sky130_fd_sc_hd__fa_1_5/CIN VDPWR VDPWR VDPWR
+ VDPWR sky130_fd_sc_hd__fa_1_6/CIN sky130_fd_sc_hd__fa_1_5/SUM a_12017_1793# a_12281_1793#
+ a_12017_2159# a_12978_2159# a_12644_1793# a_12281_2159# a_11888_2243# a_12113_2159#
+ a_13137_2243# a_12113_1793# a_12644_2159# a_12978_1793# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_15 VDPWR VDPWR sky130_fd_sc_hd__fa_1_15/CIN VDPWR VDPWR VDPWR
+ VDPWR sky130_fd_sc_hd__mux2_1_0/A0 sky130_fd_sc_hd__fa_1_15/SUM a_16275_5473# a_16539_5473#
+ a_16275_5839# a_17236_5839# a_16902_5473# a_16539_5839# a_16146_5923# a_16371_5839#
+ a_17395_5923# a_16371_5473# a_16902_5839# a_17236_5473# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_6 VDPWR VDPWR sky130_fd_sc_hd__fa_1_6/CIN VDPWR VDPWR VDPWR
+ VDPWR sky130_fd_sc_hd__fa_1_7/CIN sky130_fd_sc_hd__fa_1_6/SUM a_13969_1793# a_14233_1793#
+ a_13969_2159# a_14930_2159# a_14596_1793# a_14233_2159# a_13840_2243# a_14065_2159#
+ a_15089_2243# a_14065_1793# a_14596_2159# a_14930_1793# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_16 VDPWR VDPWR sky130_fd_sc_hd__fa_1_16/CIN VDPWR VDPWR VDPWR
+ VDPWR sky130_fd_sc_hd__fa_1_18/CIN sky130_fd_sc_hd__fa_1_16/SUM a_12559_4553# a_12823_4553#
+ a_12559_4919# a_13520_4919# a_13186_4553# a_12823_4919# a_12430_5003# a_12655_4919#
+ a_13679_5003# a_12655_4553# a_13186_4919# a_13520_4553# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__inv_1_10 sky130_fd_sc_hd__inv_1_9/Y VDPWR VDPWR VDPWR VDPWR sky130_fd_sc_hd__inv_1_11/A
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__fa_1_7 VDPWR VDPWR sky130_fd_sc_hd__fa_1_7/CIN VDPWR VDPWR VDPWR
+ VDPWR sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__fa_1_7/SUM a_16033_1793# a_16297_1793#
+ a_16033_2159# a_16994_2159# a_16660_1793# a_16297_2159# a_15904_2243# a_16129_2159#
+ a_17153_2243# a_16129_1793# a_16660_2159# a_16994_1793# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_17 VDPWR VDPWR VDPWR VDPWR VDPWR VDPWR VDPWR sky130_fd_sc_hd__fa_1_16/CIN
+ sky130_fd_sc_hd__fa_1_17/SUM a_10289_4597# a_10553_4597# a_10289_4963# a_11250_4963#
+ a_10916_4597# a_10553_4963# a_10160_5047# a_10385_4963# a_11409_5047# a_10385_4597#
+ a_10916_4963# a_11250_4597# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__inv_1_0 sky130_fd_sc_hd__inv_1_0/A VDPWR VDPWR VDPWR VDPWR sky130_fd_sc_hd__inv_1_0/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_11 sky130_fd_sc_hd__inv_1_11/A VDPWR VDPWR VDPWR VDPWR VDPWR
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__fa_1_8 VDPWR VDPWR sky130_fd_sc_hd__fa_1_8/CIN VDPWR VDPWR VDPWR
+ VDPWR sky130_fd_sc_hd__fa_1_9/CIN sky130_fd_sc_hd__fa_1_8/SUM a_4213_5043# a_4477_5043#
+ a_4213_5409# a_5174_5409# a_4840_5043# a_4477_5409# a_4084_5493# a_4309_5409# a_5333_5493#
+ a_4309_5043# a_4840_5409# a_5174_5043# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__mux2_1_0 sky130_fd_sc_hd__mux2_1_0/A0 sky130_fd_sc_hd__mux2_1_0/A1
+ sky130_fd_sc_hd__mux2_1_0/S VDPWR VDPWR VDPWR VDPWR sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__mux2_1_0/a_505_21#
+ sky130_fd_sc_hd__mux2_1_0/a_535_374# sky130_fd_sc_hd__mux2_1_0/a_439_47# sky130_fd_sc_hd__mux2_1_0/a_218_47#
+ sky130_fd_sc_hd__mux2_1_0/a_76_199# sky130_fd_sc_hd__mux2_1_0/a_218_374# sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__fa_1_18 VDPWR VDPWR sky130_fd_sc_hd__fa_1_18/CIN VDPWR VDPWR VDPWR
+ VDPWR sky130_fd_sc_hd__fa_1_19/CIN sky130_fd_sc_hd__fa_1_18/SUM a_14561_4547# a_14825_4547#
+ a_14561_4913# a_15522_4913# a_15188_4547# a_14825_4913# a_14432_4997# a_14657_4913#
+ a_15681_4997# a_14657_4547# a_15188_4913# a_15522_4547# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__inv_1_1 sky130_fd_sc_hd__inv_1_1/A VDPWR VDPWR VDPWR VDPWR sky130_fd_sc_hd__inv_1_1/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__fa_1_9 VDPWR VDPWR sky130_fd_sc_hd__fa_1_9/CIN VDPWR VDPWR VDPWR
+ VDPWR sky130_fd_sc_hd__fa_1_9/COUT sky130_fd_sc_hd__fa_1_9/SUM a_6165_5043# a_6429_5043#
+ a_6165_5409# a_7126_5409# a_6792_5043# a_6429_5409# a_6036_5493# a_6261_5409# a_7285_5493#
+ a_6261_5043# a_6792_5409# a_7126_5043# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_19 VDPWR VDPWR sky130_fd_sc_hd__fa_1_19/CIN VDPWR VDPWR VDPWR
+ VDPWR sky130_fd_sc_hd__mux2_1_0/A1 sky130_fd_sc_hd__fa_1_19/SUM a_16583_4529# a_16847_4529#
+ a_16583_4895# a_17544_4895# a_17210_4529# a_16847_4895# a_16454_4979# a_16679_4895#
+ a_17703_4979# a_16679_4529# a_17210_4895# a_17544_4529# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__inv_1_2 sky130_fd_sc_hd__inv_1_2/A VDPWR VDPWR VDPWR VDPWR sky130_fd_sc_hd__inv_1_2/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_3 VDPWR VDPWR VDPWR VDPWR VDPWR sky130_fd_sc_hd__inv_1_4/A
+ sky130_fd_sc_hd__inv_1
C0 a_16371_5473# sky130_fd_sc_hd__inv_1_1/A 0
C1 rst_n clk 0.03102f
C2 VDPWR sky130_fd_sc_hd__fa_1_6/CIN 0.5584f
C3 a_7191_2237# sky130_fd_sc_hd__fa_1_3/SUM 0
C4 VDPWR sky130_fd_sc_hd__fa_1_19/SUM 0.08552f
C5 VDPWR a_10799_13773# 0.00164f
C6 a_16454_4979# a_17395_5923# 0
C7 VDPWR a_2313_1791# 0.01237f
C8 a_6429_5043# VDPWR 0.01623f
C9 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__mux4_1_0/a_193_47# 0
C10 sky130_fd_sc_hd__fa_1_5/CIN a_12644_2159# 0
C11 VDPWR a_2175_5417# 0.0011f
C12 sky130_fd_sc_hd__mux2_1_0/S sky130_fd_sc_hd__fa_1_12/CIN 0.05343f
C13 VDPWR sky130_fd_sc_hd__mux2_1_0/a_505_21# -0.01077f
C14 sky130_fd_sc_hd__fa_1_1/CIN a_2676_1791# 0
C15 VDPWR a_3010_2157# 0
C16 a_10916_4963# sky130_fd_sc_hd__inv_1_1/A 0
C17 VDPWR CLA_0/a_153_n1483# 0.00278f
C18 VDPWR a_14930_2159# 0
C19 a_9287_5499# VDPWR 0.08325f
C20 a_12194_5909# a_10525_5837# 0
C21 a_4383_2153# a_4215_2153# 0
C22 uo_out[5] uo_out[4] 0.03102f
C23 a_16679_4895# sky130_fd_sc_hd__inv_1_1/A 0
C24 a_16129_1793# sky130_fd_sc_hd__inv_1_0/A 0
C25 a_10993_13773# CLA_1/sky130_fd_sc_hd__or2_1_0/A 0
C26 sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__inv_1_1/A 0.01006f
C27 CLA_1/sky130_fd_sc_hd__xor2_1_0/X CLA_1/sky130_fd_sc_hd__and4_1_0/B -0.00923f
C28 a_12281_2159# sky130_fd_sc_hd__inv_1_0/A 0
C29 a_12950_5459# sky130_fd_sc_hd__fa_1_12/COUT 0
C30 a_12009_15689# a_11583_15239# 0
C31 VDPWR a_8073_2159# 0
C32 CLA_0/sky130_fd_sc_hd__and4_1_1/a_197_47# CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0
C33 a_12978_2159# sky130_fd_sc_hd__inv_1_0/A 0
C34 sky130_fd_sc_hd__fa_1_12/CIN sky130_fd_sc_hd__fa_1_16/CIN 0
C35 VDPWR a_13520_4553# 0
C36 sky130_fd_sc_hd__mux2_1_0/S a_17210_4895# 0
C37 CLA_1/sky130_fd_sc_hd__or4_1_0/B CLA_0/sky130_fd_sc_hd__or4_1_0/X 0.002f
C38 sky130_fd_sc_hd__fa_1_7/SUM a_17153_2243# -0
C39 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__inv_1_1/A -0
C40 VDPWR a_16994_2159# 0
C41 a_6429_5409# sky130_fd_sc_hd__inv_1_1/A 0
C42 sky130_fd_sc_hd__fa_1_5/CIN a_12113_1793# 0
C43 a_12655_4919# VDPWR 0.00109f
C44 a_14908_5467# a_16146_5923# 0
C45 a_15089_2243# a_13840_2243# -0.00146f
C46 uio_oe[4] uio_oe[3] 0.03102f
C47 VDPWR a_9873_11747# 0.12066f
C48 VDPWR CLA_0/sky130_fd_sc_hd__or4_1_0/a_109_297# 0
C49 a_16275_5473# sky130_fd_sc_hd__inv_1_1/A 0
C50 VDPWR a_17544_4529# 0
C51 a_11409_5047# sky130_fd_sc_hd__inv_1_1/A 0
C52 sky130_fd_sc_hd__fa_1_2/SUM a_5239_2237# 0
C53 sky130_fd_sc_hd__mux2_1_0/A1 sky130_fd_sc_hd__fa_1_19/CIN 0.00125f
C54 VDPWR sky130_fd_sc_hd__fa_1_18/SUM 0.0822f
C55 ua[0] sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.00698f
C56 a_5333_5493# sky130_fd_sc_hd__inv_1_1/Y 0.00303f
C57 sky130_fd_sc_hd__fa_1_15/CIN a_15401_5917# 0.00764f
C58 VDPWR a_11381_5921# 0.14577f
C59 CLA_0/sky130_fd_sc_hd__and4_1_1/C CLA_0/sky130_fd_sc_hd__and4_1_0/B -0
C60 CLA_1/sky130_fd_sc_hd__xor2_1_0/X a_9619_16093# 0
C61 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__inv_1_0/A 0.02727f
C62 VDPWR a_4477_5409# 0.0133f
C63 sky130_fd_sc_hd__inv_1_2/Y CLA_0/sky130_fd_sc_hd__or2_1_0/A 0
C64 CLA_0/sky130_fd_sc_hd__or4_1_0/X a_9739_15799# 0
C65 a_16994_1793# a_17153_2243# 0
C66 sky130_fd_sc_hd__inv_1_1/A a_10261_5471# 0
C67 uio_in[1] uio_in[0] 0.03102f
C68 uo_out[2] uo_out[3] 0.03102f
C69 a_16146_5923# sky130_fd_sc_hd__fa_1_19/CIN 0
C70 a_9861_16543# a_9871_14979# -0
C71 CLA_0/sky130_fd_sc_hd__and3_1_0/a_27_47# CLA_0/a_n63_n2185# -0
C72 a_12281_1793# sky130_fd_sc_hd__inv_1_0/A 0
C73 VDPWR sky130_fd_sc_hd__inv_1_11/A 0.49049f
C74 a_5333_5493# a_4084_5493# -0.00146f
C75 sky130_fd_sc_hd__inv_1_2/Y CLA_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0
C76 VDPWR CLA_0/sky130_fd_sc_hd__or4_1_0/C 0.71251f
C77 a_9287_5499# a_10888_5471# 0
C78 sky130_fd_sc_hd__fa_1_6/SUM sky130_fd_sc_hd__inv_1_0/A 0.00121f
C79 CLA_0/sky130_fd_sc_hd__or4_1_0/X VDPWR 2.79848f
C80 sky130_fd_sc_hd__mux2_1_0/a_76_199# sky130_fd_sc_hd__mux2_1_0/A1 0.00891f
C81 sky130_fd_sc_hd__fa_1_18/SUM sky130_fd_sc_hd__fa_1_18/CIN 0.05169f
C82 VDPWR sky130_fd_sc_hd__fa_1_13/SUM 0.12f
C83 sky130_fd_sc_hd__mux4_1_0/a_750_97# ui_in[0] 0.19136f
C84 VDPWR a_10525_5471# 0.01773f
C85 a_14432_4997# sky130_fd_sc_hd__inv_1_0/A 0
C86 sky130_fd_sc_hd__mux2_1_0/a_505_21# sky130_fd_sc_hd__mux2_1_0/A0 0.04199f
C87 VDPWR CLA_0/a_59_n3151# 0.06721f
C88 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__inv_1_0/A 0
C89 a_14908_5833# a_13443_5909# 0
C90 a_14377_5467# VDPWR 0
C91 sky130_fd_sc_hd__inv_1_11/A sky130_fd_sc_hd__inv_1_2/A 0
C92 a_9193_2243# sky130_fd_sc_hd__fa_1_4/SUM 0
C93 VDPWR sky130_fd_sc_hd__mux2_1_0/A1 0.29859f
C94 a_12823_4553# a_11409_5047# 0
C95 sky130_fd_sc_hd__inv_1_1/A a_8431_5049# 0
C96 a_6071_1787# sky130_fd_sc_hd__inv_1_0/Y 0
C97 a_5333_5493# a_6036_5493# 0.00419f
C98 CLA_0/sky130_fd_sc_hd__or4_1_0/X sky130_fd_sc_hd__inv_1_2/A 0.14763f
C99 a_14908_5833# sky130_fd_sc_hd__inv_1_1/A 0.0019f
C100 a_16902_5473# sky130_fd_sc_hd__fa_1_19/CIN 0
C101 sky130_fd_sc_hd__inv_1_2/Y CLA_0/sky130_fd_sc_hd__or4_1_0/B 0.002f
C102 a_11409_5047# a_10525_5837# 0
C103 a_3990_2237# VDPWR 0.04367f
C104 a_3199_5501# sky130_fd_sc_hd__inv_1_1/Y 0.04725f
C105 VDPWR CLA_0/sky130_fd_sc_hd__xor2_1_0/X 0.72048f
C106 a_12587_5459# a_13679_5003# 0
C107 a_12194_5909# a_12430_5003# 0
C108 a_17153_2243# a_15904_2243# -0.00146f
C109 ui_in[4] ui_in[3] 0.03102f
C110 a_6071_1787# sky130_fd_sc_hd__fa_1_2/CIN 0
C111 a_10289_4963# sky130_fd_sc_hd__inv_1_1/A 0
C112 a_12419_5825# a_12194_5909# -0
C113 ui_in[0] sky130_fd_sc_hd__mux4_1_0/a_193_413# 0.00324f
C114 a_5080_1787# sky130_fd_sc_hd__inv_1_0/Y 0
C115 a_9896_2243# sky130_fd_sc_hd__fa_1_4/SUM 0
C116 VDPWR a_16146_5923# 0.05018f
C117 sky130_fd_sc_hd__mux4_1_0/a_757_363# ui_in[0] 0.03011f
C118 ui_in[1] ui_in[2] 0.03102f
C119 VDPWR a_10385_4597# 0
C120 a_14432_4997# a_13679_5003# 0.00352f
C121 sky130_fd_sc_hd__inv_1_1/A a_17395_5923# 0.00779f
C122 a_16679_4529# sky130_fd_sc_hd__inv_1_0/A 0
C123 VDPWR a_14596_1793# 0.02482f
C124 sky130_fd_sc_hd__fa_1_9/COUT sky130_fd_sc_hd__fa_1_11/SUM 0.05168f
C125 a_11165_13381# CLA_1/sky130_fd_sc_hd__or4_1_0/C 0
C126 uo_out[1] uo_out[0] 0.03102f
C127 VDPWR a_9751_11003# 0.07777f
C128 sky130_fd_sc_hd__fa_1_7/CIN a_15089_2243# 0.00764f
C129 a_3199_5501# a_4084_5493# 0.00286f
C130 sky130_fd_sc_hd__fa_1_14/CIN a_15401_5917# 0.00155f
C131 VDPWR sky130_fd_sc_hd__mux4_1_0/a_923_363# 0
C132 sky130_fd_sc_hd__fa_1_7/SUM VDPWR 0.08423f
C133 a_8169_1793# sky130_fd_sc_hd__inv_1_0/A 0
C134 a_14545_5833# VDPWR 0.01394f
C135 a_10995_12931# VDPWR 0.00109f
C136 sky130_fd_sc_hd__mux4_1_0/a_1290_413# ua[0] 0.00191f
C137 VDPWR a_11145_2243# 0.07858f
C138 uio_oe[2] uio_oe[1] 0.03102f
C139 VDPWR sky130_fd_sc_hd__fa_1_12/CIN 0.60715f
C140 a_7032_2153# sky130_fd_sc_hd__inv_1_0/A 0
C141 sky130_fd_sc_hd__inv_1_0/Y a_4215_1787# 0
C142 VDPWR sky130_fd_sc_hd__inv_1_0/Y 1.17812f
C143 a_16902_5473# VDPWR 0.02626f
C144 VDPWR a_10652_1793# 0.02483f
C145 VDPWR sky130_fd_sc_hd__fa_1_2/CIN 0.56183f
C146 VDPWR sky130_fd_sc_hd__mux2_1_0/a_218_374# 0
C147 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__inv_1_1/A 0.04193f
C148 a_10916_4963# a_12430_5003# 0
C149 VDPWR a_14596_2159# 0.00628f
C150 a_14377_5833# a_14152_5917# -0
C151 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__fa_1_15/SUM 0.0031f
C152 CLA_0/sky130_fd_sc_hd__or4_1_0/A CLA_0/sky130_fd_sc_hd__and4_1_0/a_27_47# -0
C153 a_16994_1793# VDPWR 0
C154 VDPWR a_10289_4597# 0
C155 a_14545_5833# sky130_fd_sc_hd__fa_1_18/CIN 0
C156 a_8700_2159# a_9193_2243# 0
C157 a_16583_4895# sky130_fd_sc_hd__inv_1_1/A 0
C158 VDPWR a_4119_1787# 0
C159 sky130_fd_sc_hd__mux4_1_0/a_27_47# VDPWR 0.0141f
C160 a_8073_1793# VDPWR 0
C161 sky130_fd_sc_hd__fa_1_15/CIN sky130_fd_sc_hd__mux2_1_0/S 0.0454f
C162 a_12587_5825# sky130_fd_sc_hd__fa_1_12/CIN 0
C163 a_9861_16543# VDPWR 0.11156f
C164 VDPWR a_17210_4895# 0.00758f
C165 VDPWR sky130_fd_sc_hd__inv_1_6/A 0.26043f
C166 a_12113_2159# sky130_fd_sc_hd__inv_1_0/A 0
C167 a_16660_1793# a_17153_2243# 0
C168 a_12587_5459# sky130_fd_sc_hd__inv_1_1/A 0
C169 sky130_fd_sc_hd__mux2_1_0/S a_8794_5049# 0
C170 CLA_0/sky130_fd_sc_hd__and4_1_1/a_303_47# CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0
C171 a_12644_2159# sky130_fd_sc_hd__inv_1_0/A 0
C172 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__mux4_1_0/a_193_413# 0
C173 a_15681_4997# a_16454_4979# 0.00271f
C174 sky130_fd_sc_hd__mux2_1_0/S a_16847_4895# 0
C175 a_14432_4997# sky130_fd_sc_hd__inv_1_1/A 0
C176 ui_in[1] sky130_fd_sc_hd__mux4_1_0/a_834_97# 0.00187f
C177 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__inv_1_1/A 0.00117f
C178 sky130_fd_sc_hd__mux2_1_0/A1 sky130_fd_sc_hd__mux2_1_0/A0 0.13254f
C179 CLA_0/sky130_fd_sc_hd__and2_1_5/a_59_75# VDPWR 0.04034f
C180 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__inv_1_2/A 0.00494f
C181 VDPWR a_16660_2159# 0
C182 sky130_fd_sc_hd__inv_1_6/A sky130_fd_sc_hd__inv_1_2/A 0
C183 a_9861_16543# sky130_fd_sc_hd__inv_1_2/A 0
C184 a_6261_5409# sky130_fd_sc_hd__inv_1_1/A 0
C185 a_4746_2153# a_5239_2237# 0
C186 a_12559_4919# VDPWR 0
C187 a_16454_4979# a_17703_4979# -0.00146f
C188 a_9749_14235# a_9739_15799# -0
C189 VDPWR sky130_fd_sc_hd__inv_1_9/A 0.42927f
C190 a_14545_5467# a_16146_5923# 0
C191 sky130_fd_sc_hd__fa_1_14/SUM a_13443_5909# 0
C192 a_11117_12361# CLA_1/sky130_fd_sc_hd__or4_1_0/C 0
C193 a_13284_5459# sky130_fd_sc_hd__inv_1_1/A 0
C194 sky130_fd_sc_hd__fa_1_4/CIN a_11145_2243# 0.00156f
C195 sky130_fd_sc_hd__inv_1_1/A a_9128_5049# 0
C196 VDPWR CLA_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 0.07537f
C197 CLA_0/sky130_fd_sc_hd__and4_1_0/B CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0.00923f
C198 a_8038_5499# sky130_fd_sc_hd__inv_1_1/A 0.00209f
C199 a_17236_5839# sky130_fd_sc_hd__inv_1_1/A 0
C200 a_7191_2237# a_5942_2237# -0.00146f
C201 VDPWR a_15904_2243# 0.04328f
C202 a_2706_5417# sky130_fd_sc_hd__inv_1_1/Y 0.00245f
C203 a_11409_5047# a_12430_5003# 0.00138f
C204 VDPWR a_17210_4529# 0.02675f
C205 sky130_fd_sc_hd__fa_1_14/SUM sky130_fd_sc_hd__inv_1_1/A 0.00306f
C206 a_14233_2159# VDPWR 0.01296f
C207 a_16297_1793# sky130_fd_sc_hd__fa_1_7/CIN 0.00339f
C208 VDPWR a_7944_2243# 0.04373f
C209 sky130_fd_sc_hd__fa_1_3/CIN a_8169_1793# 0
C210 a_2049_2157# sky130_fd_sc_hd__inv_1_0/Y 0
C211 sky130_fd_sc_hd__fa_1_5/CIN ua[5] 0
C212 CLA_0/sky130_fd_sc_hd__and4_1_1/C CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0.00252f
C213 VDPWR a_9749_14235# 0.0678f
C214 sky130_fd_sc_hd__inv_1_9/A sky130_fd_sc_hd__inv_1_2/A 0
C215 a_10888_5471# sky130_fd_sc_hd__fa_1_12/CIN 0
C216 sky130_fd_sc_hd__fa_1_1/CIN a_4383_2153# 0
C217 a_15681_4997# sky130_fd_sc_hd__inv_1_0/A 0
C218 VDPWR a_2676_1791# 0.02874f
C219 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_0/a_27_413# -0
C220 sky130_fd_sc_hd__inv_1_1/A a_11222_5837# 0
C221 a_13137_2243# sky130_fd_sc_hd__fa_1_5/SUM -0
C222 a_2706_5417# a_4084_5493# 0
C223 CLA_0/sky130_fd_sc_hd__or2_1_0/a_68_297# VDPWR 0.03601f
C224 a_12113_1793# sky130_fd_sc_hd__inv_1_0/A 0
C225 a_17703_4979# sky130_fd_sc_hd__inv_1_0/A 0
C226 sky130_fd_sc_hd__fa_1_5/CIN sky130_fd_sc_hd__inv_1_0/A 0.00285f
C227 VDPWR a_8794_5415# 0.00688f
C228 a_11165_13381# a_11225_14223# -0
C229 VDPWR a_7032_1787# 0
C230 a_9287_5499# a_10525_5471# 0
C231 a_9287_5499# sky130_fd_sc_hd__fa_1_13/SUM 0
C232 sky130_fd_sc_hd__mux2_1_0/a_505_21# sky130_fd_sc_hd__mux2_1_0/A1 0.05261f
C233 sky130_fd_sc_hd__fa_1_9/COUT a_8431_5049# 0.0034f
C234 a_13029_14207# CLA_1/sky130_fd_sc_hd__or4_1_0/A -0.00166f
C235 sky130_fd_sc_hd__fa_1_15/CIN a_14908_5467# 0
C236 a_16902_5473# sky130_fd_sc_hd__mux2_1_0/A0 0
C237 VDPWR a_10357_5471# 0
C238 sky130_fd_sc_hd__mux2_1_0/S sky130_fd_sc_hd__fa_1_14/CIN 0.00543f
C239 sky130_fd_sc_hd__fa_1_12/COUT a_13443_5909# 0.00764f
C240 uio_out[2] uio_out[3] 0.03102f
C241 sky130_fd_sc_hd__fa_1_1/CIN a_3169_2241# 0.00987f
C242 VDPWR sky130_fd_sc_hd__fa_1_5/SUM 0.07924f
C243 sky130_fd_sc_hd__mux2_1_0/S a_10160_5047# 0
C244 VDPWR sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.04455f
C245 sky130_fd_sc_hd__fa_1_12/COUT sky130_fd_sc_hd__inv_1_1/A 0.00209f
C246 a_5333_5493# sky130_fd_sc_hd__fa_1_9/CIN 0.00764f
C247 a_3199_5501# a_4477_5043# 0
C248 sky130_fd_sc_hd__fa_1_12/CIN a_12419_5459# 0
C249 sky130_fd_sc_hd__fa_1_14/CIN a_14152_5917# 0.06747f
C250 sky130_fd_sc_hd__mux4_1_0/a_750_97# ua[0] 0
C251 a_12194_5909# sky130_fd_sc_hd__fa_1_12/SUM 0
C252 a_16539_5473# sky130_fd_sc_hd__fa_1_19/CIN 0
C253 a_9619_16343# CLA_1/sky130_fd_sc_hd__and4_1_0/B -0
C254 CLA_1/sky130_fd_sc_hd__or4_1_0/A a_12793_14007# -0
C255 a_8167_5415# sky130_fd_sc_hd__inv_1_1/A 0
C256 a_11409_5047# sky130_fd_sc_hd__fa_1_17/SUM -0
C257 VDPWR a_14281_5467# 0
C258 sky130_fd_sc_hd__fa_1_15/CIN sky130_fd_sc_hd__fa_1_19/CIN 0
C259 a_16660_1793# VDPWR 0.01926f
C260 a_12950_5825# a_13443_5909# 0
C261 sky130_fd_sc_hd__mux4_1_0/a_247_21# sky130_fd_sc_hd__inv_1_2/A -0
C262 a_14432_4997# a_13186_4919# 0
C263 VDPWR a_10553_4963# 0.00819f
C264 CLA_0/sky130_fd_sc_hd__or4_1_0/a_109_297# CLA_0/sky130_fd_sc_hd__or4_1_0/C 0
C265 a_16583_4529# sky130_fd_sc_hd__inv_1_0/A 0
C266 VDPWR a_14233_1793# 0.01623f
C267 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__mux2_1_0/a_218_47# 0
C268 a_11165_13381# CLA_1/sky130_fd_sc_hd__or2_1_0/B 0
C269 sky130_fd_sc_hd__mux2_1_0/S a_12194_5909# 0
C270 a_12950_5825# sky130_fd_sc_hd__inv_1_1/A 0.00186f
C271 a_8337_2159# a_7191_2237# 0
C272 sky130_fd_sc_hd__inv_1_0/Y a_2313_1791# 0.00463f
C273 a_16847_4895# sky130_fd_sc_hd__fa_1_19/CIN 0
C274 a_2706_5051# a_3199_5501# 0
C275 CLA_0/sky130_fd_sc_hd__and2_1_5/a_59_75# CLA_0/sky130_fd_sc_hd__and4_1_0/B -0.00106f
C276 ui_in[1] VDPWR 0.14712f
C277 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__fa_1_9/SUM 0.00121f
C278 a_14377_5833# VDPWR 0.00116f
C279 a_10923_12931# VDPWR 0.00209f
C280 CLA_1/sky130_fd_sc_hd__xor2_1_0/X a_11671_15239# -0
C281 a_3010_2157# sky130_fd_sc_hd__inv_1_0/Y 0
C282 a_11381_5921# sky130_fd_sc_hd__fa_1_13/SUM -0
C283 CLA_1/sky130_fd_sc_hd__or4_1_0/B CLA_1/sky130_fd_sc_hd__and4_1_1/C -0
C284 sky130_fd_sc_hd__inv_1_0/A a_12559_4553# 0
C285 VDPWR a_10887_13773# 0.00152f
C286 a_3040_5051# sky130_fd_sc_hd__inv_1_1/Y 0
C287 clk ena 0.03102f
C288 VDPWR CLA_0/a_197_n3999# 0.00312f
C289 CLA_0/sky130_fd_sc_hd__and2_1_0/a_59_75# CLA_0/sky130_fd_sc_hd__and4_1_0/B -0
C290 a_13029_14207# CLA_1/sky130_fd_sc_hd__or4_1_0/C -0
C291 sky130_fd_sc_hd__inv_1_1/A a_17236_5473# 0
C292 a_16539_5473# VDPWR 0.01782f
C293 CLA_0/sky130_fd_sc_hd__or4_1_0/X CLA_0/sky130_fd_sc_hd__or4_1_0/C 0
C294 ui_in[1] sky130_fd_sc_hd__inv_1_2/A 0
C295 VDPWR a_10289_1793# 0.01623f
C296 VDPWR sky130_fd_sc_hd__mux2_1_0/a_535_374# -0
C297 a_4213_5043# sky130_fd_sc_hd__fa_1_8/CIN 0
C298 a_12194_5909# sky130_fd_sc_hd__fa_1_16/CIN -0
C299 a_15681_4997# sky130_fd_sc_hd__inv_1_1/A 0
C300 sky130_fd_sc_hd__fa_1_15/CIN VDPWR 0.59373f
C301 a_11165_13381# CLA_1/sky130_fd_sc_hd__and4_1_0/B 0
C302 uo_out[4] uo_out[3] 0.03102f
C303 VDPWR a_8794_5049# 0.02595f
C304 VDPWR a_11250_4963# 0
C305 sky130_fd_sc_hd__inv_1_8/A sky130_fd_sc_hd__inv_1_5/A 0
C306 CLA_1/sky130_fd_sc_hd__or4_1_0/C a_12793_14007# -0
C307 sky130_fd_sc_hd__inv_1_1/A a_17703_4979# 0
C308 ua[6] sky130_fd_sc_hd__fa_1_3/CIN 0
C309 a_9034_2159# VDPWR 0
C310 VDPWR a_16847_4895# 0.01325f
C311 a_12017_2159# sky130_fd_sc_hd__inv_1_0/A 0
C312 CLA_1/sky130_fd_sc_hd__or4_1_0/A a_12865_14007# 0
C313 CLA_1/sky130_fd_sc_hd__and4_1_1/C VDPWR 0.26746f
C314 a_14233_2159# sky130_fd_sc_hd__fa_1_6/CIN 0
C315 a_6698_2153# sky130_fd_sc_hd__inv_1_0/A 0
C316 a_6698_1787# sky130_fd_sc_hd__inv_1_0/A 0
C317 sky130_fd_sc_hd__fa_1_12/CIN a_11381_5921# 0.00989f
C318 a_8038_5499# sky130_fd_sc_hd__fa_1_9/COUT 0.06773f
C319 sky130_fd_sc_hd__fa_1_15/CIN sky130_fd_sc_hd__fa_1_18/CIN 0
C320 VDPWR sky130_fd_sc_hd__mux2_1_0/a_439_47# -0
C321 VDPWR a_15089_2243# 0.07798f
C322 CLA_1/sky130_fd_sc_hd__or4_1_0/B CLA_1/sky130_fd_sc_hd__or4_1_0/A -0.00383f
C323 sky130_fd_sc_hd__fa_1_1/CIN a_5239_2237# 0.00156f
C324 sky130_fd_sc_hd__inv_1_2/Y VDPWR 1.77772f
C325 a_5942_2237# a_5239_2237# 0.00419f
C326 a_10132_5921# sky130_fd_sc_hd__inv_1_1/A 0.00451f
C327 sky130_fd_sc_hd__inv_1_9/Y VDPWR 0.38927f
C328 sky130_fd_sc_hd__inv_1_1/A a_7285_5493# 0.00299f
C329 a_16129_1793# sky130_fd_sc_hd__fa_1_7/CIN 0
C330 a_16902_5839# sky130_fd_sc_hd__inv_1_1/A 0.00192f
C331 a_14065_2159# VDPWR 0.00104f
C332 a_6429_5409# sky130_fd_sc_hd__fa_1_9/CIN 0
C333 sky130_fd_sc_hd__fa_1_1/CIN sky130_fd_sc_hd__fa_1_1/SUM 0.05108f
C334 VDPWR sky130_fd_sc_hd__fa_1_0/SUM 0.09642f
C335 a_11810_13649# VDPWR 0
C336 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__inv_1_2/A 0.05987f
C337 a_10289_1793# sky130_fd_sc_hd__fa_1_4/CIN 0.00339f
C338 a_15401_5917# sky130_fd_sc_hd__fa_1_15/SUM 0
C339 sky130_fd_sc_hd__inv_1_1/A a_10888_5837# 0.00192f
C340 uio_in[0] ui_in[7] 0.03102f
C341 sky130_fd_sc_hd__inv_1_9/Y sky130_fd_sc_hd__inv_1_2/A 0
C342 a_12950_5459# sky130_fd_sc_hd__inv_1_1/A 0
C343 sky130_fd_sc_hd__mux2_1_0/S a_11409_5047# 0
C344 a_4383_1787# a_5239_2237# 0.00112f
C345 a_9287_5499# a_8794_5415# 0
C346 a_14561_4547# sky130_fd_sc_hd__inv_1_0/A 0
C347 a_16454_4979# sky130_fd_sc_hd__inv_1_0/A 0
C348 VDPWR a_15242_5467# 0
C349 VDPWR sky130_fd_sc_hd__fa_1_14/CIN 0.48033f
C350 CLA_1/sky130_fd_sc_hd__or4_1_0/B a_12009_15689# -0
C351 VDPWR CLA_0/a_n53_n3749# 0.11836f
C352 VDPWR a_10160_5047# 0.09998f
C353 sky130_fd_sc_hd__mux2_1_0/a_218_374# sky130_fd_sc_hd__mux2_1_0/A1 0
C354 a_3990_2237# sky130_fd_sc_hd__inv_1_0/Y 0.00211f
C355 VDPWR CLA_0/sky130_fd_sc_hd__or4_1_0/a_205_297# 0
C356 CLA_1/sky130_fd_sc_hd__or4_1_0/A VDPWR 0.5569f
C357 a_12323_5459# sky130_fd_sc_hd__inv_1_1/A 0
C358 CLA_0/sky130_fd_sc_hd__or4_1_0/X a_9861_16543# 0.00257f
C359 a_14432_4997# a_15401_5917# 0
C360 a_5333_5493# VDPWR 0.08029f
C361 a_13029_14207# a_12697_14007# -0
C362 a_13186_4553# sky130_fd_sc_hd__inv_1_0/A 0
C363 sky130_fd_sc_hd__fa_1_15/CIN sky130_fd_sc_hd__mux2_1_0/A0 0
C364 sky130_fd_sc_hd__fa_1_6/CIN a_14233_1793# 0.00339f
C365 a_11409_5047# sky130_fd_sc_hd__fa_1_16/CIN 0.01033f
C366 CLA_1/sky130_fd_sc_hd__or4_1_0/B CLA_1/sky130_fd_sc_hd__or4_1_0/C -0
C367 a_17210_4895# sky130_fd_sc_hd__mux2_1_0/A1 0
C368 VDPWR sky130_fd_sc_hd__fa_1_4/SUM 0.07933f
C369 sky130_fd_sc_hd__inv_1_1/Y sky130_fd_sc_hd__fa_1_8/CIN 0.00478f
C370 sky130_fd_sc_hd__inv_1_9/A sky130_fd_sc_hd__inv_1_11/A 0
C371 a_13029_14207# a_11225_14223# -0
C372 CLA_1/sky130_fd_sc_hd__or4_1_0/A sky130_fd_sc_hd__inv_1_2/A 0.0262f
C373 sky130_fd_sc_hd__fa_1_18/CIN sky130_fd_sc_hd__fa_1_14/CIN 0.00111f
C374 a_6698_1787# sky130_fd_sc_hd__fa_1_3/CIN 0
C375 sky130_fd_sc_hd__fa_1_14/SUM a_15401_5917# -0
C376 VDPWR a_7191_2237# 0.07989f
C377 VDPWR a_12194_5909# 0.05145f
C378 VDPWR a_15242_5833# 0
C379 a_9287_5499# a_10553_4963# 0
C380 a_16297_1793# VDPWR 0.0162f
C381 VDPWR sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.00538f
C382 a_6071_2153# VDPWR 0
C383 VDPWR a_10385_4963# 0.00101f
C384 uo_out[0] uio_in[7] 0.03102f
C385 VDPWR a_14065_1793# 0
C386 a_4084_5493# sky130_fd_sc_hd__fa_1_8/CIN 0.06766f
C387 sky130_fd_sc_hd__mux2_1_0/a_439_47# sky130_fd_sc_hd__mux2_1_0/A0 0.00191f
C388 VDPWR a_4383_2153# 0.01313f
C389 VDPWR a_6335_1787# 0.01622f
C390 CLA_0/sky130_fd_sc_hd__or4_1_0/X a_9749_14235# 0.00137f
C391 VDPWR a_12009_15689# 0.06139f
C392 a_11949_13849# CLA_1/sky130_fd_sc_hd__or4_1_0/A 0
C393 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__fa_1_2/CIN 0.00133f
C394 a_12017_1793# VDPWR 0
C395 CLA_0/sky130_fd_sc_hd__and2_1_5/a_59_75# CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0
C396 a_14281_5833# VDPWR 0
C397 ui_in[0] sky130_fd_sc_hd__inv_1_0/A 0.0357f
C398 a_13679_5003# sky130_fd_sc_hd__inv_1_0/A 0
C399 sky130_fd_sc_hd__inv_1_2/Y CLA_0/sky130_fd_sc_hd__and4_1_0/B 0
C400 a_17210_4529# sky130_fd_sc_hd__mux2_1_0/A1 0
C401 a_11222_5471# sky130_fd_sc_hd__inv_1_1/A 0
C402 uio_oe[1] uio_oe[0] 0.03102f
C403 sky130_fd_sc_hd__fa_1_15/CIN sky130_fd_sc_hd__fa_1_19/SUM 0
C404 sky130_fd_sc_hd__mux2_1_0/S a_17395_5923# 0
C405 sky130_fd_sc_hd__fa_1_10/SUM a_3199_5501# -0
C406 CLA_0/sky130_fd_sc_hd__or2_1_0/a_68_297# CLA_0/sky130_fd_sc_hd__or4_1_0/C -0
C407 VDPWR a_3199_5501# 0.0764f
C408 VDPWR sky130_fd_sc_hd__fa_1_11/SUM 0.07928f
C409 sky130_fd_sc_hd__inv_1_2/Y CLA_0/sky130_fd_sc_hd__and4_1_1/C 0.05432f
C410 CLA_0/sky130_fd_sc_hd__and2_1_0/a_59_75# CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0
C411 sky130_fd_sc_hd__inv_1_0/Y a_4119_1787# 0
C412 CLA_1/sky130_fd_sc_hd__or4_1_0/C VDPWR 0.70748f
C413 sky130_fd_sc_hd__inv_1_0/A a_8700_1793# 0
C414 a_16371_5473# VDPWR 0
C415 VDPWR a_10121_1793# 0
C416 a_13029_14207# CLA_1/sky130_fd_sc_hd__or2_1_0/A 0
C417 a_1950_5501# sky130_fd_sc_hd__inv_1_1/Y 0.03136f
C418 VDPWR a_3169_2241# 0.07686f
C419 sky130_fd_sc_hd__fa_1_12/COUT a_15401_5917# 0
C420 VDPWR sky130_fd_sc_hd__mux4_1_0/a_193_47# 0
C421 sky130_fd_sc_hd__inv_1_1/Y a_2079_5417# 0
C422 a_5333_5493# sky130_fd_sc_hd__fa_1_8/SUM -0
C423 a_16539_5839# sky130_fd_sc_hd__inv_1_1/A 0.00117f
C424 a_14545_5467# sky130_fd_sc_hd__fa_1_14/CIN 0.00339f
C425 a_11777_15239# VDPWR 0.00104f
C426 a_11888_2243# a_13137_2243# -0.00146f
C427 VDPWR a_10916_4963# 0.00686f
C428 CLA_1/sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__inv_1_2/A 0
C429 sky130_fd_sc_hd__fa_1_4/CIN sky130_fd_sc_hd__fa_1_4/SUM 0.05218f
C430 a_15089_2243# sky130_fd_sc_hd__fa_1_6/CIN 0.00156f
C431 a_8700_2159# VDPWR 0.00623f
C432 sky130_fd_sc_hd__inv_1_1/A a_16454_4979# 0
C433 a_8167_5049# sky130_fd_sc_hd__inv_1_1/A 0
C434 VDPWR a_16679_4895# 0.00127f
C435 a_11949_13849# a_12009_15689# 0
C436 sky130_fd_sc_hd__fa_1_9/CIN sky130_fd_sc_hd__fa_1_9/SUM 0.05218f
C437 VDPWR a_12644_1793# 0.02483f
C438 VDPWR sky130_fd_sc_hd__mux4_1_0/a_668_97# 0.00566f
C439 a_16847_4529# sky130_fd_sc_hd__fa_1_19/CIN 0.00339f
C440 sky130_fd_sc_hd__inv_1_8/A sky130_fd_sc_hd__inv_1_7/A 0.05599f
C441 sky130_fd_sc_hd__fa_1_3/CIN sky130_fd_sc_hd__inv_1_0/A 0.00286f
C442 VDPWR a_11888_2243# 0.0435f
C443 sky130_fd_sc_hd__fa_1_9/COUT a_7285_5493# 0.00764f
C444 CLA_1/sky130_fd_sc_hd__or4_1_0/C a_11949_13849# -0
C445 a_8431_5415# a_10132_5921# 0
C446 CLA_1/sky130_fd_sc_hd__xor2_1_0/X a_11583_15239# -0
C447 CLA_1/sky130_fd_sc_hd__or4_1_0/B a_10923_15189# -0
C448 sky130_fd_sc_hd__mux4_1_0/a_1290_413# VDPWR 0.00165f
C449 a_2676_1791# sky130_fd_sc_hd__inv_1_0/Y 0
C450 a_6335_2153# sky130_fd_sc_hd__inv_1_0/A 0
C451 a_8431_5415# a_7285_5493# 0
C452 VDPWR CLA_0/a_145_n3151# 0.00275f
C453 VDPWR a_6429_5409# 0.01299f
C454 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__inv_1_0/A 0.76181f
C455 sky130_fd_sc_hd__mux2_1_0/S a_14432_4997# 0
C456 a_12587_5459# a_14152_5917# 0
C457 a_13969_2159# VDPWR 0
C458 VDPWR a_9741_12567# 0.0685f
C459 sky130_fd_sc_hd__fa_1_8/SUM a_3199_5501# 0
C460 VDPWR a_11409_5047# 0.10372f
C461 a_16275_5473# VDPWR 0
C462 a_11145_2243# sky130_fd_sc_hd__fa_1_5/SUM 0
C463 sky130_fd_sc_hd__inv_1_7/A sky130_fd_sc_hd__inv_1_5/A 0
C464 a_10121_1793# sky130_fd_sc_hd__fa_1_4/CIN 0
C465 a_15681_4997# a_15401_5917# 0
C466 a_14432_4997# a_14152_5917# 0
C467 a_9619_16343# CLA_1/sky130_fd_sc_hd__xor2_1_0/X 0
C468 sky130_fd_sc_hd__inv_1_1/A a_17544_4895# 0
C469 a_13443_5909# a_13679_5003# 0
C470 VDPWR CLA_0/a_n55_n517# 0.1235f
C471 a_15522_4547# sky130_fd_sc_hd__inv_1_0/A 0
C472 a_12978_1793# VDPWR 0
C473 a_6036_5493# a_7285_5493# -0.00146f
C474 a_12587_5459# sky130_fd_sc_hd__fa_1_16/CIN 0
C475 VDPWR a_16847_4529# 0.01685f
C476 VDPWR a_9461_14779# 0.00528f
C477 VDPWR a_2175_5051# 0
C478 VDPWR a_10261_5471# 0
C479 a_12194_5909# a_12419_5459# -0
C480 CLA_0/sky130_fd_sc_hd__and2_1_5/a_145_75# VDPWR 0.00202f
C481 a_9034_1793# sky130_fd_sc_hd__inv_1_0/A 0
C482 ui_in[0] sky130_fd_sc_hd__inv_1_1/A 0.08382f
C483 sky130_fd_sc_hd__inv_1_1/A a_13679_5003# 0
C484 sky130_fd_sc_hd__inv_1_1/A a_13520_4919# 0
C485 a_9287_5499# a_10160_5047# 0
C486 sky130_fd_sc_hd__fa_1_19/CIN a_17395_5923# 0
C487 a_10025_1793# sky130_fd_sc_hd__inv_1_0/A 0
C488 a_11250_4597# VDPWR 0
C489 sky130_fd_sc_hd__mux2_1_0/a_535_374# sky130_fd_sc_hd__mux2_1_0/A1 0.00143f
C490 CLA_1/sky130_fd_sc_hd__and4_1_0/B a_9871_14979# -0
C491 sky130_fd_sc_hd__fa_1_3/SUM sky130_fd_sc_hd__inv_1_0/A 0.00121f
C492 sky130_fd_sc_hd__fa_1_14/SUM a_14152_5917# -0
C493 VDPWR CLA_0/sky130_fd_sc_hd__or4_1_0/a_277_297# 0
C494 VDPWR a_10923_15189# 0.04038f
C495 VDPWR a_2706_5417# 0.00641f
C496 VDPWR a_12697_14007# 0
C497 a_4477_5043# sky130_fd_sc_hd__fa_1_8/CIN 0.00339f
C498 a_12823_4553# sky130_fd_sc_hd__inv_1_0/A 0
C499 a_12281_2159# a_13137_2243# -0
C500 CLA_0/sky130_fd_sc_hd__or4_1_0/X CLA_1/sky130_fd_sc_hd__and4_1_1/C 0.05432f
C501 sky130_fd_sc_hd__fa_1_6/CIN a_14065_1793# 0
C502 a_10132_5921# a_10357_5837# -0
C503 a_11409_5047# sky130_fd_sc_hd__fa_1_16/SUM 0
C504 VDPWR a_5239_2237# 0.0789f
C505 CLA_1/sky130_fd_sc_hd__or4_1_0/B CLA_1/sky130_fd_sc_hd__or2_1_0/A -0
C506 a_16847_4895# sky130_fd_sc_hd__mux2_1_0/A1 0
C507 a_10132_5921# sky130_fd_sc_hd__fa_1_17/SUM 0
C508 a_11225_14223# VDPWR 0.06629f
C509 VDPWR a_8431_5049# 0.01653f
C510 sky130_fd_sc_hd__fa_1_15/CIN a_16146_5923# 0.06783f
C511 sky130_fd_sc_hd__inv_1_9/Y sky130_fd_sc_hd__inv_1_11/A 0.05599f
C512 CLA_0/sky130_fd_sc_hd__or2_1_0/a_150_297# VDPWR 0
C513 VDPWR CLA_0/a_n63_n2185# 0.12486f
C514 sky130_fd_sc_hd__inv_1_2/Y CLA_0/sky130_fd_sc_hd__or4_1_0/X 0.05689f
C515 a_16902_5839# a_15401_5917# 0
C516 VDPWR a_14908_5833# 0.00836f
C517 sky130_fd_sc_hd__fa_1_12/COUT sky130_fd_sc_hd__mux2_1_0/S 0.00435f
C518 a_16129_1793# VDPWR 0
C519 sky130_fd_sc_hd__fa_1_18/SUM sky130_fd_sc_hd__fa_1_14/CIN 0
C520 sky130_fd_sc_hd__fa_1_1/SUM VDPWR 0.0791f
C521 VDPWR a_10289_4963# 0
C522 sky130_fd_sc_hd__mux2_1_0/A1 sky130_fd_sc_hd__mux2_1_0/a_439_47# 0
C523 VDPWR a_12281_2159# 0.01291f
C524 sky130_fd_sc_hd__inv_1_0/A a_16297_2159# 0.00107f
C525 a_2706_5051# sky130_fd_sc_hd__fa_1_8/CIN 0
C526 VDPWR a_17395_5923# 0.0929f
C527 VDPWR CLA_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 0.06629f
C528 a_11381_5921# a_10160_5047# 0
C529 a_12978_2159# VDPWR 0
C530 sky130_fd_sc_hd__fa_1_12/COUT a_14152_5917# 0
C531 VDPWR a_9621_12861# 0.00385f
C532 ui_in[1] sky130_fd_sc_hd__mux4_1_0/a_27_47# 0
C533 sky130_fd_sc_hd__inv_1_1/A a_13443_5909# 0.00752f
C534 sky130_fd_sc_hd__inv_1_2/Y CLA_0/sky130_fd_sc_hd__xor2_1_0/X 0.22566f
C535 ui_in[0] sky130_fd_sc_hd__mux4_1_0/a_27_413# 0.00288f
C536 a_9287_5499# sky130_fd_sc_hd__fa_1_11/SUM -0
C537 sky130_fd_sc_hd__inv_1_1/Y a_4213_5409# 0
C538 a_16902_5473# sky130_fd_sc_hd__fa_1_15/CIN -0
C539 a_14908_5833# sky130_fd_sc_hd__fa_1_18/CIN 0
C540 sky130_fd_sc_hd__fa_1_9/CIN sky130_fd_sc_hd__fa_1_8/CIN 0
C541 ua[0] sky130_fd_sc_hd__inv_1_0/A 0
C542 CLA_1/sky130_fd_sc_hd__or2_1_0/B VDPWR 0.12266f
C543 a_12323_5825# sky130_fd_sc_hd__inv_1_1/A 0
C544 VDPWR CLA_1/sky130_fd_sc_hd__or2_1_0/A 0.14947f
C545 a_12644_1793# sky130_fd_sc_hd__fa_1_6/CIN 0
C546 uio_out[6] uio_out[5] 0.03102f
C547 sky130_fd_sc_hd__fa_1_7/SUM a_15089_2243# 0
C548 sky130_fd_sc_hd__fa_1_9/COUT a_8167_5049# 0
C549 sky130_fd_sc_hd__fa_1_6/SUM a_13137_2243# 0
C550 a_16371_5839# sky130_fd_sc_hd__inv_1_1/A 0
C551 a_14377_5467# sky130_fd_sc_hd__fa_1_14/CIN 0
C552 a_12194_5909# a_11381_5921# 0.00291f
C553 CLA_0/sky130_fd_sc_hd__and4_1_0/B CLA_0/a_n55_n517# -0
C554 a_14825_4913# a_16454_4979# 0
C555 a_13679_5003# a_13186_4919# 0
C556 sky130_fd_sc_hd__mux4_1_0/a_750_97# VDPWR 0.00307f
C557 sky130_fd_sc_hd__fa_1_3/CIN sky130_fd_sc_hd__fa_1_3/SUM 0.05168f
C558 VDPWR sky130_fd_sc_hd__fa_1_15/SUM 0.08255f
C559 CLA_0/sky130_fd_sc_hd__and2_1_5/a_145_75# CLA_0/sky130_fd_sc_hd__and4_1_0/B -0
C560 sky130_fd_sc_hd__inv_1_1/A a_15522_4913# 0
C561 VDPWR sky130_fd_sc_hd__fa_1_9/SUM 0.07934f
C562 CLA_1/sky130_fd_sc_hd__and4_1_0/B a_9739_15799# -0
C563 ui_in[0] ua[0] 0.38436f
C564 VDPWR a_16583_4895# 0
C565 VDPWR a_12281_1793# 0.01618f
C566 a_3040_5051# VDPWR 0
C567 sky130_fd_sc_hd__mux2_1_0/S a_15681_4997# 0
C568 a_16679_4529# sky130_fd_sc_hd__fa_1_19/CIN 0
C569 sky130_fd_sc_hd__fa_1_6/SUM VDPWR 0.07933f
C570 a_15089_2243# a_14596_2159# 0
C571 a_12587_5459# VDPWR 0.01823f
C572 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__inv_1_2/A -0
C573 CLA_1/sky130_fd_sc_hd__and4_1_0/B VDPWR 0.81349f
C574 sky130_fd_sc_hd__mux2_1_0/S a_17703_4979# 0
C575 VDPWR sky130_fd_sc_hd__mux4_1_0/a_193_413# 0.01659f
C576 CLA_1/sky130_fd_sc_hd__and4_1_0/B a_9577_15377# -0
C577 a_6261_5043# sky130_fd_sc_hd__inv_1_1/A 0
C578 sky130_fd_sc_hd__fa_1_0/SUM sky130_fd_sc_hd__inv_1_0/Y 0.0073f
C579 ua[7] VDPWR 0
C580 a_6792_5043# a_8038_5499# 0
C581 VDPWR a_14432_4997# 0.05148f
C582 CLA_1/sky130_fd_sc_hd__or2_1_0/B a_11949_13849# -0
C583 sky130_fd_sc_hd__mux4_1_0/a_757_363# VDPWR 0.00545f
C584 a_11949_13849# CLA_1/sky130_fd_sc_hd__or2_1_0/A 0
C585 a_15188_4913# a_16454_4979# 0
C586 a_14545_5833# sky130_fd_sc_hd__fa_1_14/CIN 0
C587 CLA_0/sky130_fd_sc_hd__or4_1_0/X a_12009_15689# 0.00853f
C588 sky130_fd_sc_hd__inv_1_1/A a_10525_5837# 0.0014f
C589 uio_in[3] uio_in[2] 0.03102f
C590 a_9193_2243# sky130_fd_sc_hd__inv_1_0/A 0.00304f
C591 VDPWR a_6261_5409# 0.00109f
C592 sky130_fd_sc_hd__fa_1_12/CIN sky130_fd_sc_hd__fa_1_14/CIN 0
C593 a_12430_5003# sky130_fd_sc_hd__inv_1_0/A 0
C594 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__mux4_1_0/a_27_413# 0.00138f
C595 a_11165_13381# a_9863_13311# -0
C596 VDPWR a_13284_5459# 0
C597 VDPWR a_9128_5049# 0
C598 sky130_fd_sc_hd__inv_1_5/A sky130_fd_sc_hd__inv_1_4/A 0.05599f
C599 a_8038_5499# VDPWR 0.04423f
C600 a_17236_5839# VDPWR 0
C601 a_13840_2243# sky130_fd_sc_hd__inv_1_0/A 0.00211f
C602 VDPWR sky130_fd_sc_hd__fa_1_14/SUM 0.08715f
C603 ui_in[1] sky130_fd_sc_hd__mux4_1_0/a_247_21# -0
C604 a_7285_5493# sky130_fd_sc_hd__fa_1_9/CIN 0.00156f
C605 sky130_fd_sc_hd__mux2_1_0/S a_10132_5921# 0
C606 a_16539_5839# a_15401_5917# 0
C607 a_17395_5923# sky130_fd_sc_hd__mux2_1_0/A0 0.00883f
C608 a_15188_4547# sky130_fd_sc_hd__inv_1_0/A 0
C609 a_3990_2237# a_4383_2153# 0.01182f
C610 a_9896_2243# sky130_fd_sc_hd__inv_1_0/A 0.00211f
C611 a_12823_4919# a_14432_4997# 0
C612 uio_out[6] uio_out[7] 0.03102f
C613 VDPWR CLA_0/a_69_n4715# 0.07651f
C614 CLA_0/sky130_fd_sc_hd__and4_1_0/a_27_47# CLA_0/sky130_fd_sc_hd__and4_1_0/B -0
C615 a_14432_4997# sky130_fd_sc_hd__fa_1_18/CIN 0.06767f
C616 VDPWR a_16679_4529# 0
C617 CLA_1/sky130_fd_sc_hd__and4_1_0/B a_10761_14767# -0
C618 a_9619_16093# VDPWR 0.0037f
C619 VDPWR a_9629_14779# 0.02537f
C620 uio_in[6] uio_in[7] 0.03102f
C621 a_11145_2243# sky130_fd_sc_hd__fa_1_4/SUM -0
C622 VDPWR a_11222_5837# 0
C623 a_10289_2159# sky130_fd_sc_hd__inv_1_0/A 0
C624 sky130_fd_sc_hd__inv_1_2/Y CLA_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 0
C625 sky130_fd_sc_hd__inv_1_9/Y sky130_fd_sc_hd__inv_1_9/A 0.05423f
C626 a_5174_5043# sky130_fd_sc_hd__inv_1_1/Y 0
C627 sky130_fd_sc_hd__inv_1_1/A a_13186_4919# 0
C628 a_15904_2243# a_15089_2243# 0.00358f
C629 a_13679_5003# a_12430_5003# -0.00146f
C630 VDPWR a_8169_1793# 0
C631 a_10986_2159# sky130_fd_sc_hd__inv_1_0/A 0
C632 VDPWR a_9629_14529# 0.0042f
C633 a_11225_14223# a_10799_13773# 0
C634 sky130_fd_sc_hd__fa_1_12/CIN a_12194_5909# 0.06768f
C635 a_9873_11747# a_9741_12567# 0
C636 a_7032_2153# VDPWR 0
C637 a_15188_4547# a_13679_5003# 0
C638 a_3990_2237# a_3169_2241# 0.00332f
C639 a_4309_5043# sky130_fd_sc_hd__fa_1_8/CIN 0
C640 a_12655_4553# sky130_fd_sc_hd__inv_1_0/A 0
C641 a_6071_2153# sky130_fd_sc_hd__inv_1_0/Y 0
C642 a_16371_5473# a_16146_5923# -0
C643 a_12950_5459# a_14152_5917# 0
C644 sky130_fd_sc_hd__fa_1_2/CIN a_7191_2237# 0.00156f
C645 a_16679_4895# sky130_fd_sc_hd__mux2_1_0/A1 0
C646 a_11381_5921# a_11409_5047# 0.00177f
C647 sky130_fd_sc_hd__fa_1_12/COUT VDPWR 0.09487f
C648 a_4383_2153# sky130_fd_sc_hd__inv_1_0/Y 0
C649 sky130_fd_sc_hd__fa_1_17/SUM sky130_fd_sc_hd__inv_1_0/A 0
C650 VDPWR CLA_0/sky130_fd_sc_hd__and2_1_4/a_59_75# 0.0463f
C651 a_6335_1787# sky130_fd_sc_hd__fa_1_2/CIN 0.00339f
C652 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__inv_1_1/Y 0.07047f
C653 VDPWR a_8167_5415# 0
C654 a_12950_5459# sky130_fd_sc_hd__fa_1_16/CIN 0
C655 VDPWR a_1920_2241# 0.06177f
C656 a_15681_4997# sky130_fd_sc_hd__fa_1_19/CIN 0.00786f
C657 VDPWR a_4746_1787# 0.02482f
C658 VDPWR a_12113_2159# 0.00103f
C659 sky130_fd_sc_hd__inv_1_0/A a_16129_2159# 0
C660 sky130_fd_sc_hd__fa_1_16/CIN a_12559_4553# 0
C661 a_9193_2243# sky130_fd_sc_hd__fa_1_3/CIN 0.00155f
C662 sky130_fd_sc_hd__fa_1_9/COUT sky130_fd_sc_hd__inv_1_1/A 0.00284f
C663 a_12644_2159# VDPWR 0.00623f
C664 VDPWR sky130_fd_sc_hd__mux2_1_0/a_218_47# 0
C665 sky130_fd_sc_hd__fa_1_19/CIN a_17703_4979# 0.00156f
C666 VDPWR a_9621_13111# 0.02399f
C667 a_10525_5471# a_11409_5047# 0
C668 uio_oe[7] uio_oe[6] 0.03102f
C669 a_4213_5043# sky130_fd_sc_hd__inv_1_1/Y 0
C670 a_3169_2241# sky130_fd_sc_hd__inv_1_0/Y 0.04725f
C671 VDPWR a_12950_5825# 0.00837f
C672 a_13443_5909# a_12430_5003# 0
C673 uio_oe[0] uio_out[7] 0.03102f
C674 a_14825_4913# sky130_fd_sc_hd__inv_1_1/A 0
C675 VDPWR sky130_fd_sc_hd__fa_1_8/CIN 0.57283f
C676 a_8431_5415# sky130_fd_sc_hd__inv_1_1/A 0
C677 a_16539_5473# sky130_fd_sc_hd__fa_1_15/CIN 0.0034f
C678 sky130_fd_sc_hd__fa_1_7/CIN sky130_fd_sc_hd__inv_1_0/A 0.00765f
C679 sky130_fd_sc_hd__inv_1_1/A a_12430_5003# 0
C680 a_13029_14207# CLA_1/sky130_fd_sc_hd__xor2_1_0/X -0
C681 sky130_fd_sc_hd__inv_1_0/A a_5942_2237# 0
C682 CLA_0/sky130_fd_sc_hd__or4_1_0/a_27_297# CLA_0/sky130_fd_sc_hd__or4_1_0/A -0.00166f
C683 VDPWR CLA_0/a_195_n517# 0.02537f
C684 ua[5] a_10986_1793# 0
C685 a_12419_5825# sky130_fd_sc_hd__inv_1_1/A 0
C686 sky130_fd_sc_hd__fa_1_5/CIN a_13137_2243# 0.00156f
C687 a_7944_2243# a_7191_2237# 0.0035f
C688 a_11145_2243# a_11888_2243# 0.00395f
C689 VDPWR a_17236_5473# 0
C690 CLA_0/sky130_fd_sc_hd__or4_1_0/X a_10923_15189# -0
C691 a_16275_5839# sky130_fd_sc_hd__inv_1_1/A 0
C692 sky130_fd_sc_hd__fa_1_6/SUM sky130_fd_sc_hd__fa_1_6/CIN 0.05218f
C693 sky130_fd_sc_hd__mux2_1_0/a_76_199# a_17703_4979# 0
C694 a_6036_5493# sky130_fd_sc_hd__inv_1_1/A 0
C695 VDPWR a_3010_1791# 0
C696 VDPWR a_15681_4997# 0.09897f
C697 a_9741_12567# a_9751_11003# -0
C698 CLA_1/sky130_fd_sc_hd__and4_1_0/B a_10799_13773# 0
C699 a_10986_1793# sky130_fd_sc_hd__inv_1_0/A 0
C700 a_16902_5839# sky130_fd_sc_hd__fa_1_19/CIN 0
C701 a_7944_2243# a_6335_1787# 0
C702 sky130_fd_sc_hd__inv_1_1/A a_15188_4913# 0
C703 a_14657_4547# sky130_fd_sc_hd__inv_1_0/A 0
C704 a_8337_1793# sky130_fd_sc_hd__inv_1_0/A 0
C705 CLA_0/sky130_fd_sc_hd__or2_1_0/B VDPWR 0.12266f
C706 VDPWR CLA_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# 0.00472f
C707 VDPWR a_12113_1793# 0
C708 VDPWR a_17703_4979# 0.09056f
C709 a_14281_5467# sky130_fd_sc_hd__fa_1_14/CIN 0
C710 CLA_0/sky130_fd_sc_hd__or2_1_0/a_150_297# CLA_0/sky130_fd_sc_hd__or4_1_0/C -0
C711 sky130_fd_sc_hd__fa_1_5/CIN VDPWR 0.55799f
C712 a_16583_4529# sky130_fd_sc_hd__fa_1_19/CIN 0
C713 a_9193_2243# sky130_fd_sc_hd__fa_1_3/SUM -0
C714 a_9587_13813# VDPWR 0.00293f
C715 sky130_fd_sc_hd__fa_1_12/CIN a_11409_5047# 0
C716 sky130_fd_sc_hd__fa_1_12/COUT a_14545_5467# 0
C717 sky130_fd_sc_hd__mux2_1_0/S a_16454_4979# 0
C718 VDPWR a_1950_5501# 0.06171f
C719 a_6429_5043# a_8038_5499# 0
C720 ua[6] VDPWR 0.00159f
C721 VDPWR a_2079_5417# 0
C722 CLA_0/sky130_fd_sc_hd__and4_1_0/a_27_47# CLA_0/sky130_fd_sc_hd__or4_1_0/C -0
C723 a_3990_2237# a_5239_2237# -0.00146f
C724 VDPWR a_9463_11547# 0.00557f
C725 a_15681_4997# sky130_fd_sc_hd__fa_1_18/CIN 0.00156f
C726 CLA_1/sky130_fd_sc_hd__xor2_1_0/X a_9871_14979# -0
C727 sky130_fd_sc_hd__inv_1_1/A a_10357_5837# 0
C728 VDPWR a_6165_5409# 0
C729 a_15401_5917# sky130_fd_sc_hd__inv_1_1/A 0.00768f
C730 VDPWR a_10132_5921# 0.10943f
C731 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__fa_1_17/SUM 0
C732 sky130_fd_sc_hd__fa_1_8/SUM sky130_fd_sc_hd__fa_1_8/CIN 0.05073f
C733 a_8038_5499# a_9287_5499# -0.00146f
C734 a_3169_2241# a_2676_1791# 0
C735 VDPWR a_7285_5493# 0.07952f
C736 a_16902_5839# VDPWR 0.00741f
C737 CLA_0/sky130_fd_sc_hd__or4_1_0/A CLA_0/sky130_fd_sc_hd__or2_1_0/A -0
C738 CLA_0/sky130_fd_sc_hd__or4_1_0/X CLA_1/sky130_fd_sc_hd__or2_1_0/A 0
C739 a_8337_2159# sky130_fd_sc_hd__inv_1_0/A 0
C740 a_14825_4547# sky130_fd_sc_hd__inv_1_0/A 0
C741 CLA_0/sky130_fd_sc_hd__and4_1_0/a_27_47# CLA_0/sky130_fd_sc_hd__xor2_1_0/X 0
C742 sky130_fd_sc_hd__fa_1_15/CIN sky130_fd_sc_hd__fa_1_14/CIN 0
C743 sky130_fd_sc_hd__mux2_1_0/a_218_47# sky130_fd_sc_hd__mux2_1_0/A0 0
C744 VDPWR a_9589_10581# 0.00188f
C745 VDPWR a_16583_4529# 0
C746 a_12587_5459# a_11381_5921# 0
C747 VDPWR a_10888_5837# 0.00955f
C748 a_10121_2159# sky130_fd_sc_hd__inv_1_0/A 0
C749 a_12950_5459# VDPWR 0.0281f
C750 a_16146_5923# a_17395_5923# -0.00146f
C751 a_4840_5043# sky130_fd_sc_hd__inv_1_1/Y 0
C752 a_8794_5049# a_10160_5047# 0
C753 sky130_fd_sc_hd__inv_1_0/Y a_5239_2237# 0.00305f
C754 ui_in[1] sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.02886f
C755 a_10652_2159# sky130_fd_sc_hd__inv_1_0/A 0
C756 VDPWR a_12559_4553# 0
C757 a_12559_4919# a_11409_5047# 0
C758 CLA_0/a_195_n517# CLA_0/sky130_fd_sc_hd__and4_1_0/B -0
C759 sky130_fd_sc_hd__fa_1_2/CIN a_5239_2237# 0.00764f
C760 sky130_fd_sc_hd__fa_1_5/CIN sky130_fd_sc_hd__fa_1_4/CIN 0
C761 VDPWR a_12323_5459# 0
C762 a_14825_4547# a_13679_5003# 0
C763 sky130_fd_sc_hd__mux2_1_0/A0 a_17236_5473# 0
C764 a_8263_5415# sky130_fd_sc_hd__inv_1_1/A 0
C765 sky130_fd_sc_hd__mux2_1_0/S a_13679_5003# 0
C766 sky130_fd_sc_hd__fa_1_16/CIN sky130_fd_sc_hd__inv_1_0/A 0.00102f
C767 CLA_1/sky130_fd_sc_hd__or4_1_0/B CLA_1/sky130_fd_sc_hd__xor2_1_0/X -0
C768 sky130_fd_sc_hd__fa_1_1/SUM sky130_fd_sc_hd__inv_1_0/Y 0.00121f
C769 sky130_fd_sc_hd__fa_1_3/CIN a_8337_1793# 0.0034f
C770 a_9741_12567# a_9749_14235# -0
C771 CLA_0/sky130_fd_sc_hd__or4_1_0/X CLA_1/sky130_fd_sc_hd__and4_1_0/B 0.00102f
C772 a_4084_5493# sky130_fd_sc_hd__inv_1_1/Y 0.0021f
C773 CLA_0/sky130_fd_sc_hd__or4_1_0/B CLA_0/sky130_fd_sc_hd__or4_1_0/A -0.00383f
C774 VDPWR CLA_0/sky130_fd_sc_hd__and2_1_4/a_145_75# 0.00122f
C775 a_17153_2243# sky130_fd_sc_hd__inv_1_0/A 0.02678f
C776 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__inv_1_0/A 0.00718f
C777 sky130_fd_sc_hd__mux2_1_0/A0 a_17703_4979# 0
C778 a_16146_5923# sky130_fd_sc_hd__fa_1_15/SUM 0
C779 a_16539_5839# sky130_fd_sc_hd__fa_1_19/CIN 0
C780 VDPWR a_12017_2159# 0
C781 VDPWR CLA_0/a_67_n1483# 0.06644f
C782 sky130_fd_sc_hd__inv_1_0/A a_16033_2159# 0
C783 sky130_fd_sc_hd__fa_1_9/COUT a_8431_5415# 0
C784 a_13679_5003# sky130_fd_sc_hd__fa_1_16/CIN 0.00157f
C785 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__mux4_1_0/a_247_21# -0.00452f
C786 CLA_1/sky130_fd_sc_hd__xor2_1_0/X a_9739_15799# -0
C787 a_13443_5909# sky130_fd_sc_hd__fa_1_12/SUM -0
C788 a_16454_4979# sky130_fd_sc_hd__fa_1_19/CIN 0.06766f
C789 a_6036_5493# sky130_fd_sc_hd__inv_1_1/Y 0
C790 a_7126_5043# sky130_fd_sc_hd__inv_1_1/A 0
C791 a_17210_4895# a_17395_5923# 0
C792 VDPWR a_6698_2153# 0.00627f
C793 VDPWR a_6698_1787# 0.02483f
C794 a_14657_4913# sky130_fd_sc_hd__inv_1_1/A 0
C795 ui_in[0] sky130_fd_sc_hd__mux4_1_0/a_834_97# 0.00243f
C796 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__fa_1_12/SUM 0.003f
C797 ui_in[1] sky130_fd_sc_hd__mux4_1_0/a_668_97# 0
C798 a_16371_5473# sky130_fd_sc_hd__fa_1_15/CIN 0
C799 a_11222_5471# VDPWR 0
C800 a_11671_15239# VDPWR 0.00158f
C801 CLA_1/sky130_fd_sc_hd__and4_1_1/C a_12009_15689# -0.00255f
C802 CLA_1/sky130_fd_sc_hd__xor2_1_0/X VDPWR 0.70015f
C803 VDPWR sky130_fd_sc_hd__inv_1_8/A 0.42409f
C804 a_8337_2159# sky130_fd_sc_hd__fa_1_3/CIN 0
C805 a_15681_4997# sky130_fd_sc_hd__fa_1_19/SUM 0
C806 uio_out[5] uio_out[4] 0.03102f
C807 sky130_fd_sc_hd__mux2_1_0/S a_13443_5909# 0
C808 a_11225_14223# a_9749_14235# -0
C809 sky130_fd_sc_hd__fa_1_5/CIN sky130_fd_sc_hd__fa_1_6/CIN 0
C810 a_17703_4979# sky130_fd_sc_hd__fa_1_19/SUM -0
C811 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__fa_1_9/CIN 0.00183f
C812 a_12587_5459# sky130_fd_sc_hd__fa_1_12/CIN 0.00339f
C813 a_10916_4597# sky130_fd_sc_hd__inv_1_0/A 0
C814 ui_in[1] sky130_fd_sc_hd__mux4_1_0/a_1290_413# 0.13587f
C815 a_9896_2243# a_9193_2243# 0.00419f
C816 sky130_fd_sc_hd__mux2_1_0/a_505_21# a_17703_4979# 0
C817 sky130_fd_sc_hd__fa_1_7/CIN a_16297_2159# 0
C818 sky130_fd_sc_hd__mux2_1_0/S sky130_fd_sc_hd__inv_1_1/A 0.01648f
C819 VDPWR CLA_0/sky130_fd_sc_hd__and4_1_0/a_109_47# 0.00164f
C820 uio_oe[2] uio_oe[3] 0.03102f
C821 sky130_fd_sc_hd__fa_1_19/CIN sky130_fd_sc_hd__inv_1_0/A 0.00101f
C822 a_17210_4529# a_17395_5923# 0
C823 CLA_1/sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__inv_1_2/A 0
C824 a_14152_5917# a_13443_5909# 0.00359f
C825 a_16539_5839# VDPWR 0.01438f
C826 sky130_fd_sc_hd__inv_1_8/A sky130_fd_sc_hd__inv_1_2/A 0
C827 uio_out[2] uio_out[1] 0.03102f
C828 VDPWR a_4213_5409# 0
C829 VDPWR a_14561_4547# 0
C830 a_14152_5917# sky130_fd_sc_hd__inv_1_1/A 0.0052f
C831 CLA_1/sky130_fd_sc_hd__and4_1_1/C a_11777_15239# 0
C832 VDPWR sky130_fd_sc_hd__inv_1_5/A 0.49457f
C833 uio_in[6] uio_in[5] 0.03102f
C834 VDPWR a_16454_4979# 0.05353f
C835 VDPWR a_10993_13773# 0.00144f
C836 VDPWR a_8167_5049# 0
C837 a_13137_2243# sky130_fd_sc_hd__inv_1_0/A 0.00304f
C838 a_13443_5909# sky130_fd_sc_hd__fa_1_16/CIN 0
C839 a_11117_12361# a_11165_13381# 0
C840 CLA_1/sky130_fd_sc_hd__xor2_1_0/X a_10761_14767# -0
C841 sky130_fd_sc_hd__fa_1_12/COUT a_14377_5467# 0
C842 a_4477_5409# sky130_fd_sc_hd__fa_1_8/CIN 0
C843 CLA_1/sky130_fd_sc_hd__xor2_1_0/X a_11949_13849# 0
C844 a_2676_2157# VDPWR 0.00976f
C845 CLA_1/sky130_fd_sc_hd__and4_1_0/B a_9861_16543# -0
C846 a_7126_5409# sky130_fd_sc_hd__inv_1_1/A 0
C847 ua[5] VDPWR 0.00173f
C848 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__fa_1_16/CIN 0
C849 a_11810_13649# CLA_1/sky130_fd_sc_hd__or4_1_0/C -0
C850 sky130_fd_sc_hd__inv_1_5/A sky130_fd_sc_hd__inv_1_2/A 0
C851 a_9287_5499# a_10132_5921# 0
C852 VDPWR a_9631_11547# 0.02437f
C853 a_13186_4553# VDPWR 0.02585f
C854 sky130_fd_sc_hd__inv_1_1/A a_10261_5837# 0
C855 sky130_fd_sc_hd__inv_1_0/A a_13969_1793# 0
C856 sky130_fd_sc_hd__fa_1_0/SUM a_3169_2241# -0
C857 CLA_1/sky130_fd_sc_hd__or4_1_0/A a_12009_15689# 0
C858 a_6261_5043# sky130_fd_sc_hd__fa_1_9/CIN 0
C859 a_16275_5473# sky130_fd_sc_hd__fa_1_15/CIN 0
C860 sky130_fd_sc_hd__fa_1_18/CIN a_14561_4547# 0
C861 sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__inv_1_1/A 0.00659f
C862 a_14930_1793# sky130_fd_sc_hd__inv_1_0/A 0
C863 sky130_fd_sc_hd__fa_1_18/SUM a_15681_4997# -0
C864 VDPWR sky130_fd_sc_hd__inv_1_0/A 0.87761f
C865 a_15401_5917# a_15188_4547# 0
C866 CLA_1/sky130_fd_sc_hd__or4_1_0/C CLA_1/sky130_fd_sc_hd__or4_1_0/A -0.0146f
C867 rst_n ui_in[0] 0.03102f
C868 a_8169_2159# sky130_fd_sc_hd__inv_1_0/A 0
C869 VDPWR a_17544_4895# 0
C870 a_15401_5917# a_15188_4913# 0
C871 a_10025_2159# sky130_fd_sc_hd__inv_1_0/A 0
C872 a_4477_5043# sky130_fd_sc_hd__inv_1_1/Y 0
C873 a_13186_4553# sky130_fd_sc_hd__fa_1_18/CIN 0
C874 VDPWR a_9863_13311# 0.12717f
C875 CLA_1/sky130_fd_sc_hd__and4_1_0/B a_9749_14235# 0
C876 sky130_fd_sc_hd__fa_1_12/COUT sky130_fd_sc_hd__fa_1_12/CIN 0
C877 a_14908_5467# sky130_fd_sc_hd__inv_1_1/A 0
C878 a_16033_1793# sky130_fd_sc_hd__inv_1_0/A 0
C879 ui_in[0] VDPWR 0.47798f
C880 sky130_fd_sc_hd__inv_1_1/Y a_4309_5409# 0
C881 VDPWR a_13679_5003# 0.08706f
C882 VDPWR a_6167_1787# 0
C883 VDPWR a_13520_4919# 0
C884 a_12823_4553# sky130_fd_sc_hd__fa_1_16/CIN 0.00339f
C885 sky130_fd_sc_hd__fa_1_18/CIN sky130_fd_sc_hd__inv_1_0/A 0
C886 CLA_0/sky130_fd_sc_hd__or2_1_0/B CLA_0/sky130_fd_sc_hd__or4_1_0/C -0.00108f
C887 a_10132_5921# a_11381_5921# -0.00146f
C888 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_0/a_247_21# -0
C889 a_4084_5493# a_4477_5043# 0
C890 CLA_0/a_27_n517# VDPWR 0.00528f
C891 a_1920_2241# sky130_fd_sc_hd__inv_1_0/Y 0.03136f
C892 VDPWR a_8700_1793# 0.02483f
C893 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__fa_1_16/SUM 0
C894 ui_in[0] sky130_fd_sc_hd__inv_1_2/A 0.00242f
C895 sky130_fd_sc_hd__inv_1_0/Y a_4746_1787# 0
C896 CLA_1/sky130_fd_sc_hd__and4_1_1/C a_10923_15189# -0
C897 CLA_0/sky130_fd_sc_hd__and4_1_0/a_109_47# CLA_0/sky130_fd_sc_hd__and4_1_0/B -0
C898 VDPWR sky130_fd_sc_hd__fa_1_2/SUM 0.07926f
C899 sky130_fd_sc_hd__mux2_1_0/A1 a_17703_4979# 0.01326f
C900 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__fa_1_19/CIN 0
C901 a_4746_1787# sky130_fd_sc_hd__fa_1_2/CIN 0
C902 a_2706_5051# sky130_fd_sc_hd__inv_1_1/Y 0
C903 a_12587_5825# a_13679_5003# 0
C904 VDPWR a_5174_5043# 0
C905 a_12823_4919# a_13679_5003# -0
C906 sky130_fd_sc_hd__fa_1_18/CIN a_13679_5003# 0.00766f
C907 a_8700_2159# a_7191_2237# 0
C908 a_4840_5043# sky130_fd_sc_hd__fa_1_9/CIN 0
C909 sky130_fd_sc_hd__fa_1_15/CIN a_17395_5923# 0.00155f
C910 a_12950_5459# a_11381_5921# 0
C911 sky130_fd_sc_hd__fa_1_4/CIN sky130_fd_sc_hd__inv_1_0/A 0.00282f
C912 CLA_0/sky130_fd_sc_hd__and3_1_0/a_27_47# VDPWR 0.05475f
C913 CLA_1/sky130_fd_sc_hd__and4_1_1/C a_11225_14223# -0
C914 a_11777_15239# a_12009_15689# -0
C915 VDPWR a_4119_2153# 0
C916 a_10132_5921# sky130_fd_sc_hd__fa_1_13/SUM 0
C917 a_10887_13773# CLA_1/sky130_fd_sc_hd__or2_1_0/A 0
C918 sky130_fd_sc_hd__fa_1_9/CIN sky130_fd_sc_hd__inv_1_1/Y 0.0013f
C919 sky130_fd_sc_hd__inv_1_1/A a_8263_5049# 0
C920 a_13679_5003# sky130_fd_sc_hd__fa_1_16/SUM -0
C921 ui_in[1] sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.01723f
C922 a_10160_5047# a_11409_5047# -0.00146f
C923 a_6792_5043# sky130_fd_sc_hd__inv_1_1/A 0
C924 VDPWR sky130_fd_sc_hd__fa_1_3/CIN 0.55832f
C925 a_14561_4913# sky130_fd_sc_hd__inv_1_1/A 0
C926 sky130_fd_sc_hd__mux2_1_0/a_76_199# sky130_fd_sc_hd__inv_1_1/A 0.02374f
C927 sky130_fd_sc_hd__inv_1_0/Y a_3010_1791# 0
C928 sky130_fd_sc_hd__fa_1_9/COUT sky130_fd_sc_hd__fa_1_9/CIN 0
C929 VDPWR a_13443_5909# 0.10069f
C930 sky130_fd_sc_hd__fa_1_9/COUT sky130_fd_sc_hd__mux2_1_0/S 0
C931 VDPWR a_6335_2153# 0.01299f
C932 sky130_fd_sc_hd__fa_1_5/CIN a_11145_2243# 0.00764f
C933 VDPWR sky130_fd_sc_hd__inv_1_1/A 2.79348f
C934 ui_in[1] sky130_fd_sc_hd__mux4_1_0/a_757_363# -0
C935 VDPWR a_12323_5825# 0
C936 a_10553_4597# sky130_fd_sc_hd__inv_1_0/A 0
C937 sky130_fd_sc_hd__fa_1_15/CIN sky130_fd_sc_hd__fa_1_15/SUM 0.05191f
C938 sky130_fd_sc_hd__fa_1_4/CIN a_8700_1793# 0
C939 a_13284_5825# sky130_fd_sc_hd__inv_1_1/A 0
C940 sky130_fd_sc_hd__fa_1_5/CIN a_10652_1793# 0
C941 a_8337_2159# a_9193_2243# -0
C942 VDPWR CLA_0/sky130_fd_sc_hd__and4_1_0/a_197_47# 0.00152f
C943 sky130_fd_sc_hd__mux2_1_0/S a_12430_5003# 0
C944 CLA_1/sky130_fd_sc_hd__and4_1_1/C CLA_1/sky130_fd_sc_hd__or2_1_0/B 0
C945 a_16371_5839# VDPWR 0.00114f
C946 CLA_1/sky130_fd_sc_hd__and4_1_1/C CLA_1/sky130_fd_sc_hd__or2_1_0/A -0.00389f
C947 CLA_1/sky130_fd_sc_hd__or4_1_0/A a_12697_14007# 0
C948 a_5174_5409# sky130_fd_sc_hd__inv_1_1/Y 0
C949 VDPWR a_15522_4547# 0
C950 a_12587_5825# a_13443_5909# 0
C951 VDPWR a_4213_5043# 0
C952 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__inv_1_2/A 0.00503f
C953 a_6036_5493# sky130_fd_sc_hd__fa_1_9/CIN 0.0677f
C954 VDPWR a_15522_4913# 0
C955 a_9034_1793# VDPWR 0
C956 a_9749_14235# a_9621_13111# -0
C957 a_11225_14223# CLA_1/sky130_fd_sc_hd__or4_1_0/A -0
C958 a_12823_4919# sky130_fd_sc_hd__inv_1_1/A 0
C959 a_10160_5047# a_8431_5049# 0
C960 a_12587_5825# sky130_fd_sc_hd__inv_1_1/A 0.00113f
C961 a_17210_4895# a_17703_4979# 0
C962 sky130_fd_sc_hd__fa_1_18/CIN sky130_fd_sc_hd__inv_1_1/A 0
C963 VDPWR CLA_0/a_195_n767# 0.00409f
C964 sky130_fd_sc_hd__fa_1_6/CIN sky130_fd_sc_hd__inv_1_0/A 0.00282f
C965 VDPWR a_10025_1793# 0
C966 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__fa_1_19/SUM 0
C967 VDPWR sky130_fd_sc_hd__fa_1_3/SUM 0.07924f
C968 uio_oe[6] uio_oe[5] 0.03102f
C969 CLA_0/sky130_fd_sc_hd__or4_1_0/A VDPWR 0.5643f
C970 ua[4] a_14930_1793# 0
C971 a_6792_5409# sky130_fd_sc_hd__inv_1_1/A 0
C972 VDPWR a_4215_2153# 0.00102f
C973 ua[4] VDPWR 0.00174f
C974 a_12430_5003# sky130_fd_sc_hd__fa_1_16/CIN 0.06782f
C975 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__fa_1_16/SUM 0
C976 VDPWR sky130_fd_sc_hd__inv_1_7/A 0.3874f
C977 VDPWR a_2313_2157# 0.00915f
C978 a_12823_4553# VDPWR 0.01713f
C979 VDPWR a_9631_11297# 0.00333f
C980 sky130_fd_sc_hd__fa_1_4/CIN sky130_fd_sc_hd__fa_1_3/CIN 0
C981 sky130_fd_sc_hd__inv_1_0/A a_14930_2159# 0
C982 sky130_fd_sc_hd__inv_1_1/A a_9128_5415# 0
C983 a_6261_5043# VDPWR 0
C984 CLA_1/sky130_fd_sc_hd__and4_1_0/B CLA_1/sky130_fd_sc_hd__and4_1_1/C -0
C985 a_15681_4997# a_17210_4529# 0
C986 sky130_fd_sc_hd__fa_1_12/COUT a_14281_5467# 0
C987 a_6165_5043# sky130_fd_sc_hd__fa_1_9/CIN 0
C988 VDPWR a_10525_5837# 0.01832f
C989 VDPWR a_11583_15239# 0.00102f
C990 sky130_fd_sc_hd__fa_1_6/SUM a_15089_2243# -0
C991 VDPWR CLA_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0.0196f
C992 VDPWR sky130_fd_sc_hd__mux4_1_0/a_27_413# 0.04364f
C993 CLA_0/sky130_fd_sc_hd__or4_1_0/X CLA_1/sky130_fd_sc_hd__xor2_1_0/X 0.31578f
C994 sky130_fd_sc_hd__fa_1_1/CIN a_4383_1787# 0.00428f
C995 a_4383_2153# a_5239_2237# 0.00204f
C996 sky130_fd_sc_hd__inv_1_7/A sky130_fd_sc_hd__inv_1_2/A 0
C997 sky130_fd_sc_hd__mux2_1_0/S a_15401_5917# 0
C998 a_8073_2159# sky130_fd_sc_hd__inv_1_0/A 0
C999 a_12323_5459# sky130_fd_sc_hd__fa_1_12/CIN 0
C1000 CLA_1/sky130_fd_sc_hd__or4_1_0/A CLA_1/sky130_fd_sc_hd__or2_1_0/A -0
C1001 a_10888_5471# sky130_fd_sc_hd__inv_1_1/A 0
C1002 sky130_fd_sc_hd__inv_1_0/A a_13520_4553# 0
C1003 VDPWR a_16297_2159# 0.01294f
C1004 CLA_1/sky130_fd_sc_hd__or4_1_0/C a_12697_14007# -0
C1005 a_9619_16343# VDPWR 0.0204f
C1006 a_4309_5043# sky130_fd_sc_hd__inv_1_1/Y 0
C1007 a_15401_5917# a_14152_5917# -0.00146f
C1008 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__inv_1_2/A 0.00483f
C1009 a_14545_5467# sky130_fd_sc_hd__inv_1_1/A 0
C1010 a_16994_2159# sky130_fd_sc_hd__inv_1_0/A 0
C1011 VDPWR a_13186_4919# 0.00714f
C1012 CLA_1/sky130_fd_sc_hd__or4_1_0/C a_11225_14223# -0
C1013 a_12655_4553# sky130_fd_sc_hd__fa_1_16/CIN 0
C1014 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__mux2_1_0/A0 0.00921f
C1015 VDPWR CLA_0/sky130_fd_sc_hd__and4_1_1/a_27_47# 0.06138f
C1016 a_17544_4529# sky130_fd_sc_hd__inv_1_0/A 0
C1017 a_5333_5493# sky130_fd_sc_hd__fa_1_9/SUM 0
C1018 VDPWR ua[0] 0.1976f
C1019 sky130_fd_sc_hd__fa_1_4/CIN a_10025_1793# 0
C1020 sky130_fd_sc_hd__fa_1_18/SUM sky130_fd_sc_hd__inv_1_0/A 0
C1021 VDPWR a_4746_2153# 0.00621f
C1022 a_9619_16343# sky130_fd_sc_hd__inv_1_2/A 0
C1023 ui_in[6] ui_in[5] 0.03102f
C1024 a_14432_4997# sky130_fd_sc_hd__fa_1_14/CIN 0.00135f
C1025 sky130_fd_sc_hd__fa_1_5/CIN sky130_fd_sc_hd__fa_1_5/SUM 0.05174f
C1026 CLA_1/sky130_fd_sc_hd__and4_1_0/B CLA_1/sky130_fd_sc_hd__or4_1_0/A 0
C1027 sky130_fd_sc_hd__mux2_1_0/A1 a_16454_4979# 0
C1028 sky130_fd_sc_hd__fa_1_1/SUM a_3169_2241# 0
C1029 a_2343_5051# sky130_fd_sc_hd__inv_1_1/Y 0.00447f
C1030 sky130_fd_sc_hd__inv_1_1/A a_12419_5459# 0
C1031 sky130_fd_sc_hd__fa_1_9/COUT a_8263_5049# 0
C1032 a_8794_5415# a_10132_5921# 0
C1033 VDPWR a_4840_5043# 0.02482f
C1034 a_9873_11747# a_9863_13311# -0
C1035 CLA_0/sky130_fd_sc_hd__or4_1_0/a_27_297# VDPWR 0.04614f
C1036 a_6792_5043# sky130_fd_sc_hd__fa_1_9/COUT 0
C1037 sky130_fd_sc_hd__fa_1_10/SUM sky130_fd_sc_hd__inv_1_1/Y 0.0073f
C1038 a_8794_5415# a_7285_5493# 0
C1039 VDPWR sky130_fd_sc_hd__inv_1_1/Y 1.02951f
C1040 a_15188_4547# sky130_fd_sc_hd__fa_1_19/CIN 0
C1041 sky130_fd_sc_hd__fa_1_18/SUM a_13679_5003# 0
C1042 a_16146_5923# a_16454_4979# 0
C1043 a_10357_5471# a_10132_5921# -0
C1044 sky130_fd_sc_hd__fa_1_14/SUM sky130_fd_sc_hd__fa_1_14/CIN 0.0459f
C1045 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__fa_1_19/SUM 0
C1046 CLA_1/sky130_fd_sc_hd__or4_1_0/C CLA_1/sky130_fd_sc_hd__or2_1_0/B -0.00108f
C1047 a_11165_13381# VDPWR 0.05474f
C1048 CLA_1/sky130_fd_sc_hd__or4_1_0/C CLA_1/sky130_fd_sc_hd__or2_1_0/A -0
C1049 a_6429_5043# sky130_fd_sc_hd__inv_1_1/A 0
C1050 sky130_fd_sc_hd__fa_1_9/COUT VDPWR 0.56429f
C1051 sky130_fd_sc_hd__mux2_1_0/a_505_21# sky130_fd_sc_hd__inv_1_1/A 0.00367f
C1052 a_13840_2243# a_13137_2243# 0.00419f
C1053 sky130_fd_sc_hd__mux2_1_0/A1 sky130_fd_sc_hd__inv_1_0/A 0
C1054 VDPWR a_4084_5493# 0.04455f
C1055 VDPWR a_14825_4913# 0.01519f
C1056 a_9287_5499# sky130_fd_sc_hd__inv_1_1/A 0.00302f
C1057 a_9863_13311# CLA_0/sky130_fd_sc_hd__or4_1_0/C 0
C1058 VDPWR a_8431_5415# 0.01321f
C1059 VDPWR CLA_0/a_155_n4715# 0.00186f
C1060 CLA_1/sky130_fd_sc_hd__and4_1_0/B a_12009_15689# -0
C1061 VDPWR a_9193_2243# 0.07855f
C1062 a_17153_2243# sky130_fd_sc_hd__fa_1_7/CIN 0.00156f
C1063 CLA_1/sky130_fd_sc_hd__xor2_1_0/X a_9861_16543# -0
C1064 CLA_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# CLA_0/sky130_fd_sc_hd__and4_1_0/B -0
C1065 sky130_fd_sc_hd__inv_1_8/A sky130_fd_sc_hd__inv_1_6/A 0
C1066 uio_out[4] uio_out[3] 0.03102f
C1067 VDPWR a_12430_5003# 0.05027f
C1068 sky130_fd_sc_hd__mux2_1_0/A1 a_17544_4895# 0
C1069 sky130_fd_sc_hd__fa_1_15/CIN a_15681_4997# 0
C1070 VDPWR a_12419_5825# 0.00114f
C1071 a_3040_5417# sky130_fd_sc_hd__inv_1_1/Y 0
C1072 a_10385_4597# sky130_fd_sc_hd__inv_1_0/A 0
C1073 ua[5] a_11145_2243# 0
C1074 VDPWR a_13840_2243# 0.04368f
C1075 a_14596_1793# sky130_fd_sc_hd__inv_1_0/A 0
C1076 sky130_fd_sc_hd__fa_1_15/CIN a_17703_4979# 0
C1077 a_6036_5493# VDPWR 0.04542f
C1078 a_16275_5839# VDPWR 0
C1079 VDPWR a_2145_2157# 0.00111f
C1080 a_9896_2243# VDPWR 0.04368f
C1081 VDPWR a_15188_4547# 0.0262f
C1082 sky130_fd_sc_hd__fa_1_12/COUT sky130_fd_sc_hd__fa_1_14/CIN 0.00633f
C1083 a_4840_5409# sky130_fd_sc_hd__inv_1_1/Y 0
C1084 a_2676_2157# sky130_fd_sc_hd__inv_1_0/Y 0.00222f
C1085 sky130_fd_sc_hd__fa_1_7/SUM sky130_fd_sc_hd__inv_1_0/A 0.00174f
C1086 uio_out[1] uio_out[0] 0.03102f
C1087 sky130_fd_sc_hd__inv_1_8/A sky130_fd_sc_hd__inv_1_9/A 0.05352f
C1088 a_14825_4913# sky130_fd_sc_hd__fa_1_18/CIN 0
C1089 VDPWR a_15188_4913# 0.00733f
C1090 a_6698_1787# a_7944_2243# 0
C1091 a_10289_2159# VDPWR 0.01301f
C1092 a_11145_2243# sky130_fd_sc_hd__inv_1_0/A 0.00304f
C1093 uio_in[5] uio_in[4] 0.03102f
C1094 a_13029_14207# a_12793_14007# -0
C1095 a_12655_4919# sky130_fd_sc_hd__inv_1_1/A 0
C1096 a_11225_14223# a_10923_15189# -0
C1097 sky130_fd_sc_hd__inv_1_5/A sky130_fd_sc_hd__inv_1_6/A 0.05704f
C1098 a_12823_4919# a_12430_5003# -0
C1099 CLA_0/sky130_fd_sc_hd__or2_1_0/A VDPWR 0.14946f
C1100 VDPWR a_10986_2159# 0
C1101 CLA_0/sky130_fd_sc_hd__and4_1_1/a_27_47# CLA_0/sky130_fd_sc_hd__and4_1_0/B -0
C1102 sky130_fd_sc_hd__fa_1_8/SUM sky130_fd_sc_hd__inv_1_1/Y 0.00121f
C1103 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__inv_1_0/A 0.07042f
C1104 a_2343_5417# sky130_fd_sc_hd__inv_1_1/Y 0.00637f
C1105 sky130_fd_sc_hd__fa_1_18/SUM sky130_fd_sc_hd__inv_1_1/A 0
C1106 VDPWR sky130_fd_sc_hd__inv_1_4/A 0.33922f
C1107 a_10652_1793# sky130_fd_sc_hd__inv_1_0/A 0
C1108 sky130_fd_sc_hd__mux2_1_0/S a_14152_5917# 0
C1109 sky130_fd_sc_hd__fa_1_2/CIN sky130_fd_sc_hd__inv_1_0/A 0.00234f
C1110 a_11381_5921# sky130_fd_sc_hd__inv_1_1/A 0.00739f
C1111 CLA_0/sky130_fd_sc_hd__and4_1_1/C CLA_0/sky130_fd_sc_hd__and4_1_1/a_27_47# -0.00255f
C1112 ui_in[0] sky130_fd_sc_hd__mux4_1_0/a_923_363# 0.00109f
C1113 CLA_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# VDPWR 0.11056f
C1114 a_6165_5043# VDPWR 0
C1115 a_12655_4553# VDPWR 0
C1116 sky130_fd_sc_hd__inv_1_0/A a_14596_2159# 0
C1117 VDPWR CLA_0/sky130_fd_sc_hd__and4_1_0/a_303_47# 0.00144f
C1118 VDPWR a_10955_11939# 0.00122f
C1119 a_16994_1793# sky130_fd_sc_hd__inv_1_0/A 0
C1120 a_10289_4597# sky130_fd_sc_hd__inv_1_0/A 0
C1121 a_16902_5839# sky130_fd_sc_hd__fa_1_15/CIN 0
C1122 VDPWR a_10357_5837# 0.00154f
C1123 a_2343_5417# a_4084_5493# 0
C1124 VDPWR a_15401_5917# 0.08959f
C1125 sky130_fd_sc_hd__fa_1_1/SUM a_5239_2237# -0
C1126 sky130_fd_sc_hd__mux2_1_0/S sky130_fd_sc_hd__fa_1_16/CIN 0.04098f
C1127 a_11117_12361# VDPWR 0.04632f
C1128 VDPWR CLA_0/sky130_fd_sc_hd__xor2_1_0/a_285_47# 0.00347f
C1129 VDPWR sky130_fd_sc_hd__fa_1_17/SUM 0.04118f
C1130 sky130_fd_sc_hd__fa_1_12/CIN a_13679_5003# 0
C1131 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__inv_1_2/A 0
C1132 a_8073_1793# sky130_fd_sc_hd__inv_1_0/A 0
C1133 sky130_fd_sc_hd__fa_1_4/CIN a_9193_2243# 0.00764f
C1134 a_5333_5493# sky130_fd_sc_hd__fa_1_8/CIN 0.00156f
C1135 VDPWR a_2079_5051# 0
C1136 CLA_0/sky130_fd_sc_hd__or4_1_0/B VDPWR 0.34609f
C1137 a_6167_1787# sky130_fd_sc_hd__fa_1_2/CIN 0
C1138 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__fa_1_13/SUM 0.00331f
C1139 VDPWR CLA_0/a_29_n3749# 0.00528f
C1140 a_10525_5471# sky130_fd_sc_hd__inv_1_1/A 0
C1141 VDPWR a_16129_2159# 0.00104f
C1142 a_15681_4997# sky130_fd_sc_hd__fa_1_14/CIN 0
C1143 a_14377_5467# sky130_fd_sc_hd__inv_1_1/A 0
C1144 a_9896_2243# sky130_fd_sc_hd__fa_1_4/CIN 0.0677f
C1145 a_16660_2159# sky130_fd_sc_hd__inv_1_0/A 0.00205f
C1146 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__mux2_1_0/A1 0.01989f
C1147 sky130_fd_sc_hd__fa_1_2/SUM sky130_fd_sc_hd__inv_1_0/Y 0.00121f
C1148 sky130_fd_sc_hd__fa_1_18/CIN a_15401_5917# 0.00129f
C1149 CLA_1/sky130_fd_sc_hd__or2_1_0/B a_11225_14223# -0
C1150 a_10289_2159# sky130_fd_sc_hd__fa_1_4/CIN 0
C1151 a_11225_14223# CLA_1/sky130_fd_sc_hd__or2_1_0/A 0
C1152 sky130_fd_sc_hd__fa_1_1/CIN a_4215_1787# 0
C1153 VDPWR CLA_0/sky130_fd_sc_hd__and4_1_1/a_109_47# 0.00102f
C1154 sky130_fd_sc_hd__fa_1_2/SUM sky130_fd_sc_hd__fa_1_2/CIN 0.05218f
C1155 sky130_fd_sc_hd__fa_1_7/CIN VDPWR 0.54328f
C1156 a_17210_4529# sky130_fd_sc_hd__inv_1_0/A 0
C1157 sky130_fd_sc_hd__fa_1_1/CIN VDPWR 0.5665f
C1158 a_15904_2243# sky130_fd_sc_hd__inv_1_0/A 0.00324f
C1159 a_14233_2159# sky130_fd_sc_hd__inv_1_0/A 0
C1160 VDPWR a_5942_2237# 0.04634f
C1161 a_7944_2243# sky130_fd_sc_hd__inv_1_0/A 0.00211f
C1162 a_16146_5923# sky130_fd_sc_hd__inv_1_1/A 0.00525f
C1163 a_13029_14207# a_12865_14007# -0
C1164 sky130_fd_sc_hd__inv_1_0/Y a_4119_2153# 0
C1165 VDPWR a_8263_5415# 0.00104f
C1166 a_2175_5417# sky130_fd_sc_hd__inv_1_1/Y 0
C1167 a_14545_5833# a_13443_5909# 0
C1168 a_3169_2241# a_1920_2241# -0.00146f
C1169 CLA_0/sky130_fd_sc_hd__or4_1_0/A CLA_0/sky130_fd_sc_hd__or4_1_0/C -0.0146f
C1170 CLA_0/sky130_fd_sc_hd__or4_1_0/X CLA_0/sky130_fd_sc_hd__or4_1_0/A 0.02609f
C1171 CLA_1/sky130_fd_sc_hd__and4_1_0/B a_10923_15189# -0.00106f
C1172 CLA_1/sky130_fd_sc_hd__or4_1_0/B a_13029_14207# -0
C1173 a_10986_1793# VDPWR 0
C1174 VDPWR a_4477_5043# 0.01626f
C1175 sky130_fd_sc_hd__fa_1_12/CIN a_13443_5909# 0.00156f
C1176 a_16371_5839# a_16146_5923# -0
C1177 sky130_fd_sc_hd__fa_1_7/CIN a_16033_1793# 0
C1178 a_14545_5833# sky130_fd_sc_hd__inv_1_1/A 0.00115f
C1179 a_3199_5501# sky130_fd_sc_hd__fa_1_8/CIN 0.00988f
C1180 VDPWR a_14657_4547# 0
C1181 CLA_1/sky130_fd_sc_hd__xor2_1_0/X a_10887_13773# -0
C1182 VDPWR a_4309_5409# 0.00104f
C1183 sky130_fd_sc_hd__fa_1_3/CIN sky130_fd_sc_hd__fa_1_2/CIN 0
C1184 a_10132_5921# a_10160_5047# 0
C1185 VDPWR a_5080_2153# 0
C1186 VDPWR a_8337_1793# 0.01619f
C1187 a_7032_1787# sky130_fd_sc_hd__inv_1_0/A 0
C1188 a_4383_1787# a_4215_1787# 0
C1189 sky130_fd_sc_hd__mux2_1_0/S sky130_fd_sc_hd__fa_1_19/CIN 0.03084f
C1190 sky130_fd_sc_hd__fa_1_12/CIN sky130_fd_sc_hd__inv_1_1/A 0.00685f
C1191 a_9749_14235# a_9863_13311# -0
C1192 CLA_1/sky130_fd_sc_hd__and4_1_0/B a_11225_14223# -0
C1193 a_4383_1787# VDPWR 0.01876f
C1194 a_17395_5923# sky130_fd_sc_hd__fa_1_15/SUM -0
C1195 a_9287_5499# sky130_fd_sc_hd__fa_1_9/COUT 0.00155f
C1196 VDPWR a_9453_13111# 0.00559f
C1197 CLA_0/sky130_fd_sc_hd__or4_1_0/A CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0
C1198 a_16902_5473# sky130_fd_sc_hd__inv_1_1/A 0
C1199 a_6335_2153# sky130_fd_sc_hd__fa_1_2/CIN 0
C1200 VDPWR a_6167_2153# 0.00119f
C1201 CLA_1/sky130_fd_sc_hd__or2_1_0/B CLA_1/sky130_fd_sc_hd__or2_1_0/A -0
C1202 CLA_0/sky130_fd_sc_hd__and4_1_1/C CLA_0/sky130_fd_sc_hd__or2_1_0/A -0.00389f
C1203 sky130_fd_sc_hd__fa_1_5/SUM sky130_fd_sc_hd__inv_1_0/A 0.00121f
C1204 sky130_fd_sc_hd__mux2_1_0/a_218_374# sky130_fd_sc_hd__inv_1_1/A 0.0023f
C1205 a_8073_1793# sky130_fd_sc_hd__fa_1_3/CIN 0
C1206 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__mux4_1_0/a_247_21# -0.00115f
C1207 CLA_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# CLA_0/sky130_fd_sc_hd__and4_1_0/B -0
C1208 ua[6] a_7191_2237# 0
C1209 a_13840_2243# sky130_fd_sc_hd__fa_1_6/CIN 0.0677f
C1210 a_7126_5043# VDPWR 0
C1211 a_9287_5499# a_8431_5415# 0
C1212 sky130_fd_sc_hd__fa_1_5/CIN a_12017_1793# 0
C1213 VDPWR a_14657_4913# 0.00113f
C1214 a_9619_16343# CLA_0/sky130_fd_sc_hd__or4_1_0/X 0
C1215 VDPWR a_2706_5051# 0.02496f
C1216 VDPWR sky130_fd_sc_hd__fa_1_12/SUM 0.08286f
C1217 sky130_fd_sc_hd__fa_1_18/CIN a_14657_4547# 0
C1218 a_10916_4597# sky130_fd_sc_hd__fa_1_16/CIN 0
C1219 sky130_fd_sc_hd__mux4_1_0/a_27_47# sky130_fd_sc_hd__inv_1_1/A 0.00542f
C1220 uo_out[6] uo_out[5] 0.03102f
C1221 a_17210_4895# sky130_fd_sc_hd__inv_1_1/A 0
C1222 CLA_0/sky130_fd_sc_hd__and3_1_0/a_109_47# VDPWR 0.00209f
C1223 a_13029_14207# VDPWR 0.03959f
C1224 a_16660_1793# sky130_fd_sc_hd__inv_1_0/A 0.00236f
C1225 a_16539_5839# sky130_fd_sc_hd__fa_1_15/CIN 0
C1226 CLA_1/sky130_fd_sc_hd__and4_1_1/C a_11671_15239# 0
C1227 CLA_1/sky130_fd_sc_hd__xor2_1_0/X CLA_1/sky130_fd_sc_hd__and4_1_1/C -0.00252f
C1228 VDPWR sky130_fd_sc_hd__fa_1_9/CIN 0.56509f
C1229 a_14233_1793# sky130_fd_sc_hd__inv_1_0/A 0
C1230 ui_in[0] sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.09466f
C1231 a_1950_5501# a_3199_5501# -0.00146f
C1232 VDPWR a_8337_2159# 0.01291f
C1233 VDPWR a_14825_4547# 0.01799f
C1234 sky130_fd_sc_hd__fa_1_15/CIN a_16454_4979# 0
C1235 VDPWR sky130_fd_sc_hd__mux2_1_0/S 4.25114f
C1236 CLA_1/sky130_fd_sc_hd__and4_1_0/B CLA_1/sky130_fd_sc_hd__or2_1_0/A -0
C1237 a_4477_5409# sky130_fd_sc_hd__inv_1_1/Y 0
C1238 a_4215_2153# sky130_fd_sc_hd__inv_1_0/Y 0
C1239 ui_in[1] sky130_fd_sc_hd__inv_1_0/A 0.1618f
C1240 a_12194_5909# a_10888_5837# 0
C1241 CLA_0/sky130_fd_sc_hd__and4_1_1/C CLA_0/sky130_fd_sc_hd__or4_1_0/B -0
C1242 a_2313_2157# sky130_fd_sc_hd__inv_1_0/Y 0.00666f
C1243 a_7944_2243# sky130_fd_sc_hd__fa_1_3/CIN 0.06773f
C1244 VDPWR a_12793_14007# 0
C1245 a_10121_2159# VDPWR 0.00104f
C1246 a_13029_14207# sky130_fd_sc_hd__inv_1_2/A 0.00913f
C1247 sky130_fd_sc_hd__inv_1_9/Y sky130_fd_sc_hd__inv_1_8/A 0
C1248 a_12559_4919# sky130_fd_sc_hd__inv_1_1/A 0
C1249 CLA_0/a_187_n2435# VDPWR 0.00364f
C1250 VDPWR a_14152_5917# 0.05342f
C1251 CLA_0/sky130_fd_sc_hd__or4_1_0/a_27_297# CLA_0/sky130_fd_sc_hd__or4_1_0/C -0
C1252 CLA_0/sky130_fd_sc_hd__or4_1_0/X CLA_0/sky130_fd_sc_hd__or4_1_0/a_27_297# 0.00887f
C1253 VDPWR a_10652_2159# 0.00629f
C1254 CLA_0/sky130_fd_sc_hd__and4_1_1/a_27_47# CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0.00369f
C1255 sky130_fd_sc_hd__fa_1_11/SUM a_7285_5493# 0
C1256 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_0/a_193_413# -0
C1257 uio_oe[5] uio_oe[4] 0.03102f
C1258 a_2049_1791# VDPWR 0
C1259 a_4084_5493# a_4477_5409# -0
C1260 a_9871_14979# a_9739_15799# 0
C1261 a_10289_1793# sky130_fd_sc_hd__inv_1_0/A 0
C1262 ui_in[1] ui_in[0] 5.54868f
C1263 a_7126_5409# VDPWR 0
C1264 VDPWR sky130_fd_sc_hd__fa_1_16/CIN 0.8062f
C1265 sky130_fd_sc_hd__fa_1_5/CIN a_11888_2243# 0.06767f
C1266 sky130_fd_sc_hd__mux2_1_0/S sky130_fd_sc_hd__fa_1_18/CIN 0.0303f
C1267 sky130_fd_sc_hd__fa_1_18/CIN a_14825_4547# 0.00339f
C1268 a_13029_14207# a_11949_13849# -0
C1269 sky130_fd_sc_hd__inv_1_7/A sky130_fd_sc_hd__inv_1_6/A 0.05615f
C1270 a_9287_5499# sky130_fd_sc_hd__fa_1_17/SUM 0
C1271 VDPWR a_10261_5837# 0
C1272 VDPWR a_5174_5409# 0
C1273 CLA_0/sky130_fd_sc_hd__or4_1_0/a_27_297# CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0
C1274 CLA_0/sky130_fd_sc_hd__and2_1_0/a_145_75# VDPWR 0.0031f
C1275 uio_in[2] uio_in[1] 0.03102f
C1276 VDPWR a_9871_14979# 0.12398f
C1277 a_9034_2159# sky130_fd_sc_hd__inv_1_0/A 0
C1278 sky130_fd_sc_hd__fa_1_12/CIN a_13186_4919# 0
C1279 a_8794_5415# sky130_fd_sc_hd__inv_1_1/A 0
C1280 a_17153_2243# VDPWR 0.04562f
C1281 sky130_fd_sc_hd__fa_1_18/CIN a_14152_5917# 0
C1282 VDPWR sky130_fd_sc_hd__mux4_1_0/a_834_97# 0
C1283 CLA_1/sky130_fd_sc_hd__xor2_1_0/X CLA_1/sky130_fd_sc_hd__or4_1_0/A -0
C1284 a_15681_4997# a_16847_4529# 0
C1285 sky130_fd_sc_hd__fa_1_7/CIN sky130_fd_sc_hd__fa_1_6/CIN 0
C1286 VDPWR CLA_0/a_197_n3749# 0.02361f
C1287 a_10357_5471# sky130_fd_sc_hd__inv_1_1/A 0
C1288 sky130_fd_sc_hd__inv_1_7/A sky130_fd_sc_hd__inv_1_9/A 0
C1289 VDPWR a_16033_2159# 0
C1290 a_12587_5825# sky130_fd_sc_hd__fa_1_16/CIN 0
C1291 sky130_fd_sc_hd__inv_1_0/Y a_4746_2153# 0
C1292 a_12823_4919# sky130_fd_sc_hd__fa_1_16/CIN 0
C1293 CLA_0/sky130_fd_sc_hd__and4_1_1/a_197_47# VDPWR 0.00158f
C1294 sky130_fd_sc_hd__fa_1_18/CIN sky130_fd_sc_hd__fa_1_16/CIN 0
C1295 a_15089_2243# sky130_fd_sc_hd__inv_1_0/A 0.00304f
C1296 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.02964f
C1297 CLA_0/sky130_fd_sc_hd__or4_1_0/A a_9749_14235# 0
C1298 uo_out[7] uo_out[6] 0.03102f
C1299 a_14908_5467# VDPWR 0.02801f
C1300 sky130_fd_sc_hd__fa_1_16/CIN sky130_fd_sc_hd__fa_1_16/SUM 0.04873f
C1301 CLA_1/sky130_fd_sc_hd__and4_1_0/B a_9629_14779# -0
C1302 a_14065_2159# sky130_fd_sc_hd__inv_1_0/A 0
C1303 a_14281_5467# sky130_fd_sc_hd__inv_1_1/A 0
C1304 CLA_0/sky130_fd_sc_hd__or2_1_0/A CLA_0/sky130_fd_sc_hd__or4_1_0/C -0
C1305 VDPWR a_12865_14007# 0
C1306 ui_in[5] ui_in[4] 0.03102f
C1307 a_10553_4963# sky130_fd_sc_hd__inv_1_1/A 0
C1308 CLA_1/sky130_fd_sc_hd__xor2_1_0/X a_12009_15689# -0.00369f
C1309 VDPWR a_10916_4597# 0.02835f
C1310 sky130_fd_sc_hd__mux2_1_0/S sky130_fd_sc_hd__mux2_1_0/A0 0.2153f
C1311 VDPWR a_9451_16343# 0.00472f
C1312 CLA_1/sky130_fd_sc_hd__or4_1_0/B VDPWR 0.34374f
C1313 VDPWR a_4309_5043# 0
C1314 VDPWR sky130_fd_sc_hd__fa_1_19/CIN 0.61872f
C1315 uo_out[2] uo_out[1] 0.03102f
C1316 VDPWR a_6071_1787# 0
C1317 ui_in[1] sky130_fd_sc_hd__inv_1_1/A 0.06114f
C1318 a_14377_5833# sky130_fd_sc_hd__inv_1_1/A 0
C1319 a_14908_5467# sky130_fd_sc_hd__fa_1_18/CIN 0
C1320 sky130_fd_sc_hd__fa_1_12/CIN a_12430_5003# 0
C1321 a_5080_1787# VDPWR 0
C1322 a_10160_5047# sky130_fd_sc_hd__inv_1_0/A 0
C1323 CLA_1/sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__inv_1_2/A 0.04052f
C1324 VDPWR a_13137_2243# 0.07855f
C1325 CLA_0/a_19_n2185# VDPWR 0.00529f
C1326 a_16539_5473# sky130_fd_sc_hd__inv_1_1/A 0
C1327 VDPWR a_8263_5049# 0
C1328 a_17395_5923# a_17703_4979# 0
C1329 sky130_fd_sc_hd__fa_1_5/CIN a_12281_2159# 0
C1330 a_9896_2243# a_11145_2243# -0.00146f
C1331 sky130_fd_sc_hd__mux2_1_0/a_535_374# sky130_fd_sc_hd__inv_1_1/A 0
C1332 CLA_0/sky130_fd_sc_hd__or4_1_0/B CLA_0/sky130_fd_sc_hd__or4_1_0/C -0
C1333 CLA_0/sky130_fd_sc_hd__or4_1_0/X CLA_0/sky130_fd_sc_hd__or4_1_0/B 0.03899f
C1334 a_2145_1791# VDPWR 0
C1335 CLA_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0
C1336 VDPWR a_9739_15799# 0.07542f
C1337 CLA_1/sky130_fd_sc_hd__xor2_1_0/X a_11777_15239# -0
C1338 a_6792_5043# VDPWR 0.02485f
C1339 sky130_fd_sc_hd__fa_1_15/CIN sky130_fd_sc_hd__inv_1_1/A 0.00685f
C1340 VDPWR sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.03032f
C1341 VDPWR a_14561_4913# 0
C1342 sky130_fd_sc_hd__fa_1_18/CIN sky130_fd_sc_hd__fa_1_19/CIN 0
C1343 VDPWR a_2343_5051# 0.01606f
C1344 a_6429_5043# sky130_fd_sc_hd__fa_1_9/CIN 0.00339f
C1345 a_9577_15377# a_9739_15799# -0
C1346 a_2145_2157# sky130_fd_sc_hd__inv_1_0/Y 0
C1347 a_8794_5049# sky130_fd_sc_hd__inv_1_1/A 0
C1348 sky130_fd_sc_hd__fa_1_4/SUM sky130_fd_sc_hd__inv_1_0/A 0.00121f
C1349 VDPWR a_13969_1793# 0
C1350 sky130_fd_sc_hd__fa_1_12/COUT sky130_fd_sc_hd__fa_1_14/SUM 0.00621f
C1351 sky130_fd_sc_hd__fa_1_10/SUM VDPWR 0.09157f
C1352 a_9579_12145# VDPWR 0.00291f
C1353 VDPWR a_4215_1787# 0
C1354 a_7191_2237# sky130_fd_sc_hd__inv_1_0/A 0.00307f
C1355 sky130_fd_sc_hd__mux2_1_0/S sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.05171f
C1356 a_16847_4895# sky130_fd_sc_hd__inv_1_1/A 0
C1357 VDPWR a_14930_1793# 0
C1358 a_16146_5923# a_15401_5917# 0.00354f
C1359 CLA_0/sky130_fd_sc_hd__and3_1_0/a_181_47# VDPWR 0.00109f
C1360 a_16297_1793# sky130_fd_sc_hd__inv_1_0/A 0
C1361 sky130_fd_sc_hd__mux4_1_0/a_1478_413# sky130_fd_sc_hd__inv_1_0/A 0.00234f
C1362 CLA_0/sky130_fd_sc_hd__or4_1_0/a_27_297# a_9749_14235# 0
C1363 a_9287_5499# sky130_fd_sc_hd__mux2_1_0/S 0.00783f
C1364 CLA_0/sky130_fd_sc_hd__or4_1_0/B CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0
C1365 a_9577_15377# VDPWR 0.0031f
C1366 a_14065_1793# sky130_fd_sc_hd__inv_1_0/A 0
C1367 VDPWR a_13284_5825# 0
C1368 a_6335_1787# sky130_fd_sc_hd__inv_1_0/A 0
C1369 VDPWR a_8169_2159# 0.00103f
C1370 a_12017_1793# sky130_fd_sc_hd__inv_1_0/A 0
C1371 uio_out[0] uo_out[7] 0.03102f
C1372 sky130_fd_sc_hd__inv_1_1/A sky130_fd_sc_hd__mux2_1_0/a_439_47# 0
C1373 CLA_0/sky130_fd_sc_hd__or2_1_0/a_68_297# CLA_0/sky130_fd_sc_hd__or4_1_0/a_27_297# -0
C1374 a_10025_2159# VDPWR 0
C1375 uio_in[4] uio_in[3] 0.03102f
C1376 VDPWR sky130_fd_sc_hd__inv_1_2/A 2.1608f
C1377 VDPWR a_16033_1793# 0
C1378 CLA_0/sky130_fd_sc_hd__and4_1_1/a_109_47# CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0
C1379 ui_in[0] sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.02482f
C1380 sky130_fd_sc_hd__fa_1_1/CIN a_3990_2237# 0.06765f
C1381 sky130_fd_sc_hd__fa_1_5/CIN a_12281_1793# 0.00339f
C1382 a_12823_4919# VDPWR 0.01428f
C1383 a_12587_5825# VDPWR 0.01457f
C1384 VDPWR sky130_fd_sc_hd__fa_1_18/CIN 0.57908f
C1385 a_7944_2243# a_9193_2243# -0.00146f
C1386 a_11381_5921# sky130_fd_sc_hd__fa_1_12/SUM 0
C1387 a_14432_4997# a_15681_4997# -0.00146f
C1388 ui_in[2] ui_in[3] 0.03102f
C1389 a_10121_1793# sky130_fd_sc_hd__inv_1_0/A 0
C1390 VDPWR a_3040_5417# 0
C1391 VDPWR a_10761_14767# 0.00202f
C1392 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__inv_1_6/A 0
C1393 a_6792_5409# VDPWR 0.00627f
C1394 VDPWR sky130_fd_sc_hd__fa_1_16/SUM 0.08488f
C1395 a_11949_13849# VDPWR 0.03598f
C1396 sky130_fd_sc_hd__fa_1_7/CIN a_14596_1793# 0
C1397 a_14233_2159# a_13840_2243# -0
C1398 sky130_fd_sc_hd__fa_1_19/CIN sky130_fd_sc_hd__mux2_1_0/A0 0
C1399 sky130_fd_sc_hd__fa_1_14/CIN a_13443_5909# 0
C1400 VDPWR a_4840_5409# 0.00656f
C1401 VDPWR a_9128_5415# 0
C1402 sky130_fd_sc_hd__fa_1_2/SUM a_7191_2237# -0
C1403 sky130_fd_sc_hd__fa_1_7/SUM sky130_fd_sc_hd__fa_1_7/CIN 0.05087f
C1404 ui_in[1] ua[0] 0.48906f
C1405 a_8700_2159# sky130_fd_sc_hd__inv_1_0/A 0
C1406 a_7285_5493# sky130_fd_sc_hd__fa_1_9/SUM -0
C1407 sky130_fd_sc_hd__inv_1_1/A a_15242_5467# 0
C1408 sky130_fd_sc_hd__mux2_1_0/S a_11381_5921# 0
C1409 sky130_fd_sc_hd__fa_1_14/CIN sky130_fd_sc_hd__inv_1_1/A 0.00398f
C1410 a_12644_1793# sky130_fd_sc_hd__inv_1_0/A 0
C1411 ua[4] a_15089_2243# 0
C1412 a_3990_2237# a_4383_1787# 0.01174f
C1413 CLA_1/sky130_fd_sc_hd__xor2_1_0/X a_10923_15189# -0
C1414 a_10160_5047# sky130_fd_sc_hd__inv_1_1/A 0
C1415 CLA_1/sky130_fd_sc_hd__and4_1_1/C a_11583_15239# -0
C1416 VDPWR sky130_fd_sc_hd__fa_1_4/CIN 0.55836f
C1417 VDPWR sky130_fd_sc_hd__fa_1_8/SUM 0.07919f
C1418 a_2049_2157# VDPWR 0
C1419 sky130_fd_sc_hd__fa_1_1/CIN sky130_fd_sc_hd__inv_1_0/Y 0.00472f
C1420 VDPWR a_2343_5417# 0.01298f
C1421 sky130_fd_sc_hd__inv_1_0/Y a_5942_2237# 0.001f
C1422 CLA_0/sky130_fd_sc_hd__and4_1_1/a_303_47# VDPWR 0.00104f
C1423 a_11888_2243# sky130_fd_sc_hd__inv_1_0/A 0.00211f
C1424 ui_in[6] ui_in[7] 0.03102f
C1425 VDPWR a_10888_5471# 0.02669f
C1426 sky130_fd_sc_hd__fa_1_1/CIN sky130_fd_sc_hd__fa_1_2/CIN 0
C1427 sky130_fd_sc_hd__mux2_1_0/a_76_199# sky130_fd_sc_hd__mux2_1_0/A0 0.01474f
C1428 sky130_fd_sc_hd__fa_1_2/CIN a_5942_2237# 0.0677f
C1429 sky130_fd_sc_hd__fa_1_3/CIN a_7191_2237# 0.00764f
C1430 CLA_0/a_187_n2185# VDPWR 0.02321f
C1431 sky130_fd_sc_hd__inv_1_2/Y CLA_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0
C1432 CLA_0/sky130_fd_sc_hd__and4_1_0/a_27_47# CLA_0/a_67_n1483# -0
C1433 CLA_1/sky130_fd_sc_hd__xor2_1_0/X a_11225_14223# -0
C1434 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__inv_1_0/A 0
C1435 a_4383_2153# a_4119_2153# 0
C1436 a_17153_2243# a_16994_2159# -0
C1437 a_12194_5909# a_13443_5909# -0.00146f
C1438 a_14545_5467# VDPWR 0.01734f
C1439 CLA_0/sky130_fd_sc_hd__or2_1_0/a_68_297# CLA_0/sky130_fd_sc_hd__or2_1_0/A 0
C1440 sky130_fd_sc_hd__mux2_1_0/S sky130_fd_sc_hd__fa_1_13/SUM -0
C1441 sky130_fd_sc_hd__fa_1_19/CIN sky130_fd_sc_hd__fa_1_19/SUM 0.05149f
C1442 ui_in[0] sky130_fd_sc_hd__mux4_1_0/a_668_97# 0.00464f
C1443 sky130_fd_sc_hd__fa_1_1/CIN a_4119_1787# 0
C1444 a_13969_2159# sky130_fd_sc_hd__inv_1_0/A 0
C1445 VDPWR sky130_fd_sc_hd__mux2_1_0/A0 0.4376f
C1446 a_15242_5833# sky130_fd_sc_hd__inv_1_1/A 0
C1447 a_12194_5909# sky130_fd_sc_hd__inv_1_1/A 0.0051f
C1448 VDPWR CLA_0/sky130_fd_sc_hd__and4_1_0/B 0.81349f
C1449 sky130_fd_sc_hd__inv_1_0/Y a_5080_2153# 0
C1450 a_11409_5047# sky130_fd_sc_hd__inv_1_0/A 0
C1451 a_8038_5499# a_7285_5493# 0.0035f
C1452 sky130_fd_sc_hd__mux2_1_0/S sky130_fd_sc_hd__mux2_1_0/A1 0.2868f
C1453 a_10385_4963# sky130_fd_sc_hd__inv_1_1/A 0
C1454 a_4383_1787# sky130_fd_sc_hd__inv_1_0/Y 0
C1455 sky130_fd_sc_hd__fa_1_6/CIN a_13137_2243# 0.00764f
C1456 VDPWR a_10553_4597# 0.02335f
C1457 CLA_0/sky130_fd_sc_hd__and4_1_1/C VDPWR 0.26677f
C1458 a_12978_1793# sky130_fd_sc_hd__inv_1_0/A 0
C1459 ui_in[0] sky130_fd_sc_hd__mux4_1_0/a_1290_413# 0.02515f
C1460 a_14377_5467# a_14152_5917# -0
C1461 a_16847_4529# sky130_fd_sc_hd__inv_1_0/A 0
C1462 CLA_0/sky130_fd_sc_hd__or4_1_0/B a_9749_14235# 0
C1463 a_14281_5833# sky130_fd_sc_hd__inv_1_1/A 0
C1464 VDPWR a_12419_5459# 0
C1465 a_11225_14223# a_10993_13773# -0
C1466 sky130_fd_sc_hd__inv_1_2/Y CLA_0/sky130_fd_sc_hd__and4_1_1/a_27_47# 0.00853f
C1467 a_14545_5467# sky130_fd_sc_hd__fa_1_18/CIN 0
C1468 sky130_fd_sc_hd__mux2_1_0/S a_16146_5923# 0
C1469 sky130_fd_sc_hd__fa_1_12/CIN sky130_fd_sc_hd__fa_1_12/SUM 0.05122f
C1470 sky130_fd_sc_hd__fa_1_6/CIN a_13969_1793# 0
C1471 CLA_0/sky130_fd_sc_hd__or4_1_0/X a_9871_14979# 0.00206f
C1472 a_11250_4597# sky130_fd_sc_hd__inv_1_0/A 0
C1473 a_4383_1787# a_4119_1787# 0
C1474 a_16539_5839# a_17395_5923# -0
C1475 sky130_fd_sc_hd__fa_1_11/SUM sky130_fd_sc_hd__inv_1_1/A 0.00121f
C1476 CLA_1/sky130_fd_sc_hd__xor2_1_0/X CLA_1/sky130_fd_sc_hd__or2_1_0/A -0
C1477 sky130_fd_sc_hd__fa_1_7/CIN a_15904_2243# 0.06765f
C1478 ua[1] 0 0.14696f
C1479 ua[2] 0 0.14696f
C1480 ua[3] 0 0.14696f
C1481 ua[4] 0 0.1448f
C1482 ua[5] 0 0.1448f
C1483 ua[6] 0 0.1449f
C1484 ua[7] 0 0.14552f
C1485 ena 0 0.07038f
C1486 clk 0 0.04288f
C1487 rst_n 0 0.04288f
C1488 ui_in[2] 0 0.04288f
C1489 ui_in[3] 0 0.04288f
C1490 ui_in[4] 0 0.04288f
C1491 ui_in[5] 0 0.04288f
C1492 ui_in[6] 0 0.04288f
C1493 ui_in[7] 0 0.04288f
C1494 uio_in[0] 0 0.04288f
C1495 uio_in[1] 0 0.04288f
C1496 uio_in[2] 0 0.04288f
C1497 uio_in[3] 0 0.04288f
C1498 uio_in[4] 0 0.04288f
C1499 uio_in[5] 0 0.04288f
C1500 uio_in[6] 0 0.04288f
C1501 uio_in[7] 0 0.04288f
C1502 uo_out[0] 0 0.04288f
C1503 uo_out[1] 0 0.04288f
C1504 uo_out[2] 0 0.04288f
C1505 uo_out[3] 0 0.04288f
C1506 uo_out[4] 0 0.04288f
C1507 uo_out[5] 0 0.04288f
C1508 uo_out[6] 0 0.04288f
C1509 uo_out[7] 0 0.04288f
C1510 uio_out[0] 0 0.04288f
C1511 uio_out[1] 0 0.04288f
C1512 uio_out[2] 0 0.04288f
C1513 uio_out[3] 0 0.04288f
C1514 uio_out[4] 0 0.04288f
C1515 uio_out[5] 0 0.04288f
C1516 uio_out[6] 0 0.04288f
C1517 uio_out[7] 0 0.04288f
C1518 uio_oe[0] 0 0.04288f
C1519 uio_oe[1] 0 0.04288f
C1520 uio_oe[2] 0 0.04288f
C1521 uio_oe[3] 0 0.04288f
C1522 uio_oe[4] 0 0.04288f
C1523 uio_oe[5] 0 0.04288f
C1524 uio_oe[6] 0 0.04288f
C1525 uio_oe[7] 0 0.07038f
C1526 a_15904_2243# 0 0.12936f
C1527 a_15089_2243# 0 0.26671f
C1528 a_13840_2243# 0 0.12858f
C1529 a_13137_2243# 0 0.2654f
C1530 a_11888_2243# 0 0.12885f
C1531 a_9896_2243# 0 0.12858f
C1532 a_9193_2243# 0 0.2654f
C1533 a_7944_2243# 0 0.12915f
C1534 a_5942_2237# 0 0.12819f
C1535 a_5239_2237# 0 0.2654f
C1536 a_3990_2237# 0 0.12941f
C1537 a_17153_2243# 0 0.27343f
C1538 sky130_fd_sc_hd__fa_1_7/CIN 0 0.58889f
C1539 sky130_fd_sc_hd__fa_1_6/CIN 0 0.52882f
C1540 sky130_fd_sc_hd__fa_1_5/CIN 0 0.54908f
C1541 a_11145_2243# 0 0.26591f
C1542 sky130_fd_sc_hd__fa_1_3/CIN 0 0.55449f
C1543 a_7191_2237# 0 0.26537f
C1544 sky130_fd_sc_hd__fa_1_2/CIN 0 0.52732f
C1545 sky130_fd_sc_hd__fa_1_1/CIN 0 0.58865f
C1546 a_1920_2241# 0 0.13344f
C1547 a_3169_2241# 0 0.26688f
C1548 VDPWR 0 0.28429p
C1549 sky130_fd_sc_hd__inv_1_0/Y 0 2.2293f
C1550 a_17703_4979# 0 0.267f
C1551 a_16454_4979# 0 0.128f
C1552 sky130_fd_sc_hd__fa_1_19/CIN 0 0.52835f
C1553 a_14432_4997# 0 0.12725f
C1554 a_15681_4997# 0 0.26489f
C1555 sky130_fd_sc_hd__fa_1_18/CIN 0 0.51698f
C1556 a_13679_5003# 0 0.26503f
C1557 a_12430_5003# 0 0.12883f
C1558 sky130_fd_sc_hd__fa_1_16/CIN 0 0.54105f
C1559 a_10160_5047# 0 0.1338f
C1560 a_11409_5047# 0 0.26105f
C1561 a_17395_5923# 0 0.27223f
C1562 a_16146_5923# 0 0.12888f
C1563 a_15401_5917# 0 0.26397f
C1564 sky130_fd_sc_hd__fa_1_14/CIN 0 0.3414f
C1565 a_14152_5917# 0 0.12861f
C1566 a_13443_5909# 0 0.26345f
C1567 a_12194_5909# 0 0.12922f
C1568 a_11381_5921# 0 0.26503f
C1569 a_10132_5921# 0 0.13251f
C1570 a_9287_5499# 0 0.27121f
C1571 a_8038_5499# 0 0.12915f
C1572 a_6036_5493# 0 0.12846f
C1573 a_5333_5493# 0 0.2654f
C1574 a_4084_5493# 0 0.12981f
C1575 sky130_fd_sc_hd__fa_1_9/COUT 0 0.55404f
C1576 a_7285_5493# 0 0.2656f
C1577 sky130_fd_sc_hd__fa_1_9/CIN 0 0.52729f
C1578 sky130_fd_sc_hd__fa_1_8/CIN 0 0.61983f
C1579 a_3199_5501# 0 0.26755f
C1580 a_1950_5501# 0 0.13325f
C1581 sky130_fd_sc_hd__inv_1_1/Y 0 2.29088f
C1582 a_11117_12361# 0 0.15959f
C1583 a_11165_13381# 0 0.15893f
C1584 a_13029_14207# 0 0.15924f
C1585 a_11949_13849# 0 0.15168f
C1586 a_11225_14223# 0 0.16017f
C1587 a_10923_15189# 0 0.1611f
C1588 a_12009_15689# 0 0.15596f
C1589 a_9739_15799# 0 0.1563f
C1590 a_9861_16543# 0 0.20741f
C1591 sky130_fd_sc_hd__fa_1_19/SUM 0 0.03818f
C1592 sky130_fd_sc_hd__mux2_1_0/A1 0 0.47115f
C1593 a_16847_4895# 0 0.01584f
C1594 a_17210_4895# 0 0.01578f
C1595 a_16847_4529# 0 0.00484f
C1596 a_17210_4529# 0 0.00345f
C1597 sky130_fd_sc_hd__fa_1_9/SUM 0 0.03738f
C1598 a_6429_5409# 0 0.01584f
C1599 a_6792_5409# 0 0.01578f
C1600 a_6429_5043# 0 0.00484f
C1601 a_6792_5043# 0 0.00345f
C1602 sky130_fd_sc_hd__fa_1_18/SUM 0 0.038f
C1603 a_14825_4913# 0 0.01584f
C1604 a_15188_4913# 0 0.01578f
C1605 a_14825_4547# 0 0.00484f
C1606 a_15188_4547# 0 0.00345f
C1607 sky130_fd_sc_hd__inv_1_1/A 0 7.12086f
C1608 sky130_fd_sc_hd__mux2_1_0/a_505_21# 0 0.24676f
C1609 sky130_fd_sc_hd__mux2_1_0/a_76_199# 0 0.13947f
C1610 sky130_fd_sc_hd__fa_1_8/SUM 0 0.03934f
C1611 a_4477_5409# 0 0.01584f
C1612 a_4840_5409# 0 0.01578f
C1613 a_4477_5043# 0 0.00484f
C1614 a_4840_5043# 0 0.00345f
C1615 sky130_fd_sc_hd__fa_1_17/SUM 0 0.09665f
C1616 a_10553_4963# 0 0.01584f
C1617 a_10916_4963# 0 0.01578f
C1618 a_10553_4597# 0 0.00484f
C1619 a_10916_4597# 0 0.00345f
C1620 sky130_fd_sc_hd__fa_1_7/SUM 0 0.03833f
C1621 sky130_fd_sc_hd__inv_1_0/A 0 8.84248f
C1622 a_16297_2159# 0 0.01584f
C1623 a_16660_2159# 0 0.01578f
C1624 a_16297_1793# 0 0.00484f
C1625 a_16660_1793# 0 0.00345f
C1626 sky130_fd_sc_hd__inv_1_11/A 0 0.37553f
C1627 sky130_fd_sc_hd__inv_1_9/Y 0 0.33162f
C1628 sky130_fd_sc_hd__fa_1_16/SUM 0 0.03939f
C1629 a_12823_4919# 0 0.01584f
C1630 a_13186_4919# 0 0.01578f
C1631 a_12823_4553# 0 0.00484f
C1632 a_13186_4553# 0 0.00345f
C1633 sky130_fd_sc_hd__fa_1_6/SUM 0 0.03738f
C1634 a_14233_2159# 0 0.01584f
C1635 a_14596_2159# 0 0.01578f
C1636 a_14233_1793# 0 0.00484f
C1637 a_14596_1793# 0 0.00345f
C1638 sky130_fd_sc_hd__fa_1_15/SUM 0 0.03797f
C1639 sky130_fd_sc_hd__mux2_1_0/A0 0 0.58507f
C1640 a_16539_5839# 0 0.01584f
C1641 a_16902_5839# 0 0.01578f
C1642 a_16539_5473# 0 0.00484f
C1643 a_16902_5473# 0 0.00345f
C1644 sky130_fd_sc_hd__fa_1_5/SUM 0 0.03791f
C1645 a_12281_2159# 0 0.01584f
C1646 a_12644_2159# 0 0.01578f
C1647 a_12281_1793# 0 0.00484f
C1648 a_12644_1793# 0 0.00345f
C1649 sky130_fd_sc_hd__fa_1_14/SUM 0 0.03751f
C1650 sky130_fd_sc_hd__fa_1_15/CIN 0 0.50457f
C1651 a_14545_5833# 0 0.01584f
C1652 a_14908_5833# 0 0.01578f
C1653 a_14545_5467# 0 0.00484f
C1654 a_14908_5467# 0 0.00345f
C1655 sky130_fd_sc_hd__fa_1_4/SUM 0 0.03738f
C1656 a_10289_2159# 0 0.01584f
C1657 a_10652_2159# 0 0.01578f
C1658 a_10289_1793# 0 0.00484f
C1659 a_10652_1793# 0 0.00345f
C1660 sky130_fd_sc_hd__fa_1_13/SUM 0 0.04554f
C1661 sky130_fd_sc_hd__fa_1_12/CIN 0 0.53079f
C1662 a_10525_5837# 0 0.01584f
C1663 a_10888_5837# 0 0.01578f
C1664 a_10525_5471# 0 0.00484f
C1665 a_10888_5471# 0 0.00345f
C1666 sky130_fd_sc_hd__fa_1_3/SUM 0 0.03806f
C1667 sky130_fd_sc_hd__fa_1_4/CIN 0 0.52882f
C1668 a_8337_2159# 0 0.01584f
C1669 a_8700_2159# 0 0.01578f
C1670 a_8337_1793# 0 0.00484f
C1671 a_8700_1793# 0 0.00345f
C1672 sky130_fd_sc_hd__fa_1_12/SUM 0 0.03865f
C1673 sky130_fd_sc_hd__fa_1_12/COUT 0 0.06859f
C1674 a_12587_5825# 0 0.01584f
C1675 a_12950_5825# 0 0.01578f
C1676 a_12587_5459# 0 0.00484f
C1677 a_12950_5459# 0 0.00345f
C1678 sky130_fd_sc_hd__fa_1_2/SUM 0 0.03738f
C1679 a_6335_2153# 0 0.01584f
C1680 a_6698_2153# 0 0.01578f
C1681 a_6335_1787# 0 0.00484f
C1682 a_6698_1787# 0 0.00345f
C1683 sky130_fd_sc_hd__fa_1_11/SUM 0 0.03806f
C1684 sky130_fd_sc_hd__mux2_1_0/S 0 1.14547f
C1685 a_8431_5415# 0 0.01584f
C1686 a_8794_5415# 0 0.01578f
C1687 a_8431_5049# 0 0.00484f
C1688 a_8794_5049# 0 0.00345f
C1689 sky130_fd_sc_hd__fa_1_1/SUM 0 0.03876f
C1690 a_4383_2153# 0 -0.02403f
C1691 a_4746_2153# 0 0.01578f
C1692 a_4383_1787# 0 -0.03724f
C1693 a_4746_1787# 0 0.00345f
C1694 sky130_fd_sc_hd__fa_1_10/SUM 0 0.04606f
C1695 a_2343_5417# 0 0.01584f
C1696 a_2706_5417# 0 0.01578f
C1697 a_2343_5051# 0 0.00484f
C1698 a_2706_5051# 0 0.00345f
C1699 sky130_fd_sc_hd__fa_1_0/SUM 0 0.0457f
C1700 a_2313_2157# 0 0.01584f
C1701 a_2676_2157# 0 0.01578f
C1702 a_2313_1791# 0 0.00484f
C1703 a_2676_1791# 0 0.00345f
C1704 a_9751_11003# 0 0.15405f
C1705 a_9873_11747# 0 0.20027f
C1706 a_9741_12567# 0 0.15062f
C1707 a_9863_13311# 0 0.19705f
C1708 a_9749_14235# 0 0.14822f
C1709 a_9871_14979# 0 0.19797f
C1710 a_9631_11547# 0 0.00137f
C1711 a_9629_14779# 0 0.00137f
C1712 a_9619_16343# 0 0.00137f
C1713 CLA_1/sky130_fd_sc_hd__or2_1_0/B 0 0.45897f
C1714 sky130_fd_sc_hd__inv_1_2/A 0 4.21407f
C1715 CLA_1/sky130_fd_sc_hd__or4_1_0/B 0 0.76691f
C1716 CLA_1/sky130_fd_sc_hd__or2_1_0/A 0 0.31659f
C1717 CLA_1/sky130_fd_sc_hd__xor2_1_0/X 0 1.57103f
C1718 CLA_1/sky130_fd_sc_hd__and4_1_0/B 0 0.65098f
C1719 CLA_1/sky130_fd_sc_hd__or4_1_0/A 0 0.31745f
C1720 CLA_1/sky130_fd_sc_hd__and4_1_1/C 0 0.30772f
C1721 CLA_1/sky130_fd_sc_hd__or4_1_0/C 0 1.1412f
C1722 a_9621_13111# 0 0.00137f
C1723 CLA_0/a_69_n4715# 0 0.1752f
C1724 CLA_0/a_n53_n3749# 0 0.24712f
C1725 CLA_0/a_59_n3151# 0 0.17114f
C1726 CLA_0/a_n63_n2185# 0 0.24424f
C1727 CLA_0/a_67_n1483# 0 0.17003f
C1728 CLA_0/a_n55_n517# 0 0.24496f
C1729 CLA_0/a_197_n3749# 0 0.00137f
C1730 CLA_0/a_195_n517# 0 0.00137f
C1731 CLA_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C1732 CLA_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.25457f
C1733 CLA_0/sky130_fd_sc_hd__or2_1_0/B 0 0.46058f
C1734 CLA_0/sky130_fd_sc_hd__and3_1_0/a_27_47# 0 0.17719f
C1735 CLA_0/sky130_fd_sc_hd__or4_1_0/X 0 2.79329f
C1736 CLA_0/sky130_fd_sc_hd__or4_1_0/B 0 0.82103f
C1737 CLA_0/sky130_fd_sc_hd__or4_1_0/a_27_297# 0 0.16291f
C1738 sky130_fd_sc_hd__inv_1_2/Y 0 2.40508f
C1739 CLA_0/sky130_fd_sc_hd__and4_1_1/a_27_47# 0 0.17489f
C1740 CLA_0/sky130_fd_sc_hd__or2_1_0/A 0 0.322f
C1741 CLA_0/sky130_fd_sc_hd__xor2_1_0/X 0 1.89172f
C1742 CLA_0/sky130_fd_sc_hd__and4_1_0/B 0 0.74819f
C1743 CLA_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 0 0.17489f
C1744 CLA_0/sky130_fd_sc_hd__or4_1_0/A 0 0.45644f
C1745 CLA_0/sky130_fd_sc_hd__or2_1_0/a_68_297# 0 0.15387f
C1746 CLA_0/sky130_fd_sc_hd__and4_1_1/C 0 0.33836f
C1747 CLA_0/sky130_fd_sc_hd__and2_1_5/a_59_75# 0 0.17706f
C1748 CLA_0/sky130_fd_sc_hd__or4_1_0/C 0 1.46406f
C1749 CLA_0/sky130_fd_sc_hd__and2_1_4/a_59_75# 0 0.17706f
C1750 CLA_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 0 0.17706f
C1751 CLA_0/a_187_n2185# 0 0.00137f
C1752 ua[0] 0 9.43909f
C1753 ui_in[1] 0 7.45535f
C1754 ui_in[0] 0 9.0828f
C1755 sky130_fd_sc_hd__mux4_1_0/a_834_97# 0 0.02499f
C1756 sky130_fd_sc_hd__mux4_1_0/a_668_97# 0 0.02039f
C1757 sky130_fd_sc_hd__mux4_1_0/a_27_47# 0 0.04207f
C1758 sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0 0.16413f
C1759 sky130_fd_sc_hd__mux4_1_0/a_1290_413# 0 0.2199f
C1760 sky130_fd_sc_hd__mux4_1_0/a_750_97# 0 0.04192f
C1761 sky130_fd_sc_hd__mux4_1_0/a_757_363# 0 0.00666f
C1762 sky130_fd_sc_hd__mux4_1_0/a_247_21# 0 0.34344f
C1763 sky130_fd_sc_hd__mux4_1_0/a_193_413# 0 0.00373f
C1764 sky130_fd_sc_hd__mux4_1_0/a_27_413# 0 0.02865f
C1765 sky130_fd_sc_hd__inv_1_9/A 0 0.45841f
C1766 sky130_fd_sc_hd__inv_1_8/A 0 0.38043f
C1767 sky130_fd_sc_hd__inv_1_7/A 0 0.32958f
C1768 sky130_fd_sc_hd__inv_1_6/A 0 0.33556f
C1769 sky130_fd_sc_hd__inv_1_5/A 0 0.33848f
C1770 sky130_fd_sc_hd__inv_1_4/A 0 0.40061f
.ends

