* SPICE3 file created from tt_um_ohmy90_adders.ext - technology: sky130A

.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
C0 VGND VPWR 0.03382f
C1 VPB A 0.04506f
C2 VPB VPWR 0.05448f
C3 VPB VGND 0.00948f
C4 Y A 0.0476f
C5 Y VPWR 0.12758f
C6 Y VGND 0.09984f
C7 Y VPB 0.01774f
C8 A VPWR 0.03703f
C9 VGND A 0.04004f
C10 VGND VNB 0.25113f
C11 Y VNB 0.0961f
C12 VPWR VNB 0.21892f
C13 A VNB 0.16664f
C14 VPB VNB 0.33898f
.ends

.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X a_1290_413#
+ a_757_363# a_1478_413# a_277_47# a_750_97# a_27_413# a_923_363# a_193_47# a_834_97#
+ a_247_21# a_668_97# a_193_413# a_27_47#
X0 a_277_47# a_247_21# a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VGND S0 a_247_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_834_97# a_247_21# a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=0.10795 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VGND A3 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1079 ps=1.36 w=0.42 l=0.15
X4 a_1290_413# S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_834_97# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_750_97# S0 a_757_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1079 ps=1.36 w=0.42 l=0.15
X7 a_27_47# S0 a_277_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.08523 ps=0.925 w=0.42 l=0.15
X8 X a_1478_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X9 VPWR A1 a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VPWR S0 a_247_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1079 pd=1.36 as=0.1083 ps=1.36 w=0.42 l=0.15
X11 X a_1478_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X12 a_193_47# A0 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_750_97# a_1290_413# a_1478_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2688 pd=2.12 as=0.09207 ps=0.99 w=0.42 l=0.15
X14 a_1478_413# S1 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09207 pd=0.99 as=0.1092 ps=1.36 w=0.42 l=0.15
X15 a_1290_413# S1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X16 a_277_47# a_247_21# a_193_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08523 pd=0.925 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_750_97# S0 a_668_97# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X18 a_923_363# a_247_21# a_750_97# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09013 pd=0.995 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 a_757_363# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X20 VPWR A3 a_923_363# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.09013 ps=0.995 w=0.42 l=0.15
X21 a_277_47# a_1290_413# a_1478_413# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.15102 ps=1.285 w=0.42 l=0.15
X22 a_193_413# A0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X23 a_193_413# S0 a_277_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1079 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X24 VGND A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X25 a_1478_413# S1 a_750_97# VNB sky130_fd_pr__nfet_01v8 ad=0.15102 pd=1.285 as=0.1092 ps=1.36 w=0.42 l=0.15
C0 A3 a_923_363# 0
C1 a_668_97# VPB 0.00146f
C2 A3 VPWR 0.012f
C3 A1 a_27_47# 0.03909f
C4 a_277_47# a_757_363# 0
C5 a_750_97# A2 0.01619f
C6 VGND a_27_413# 0.00189f
C7 a_750_97# VGND 0.05676f
C8 a_668_97# VPWR 0.00181f
C9 A2 a_757_363# 0.03541f
C10 VPB S1 0.21534f
C11 S0 a_27_413# 0
C12 a_750_97# S0 0.09449f
C13 A3 a_247_21# 0.07395f
C14 a_750_97# a_834_97# 0.0296f
C15 S0 a_757_363# 0.03305f
C16 VPWR S1 0.0409f
C17 a_668_97# a_247_21# 0.01881f
C18 a_834_97# a_757_363# 0.01352f
C19 a_277_47# A2 0.01375f
C20 X a_1290_413# 0.00208f
C21 a_277_47# VGND 0.41112f
C22 VPB a_27_47# 0.00324f
C23 a_247_21# S1 0
C24 a_277_47# S0 0.03381f
C25 A2 VGND 0.0122f
C26 a_277_47# a_834_97# 0.04391f
C27 VPWR a_27_47# 0.0018f
C28 A0 a_27_47# 0.04574f
C29 VGND S0 0.06675f
C30 X a_1478_413# 0.12698f
C31 a_834_97# A2 0.04394f
C32 VPB a_1290_413# 0.14223f
C33 a_834_97# VGND 0.09477f
C34 a_193_413# a_27_413# 0.05551f
C35 a_193_413# a_750_97# 0
C36 a_247_21# a_27_47# 0.0457f
C37 a_834_97# S0 0
C38 a_923_363# a_1290_413# 0
C39 A1 a_27_413# 0.0413f
C40 A1 a_750_97# 0
C41 VPWR a_1290_413# 0.0823f
C42 X a_750_97# 0
C43 a_1478_413# VPB 0.07712f
C44 a_247_21# a_1290_413# 0.00705f
C45 a_193_413# a_277_47# 0.0594f
C46 a_1478_413# VPWR 0.21151f
C47 A1 a_277_47# 0.00101f
C48 a_193_413# VGND 0
C49 VPB a_27_413# 0.02285f
C50 a_750_97# VPB 0.05933f
C51 a_277_47# X 0
C52 a_193_413# S0 0.01772f
C53 A1 VGND 0.01705f
C54 a_247_21# a_1478_413# 0
C55 VPB a_757_363# 0.0237f
C56 a_923_363# a_750_97# 0.00222f
C57 VPWR a_27_413# 0.08385f
C58 A0 a_27_413# 0.04892f
C59 a_750_97# A0 0
C60 a_750_97# VPWR 0.22609f
C61 X VGND 0.05939f
C62 a_923_363# a_757_363# 0.00988f
C63 VPWR a_757_363# 0.24812f
C64 A3 a_668_97# 0.0033f
C65 a_247_21# a_27_413# 0.00549f
C66 a_277_47# VPB 0.03677f
C67 a_750_97# a_247_21# 0.12371f
C68 A3 S1 0
C69 A2 VPB 0.07872f
C70 a_247_21# a_757_363# 0.02645f
C71 VGND VPB 0.01387f
C72 a_277_47# A0 0.05427f
C73 a_277_47# VPWR 0.05706f
C74 VPB S0 0.31074f
C75 A2 VPWR 0.0129f
C76 VGND VPWR 0.05896f
C77 A0 VGND 0.01709f
C78 a_834_97# VPB 0.00426f
C79 a_27_47# a_193_47# 0.00648f
C80 a_277_47# a_247_21# 0.35203f
C81 A0 S0 0.00186f
C82 VPWR S0 0.0687f
C83 A3 a_27_47# 0
C84 A1 a_193_413# 0
C85 a_923_363# a_834_97# 0
C86 a_247_21# A2 0.00145f
C87 a_834_97# VPWR 0
C88 a_247_21# VGND 0.09412f
C89 a_247_21# S0 0.39319f
C90 a_834_97# a_247_21# 0.02707f
C91 A3 a_1290_413# 0
C92 a_668_97# a_1290_413# 0
C93 a_193_413# VPB 0.01733f
C94 A1 VPB 0.0741f
C95 S1 a_1290_413# 0.15612f
C96 a_193_413# VPWR 0.18442f
C97 a_193_413# A0 0.00145f
C98 X VPB 0.01181f
C99 A1 A0 0.14123f
C100 A1 VPWR 0.01712f
C101 a_193_413# a_247_21# 0.09132f
C102 X VPWR 0.05937f
C103 a_1478_413# S1 0.00517f
C104 A3 a_750_97# 0.03406f
C105 A1 a_247_21# 0
C106 A3 a_757_363# 0.03224f
C107 a_668_97# a_750_97# 0.04662f
C108 X a_247_21# 0
C109 VPB VPWR 0.22689f
C110 A0 VPB 0.08019f
C111 a_277_47# a_193_47# 0
C112 a_750_97# S1 0.06323f
C113 A3 a_277_47# 0.0121f
C114 a_923_363# VPWR 0.00225f
C115 S1 a_757_363# 0.00151f
C116 A0 VPWR 0.01747f
C117 VGND a_193_47# 0.00175f
C118 A3 A2 0.15492f
C119 a_277_47# a_668_97# 0.02235f
C120 a_247_21# VPB 0.22297f
C121 A3 VGND 0.01161f
C122 A3 S0 0.00317f
C123 a_1478_413# a_1290_413# 0.10432f
C124 a_27_47# a_27_413# 0.00987f
C125 a_668_97# VGND 0.22352f
C126 a_247_21# VPWR 0.15063f
C127 a_277_47# S1 0.06116f
C128 a_247_21# A0 0.07359f
C129 A3 a_834_97# 0.03609f
C130 a_668_97# S0 0.03f
C131 A2 S1 0.06853f
C132 VGND S1 0.04087f
C133 a_668_97# a_834_97# 0.05583f
C134 a_750_97# a_1290_413# 0.17579f
C135 a_834_97# S1 0.00189f
C136 a_277_47# a_27_47# 0.08551f
C137 a_757_363# a_1290_413# 0.0098f
C138 VGND a_27_47# 0.22952f
C139 a_750_97# a_1478_413# 0.1456f
C140 S0 a_27_47# 0.01792f
C141 a_277_47# a_1290_413# 0.33858f
C142 A2 a_1290_413# 0.00165f
C143 VGND a_1290_413# 0.06373f
C144 a_750_97# a_27_413# 0
C145 a_277_47# a_1478_413# 0.09435f
C146 a_834_97# a_1290_413# 0.01242f
C147 a_750_97# a_757_363# 0.13413f
C148 a_1478_413# VGND 0.18885f
C149 X S1 0
C150 A3 VPB 0.07252f
C151 a_277_47# a_27_413# 0.05408f
C152 a_277_47# a_750_97# 0.26678f
C153 A0 a_193_47# 0
C154 VPWR a_193_47# 0
C155 VGND VNB 1.07507f
C156 X VNB 0.09236f
C157 S1 VNB 0.32062f
C158 A2 VNB 0.11249f
C159 A3 VNB 0.11926f
C160 S0 VNB 0.46486f
C161 VPWR VNB 0.86887f
C162 A0 VNB 0.10257f
C163 A1 VNB 0.17585f
C164 VPB VNB 1.9337f
C165 a_834_97# VNB 0.02499f
C166 a_668_97# VNB 0.02039f
C167 a_27_47# VNB 0.04207f
C168 a_1478_413# VNB 0.16413f
C169 a_1290_413# VNB 0.2199f
C170 a_750_97# VNB 0.04192f
C171 a_757_363# VNB 0.00666f
C172 a_277_47# VNB 0.07984f
C173 a_247_21# VNB 0.34344f
C174 a_193_413# VNB 0.00373f
C175 a_27_413# VNB 0.02865f
.ends

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X a_117_297# a_285_297# a_285_47#
+ a_35_297#
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
C0 a_285_297# a_35_297# 0.02504f
C1 a_285_47# VPWR 0
C2 B VPWR 0.07031f
C3 a_117_297# VPWR 0.00852f
C4 a_285_297# VGND 0.00394f
C5 a_285_47# B 0
C6 B a_117_297# 0.00777f
C7 X VPWR 0.05365f
C8 A VPWR 0.03484f
C9 VPB VPWR 0.06891f
C10 X a_285_47# 0.00206f
C11 X B 0.01488f
C12 X a_117_297# 0
C13 A B 0.22134f
C14 a_35_297# VPWR 0.09604f
C15 VPB B 0.06969f
C16 VGND VPWR 0.06426f
C17 a_285_47# a_35_297# 0.00723f
C18 B a_35_297# 0.203f
C19 a_35_297# a_117_297# 0.00641f
C20 A X 0.00166f
C21 VGND a_285_47# 0.00552f
C22 VGND B 0.03045f
C23 X VPB 0.01541f
C24 VGND a_117_297# 0.00177f
C25 A VPB 0.05101f
C26 X a_35_297# 0.166f
C27 A a_35_297# 0.06334f
C28 X VGND 0.1729f
C29 VPB a_35_297# 0.06993f
C30 a_285_297# VPWR 0.24631f
C31 A VGND 0.03254f
C32 VPB VGND 0.00696f
C33 a_285_297# B 0.05532f
C34 VGND a_35_297# 0.17666f
C35 a_285_297# X 0.07125f
C36 a_285_297# A 0.00749f
C37 a_285_297# VPB 0.01327f
C38 VGND VNB 0.43488f
C39 X VNB 0.06491f
C40 VPWR VNB 0.33278f
C41 A VNB 0.16672f
C42 B VNB 0.21337f
C43 VPB VNB 0.69336f
C44 a_285_297# VNB 0.00137f
C45 a_35_297# VNB 0.25457f
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X a_145_75# a_59_75#
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
C0 VPWR B 0.01175f
C1 VPB A 0.08057f
C2 X A 0
C3 A VGND 0.01472f
C4 VPB a_59_75# 0.05631f
C5 a_145_75# a_59_75# 0.00658f
C6 VPWR A 0.03623f
C7 X a_59_75# 0.10872f
C8 a_59_75# VGND 0.11564f
C9 VPWR a_59_75# 0.15028f
C10 VPB X 0.01265f
C11 a_145_75# X 0
C12 A B 0.09709f
C13 VPB VGND 0.008f
C14 a_145_75# VGND 0.00468f
C15 VPB VPWR 0.07293f
C16 X VGND 0.09933f
C17 a_145_75# VPWR 0
C18 X VPWR 0.11122f
C19 a_59_75# B 0.14331f
C20 VPWR VGND 0.04608f
C21 VPB B 0.06287f
C22 X B 0.00276f
C23 A a_59_75# 0.08088f
C24 VGND B 0.01146f
C25 VGND VNB 0.3114f
C26 X VNB 0.10018f
C27 B VNB 0.11287f
C28 A VNB 0.17379f
C29 VPWR VNB 0.27345f
C30 VPB VNB 0.51617f
C31 a_59_75# VNB 0.17706f
.ends

.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X a_150_297# a_68_297#
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
C0 B VPB 0.0462f
C1 X a_150_297# 0
C2 B X 0
C3 VPB A 0.03097f
C4 X A 0.01305f
C5 VGND VPWR 0.04645f
C6 a_68_297# VPB 0.06114f
C7 X a_68_297# 0.10534f
C8 B A 0.07509f
C9 VGND VPB 0.0112f
C10 VPB VPWR 0.08053f
C11 X VGND 0.11395f
C12 X VPWR 0.12857f
C13 a_68_297# a_150_297# 0.00477f
C14 B a_68_297# 0.09843f
C15 a_68_297# A 0.15786f
C16 VGND a_150_297# 0
C17 B VGND 0.04365f
C18 VPWR a_150_297# 0.00193f
C19 B VPWR 0.00855f
C20 X VPB 0.0209f
C21 VGND A 0.03465f
C22 A VPWR 0.00846f
C23 a_68_297# VGND 0.11796f
C24 a_68_297# VPWR 0.08898f
C25 VGND VNB 0.32043f
C26 X VNB 0.10095f
C27 A VNB 0.11072f
C28 B VNB 0.18272f
C29 VPWR VNB 0.26856f
C30 VPB VNB 0.51617f
C31 a_68_297# VNB 0.15387f
.ends

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X a_109_47# a_197_47# a_303_47#
+ a_27_47#
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.19627 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.19627 ps=1.33 w=0.65 l=0.15
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
C0 a_27_47# X 0.07537f
C1 VGND a_303_47# 0.00381f
C2 B VPB 0.06433f
C3 VGND B 0.04527f
C4 a_27_47# a_197_47# 0.00167f
C5 VPWR C 0.02103f
C6 A VPB 0.09066f
C7 A VGND 0.01512f
C8 VPWR VPB 0.07695f
C9 VPWR VGND 0.06618f
C10 A B 0.08391f
C11 a_197_47# C 0.00123f
C12 a_27_47# D 0.10658f
C13 X VPB 0.01107f
C14 VGND X 0.09025f
C15 VPWR a_303_47# 0
C16 VPWR B 0.02308f
C17 VGND a_197_47# 0.00387f
C18 a_27_47# a_109_47# 0.00578f
C19 A VPWR 0.044f
C20 a_197_47# B 0.00623f
C21 C D 0.18016f
C22 a_27_47# C 0.05159f
C23 D VPB 0.07823f
C24 VGND D 0.0898f
C25 VPWR X 0.09451f
C26 C a_109_47# 0
C27 a_27_47# VPB 0.08205f
C28 a_27_47# VGND 0.13176f
C29 VPWR a_197_47# 0
C30 VGND a_109_47# 0.00223f
C31 a_303_47# D 0.00119f
C32 a_27_47# a_303_47# 0.00119f
C33 a_27_47# B 0.12972f
C34 a_109_47# B 0.00153f
C35 C VPB 0.06088f
C36 VGND C 0.04082f
C37 a_27_47# A 0.15343f
C38 VPWR D 0.02073f
C39 a_27_47# VPWR 0.32628f
C40 VGND VPB 0.00852f
C41 C a_303_47# 0.00527f
C42 VPWR a_109_47# 0
C43 C B 0.16061f
C44 X D 0.00746f
C45 VGND VNB 0.39291f
C46 X VNB 0.09332f
C47 VPWR VNB 0.33454f
C48 D VNB 0.13027f
C49 C VNB 0.10983f
C50 B VNB 0.11212f
C51 A VNB 0.22098f
C52 VPB VNB 0.69336f
C53 a_27_47# VNB 0.17489f
.ends

.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X a_277_297# a_205_297# a_27_297#
+ a_109_297#
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.10187 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
C0 D VPWR 0.00503f
C1 X a_27_297# 0.0991f
C2 a_205_297# a_27_297# 0.00412f
C3 X VGND 0.03541f
C4 D A 0
C5 a_205_297# VGND 0
C6 VPWR C 0.00723f
C7 A C 0.02804f
C8 B a_277_297# 0
C9 a_109_297# a_27_297# 0.00695f
C10 B a_27_297# 0.15929f
C11 a_109_297# VGND 0
C12 VPB a_27_297# 0.05168f
C13 B VGND 0.01587f
C14 VPB VGND 0.00796f
C15 a_277_297# VPWR 0
C16 B X 0
C17 A a_277_297# 0
C18 VPWR a_27_297# 0.08397f
C19 VPB X 0.01089f
C20 VPWR VGND 0.05464f
C21 A a_27_297# 0.16258f
C22 D C 0.09543f
C23 A VGND 0.01596f
C24 X VPWR 0.08784f
C25 VPWR a_205_297# 0
C26 A X 0.00133f
C27 B VPB 0.10612f
C28 a_109_297# VPWR 0
C29 B VPWR 0.19276f
C30 VPB VPWR 0.07497f
C31 D a_27_297# 0.05404f
C32 a_277_297# C 0
C33 B A 0.06391f
C34 D VGND 0.05172f
C35 VPB A 0.03298f
C36 C a_27_297# 0.15835f
C37 C VGND 0.0191f
C38 A VPWR 0.00769f
C39 C a_205_297# 0.00261f
C40 a_277_297# a_27_297# 0.00876f
C41 a_277_297# VGND 0
C42 D B 0.00287f
C43 D VPB 0.04052f
C44 a_109_297# C 0.00356f
C45 VGND a_27_297# 0.23515f
C46 B C 0.09165f
C47 a_277_297# X 0
C48 VPB C 0.03382f
C49 VGND VNB 0.36697f
C50 X VNB 0.08835f
C51 A VNB 0.10929f
C52 C VNB 0.10488f
C53 D VNB 0.17526f
C54 B VNB 0.11467f
C55 VPWR VNB 0.28998f
C56 VPB VNB 0.60476f
C57 a_27_297# VNB 0.16291f
.ends

.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X a_181_47# a_109_47# a_27_47#
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14222 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14222 ps=1.335 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
C0 VPWR C 0.00464f
C1 VGND C 0.07031f
C2 B A 0.08692f
C3 B VPB 0.08363f
C4 VPWR VGND 0.04751f
C5 X C 0.01492f
C6 a_181_47# C 0.00151f
C7 a_27_47# C 0.1862f
C8 X VPWR 0.07662f
C9 X VGND 0.07078f
C10 a_181_47# VPWR 0
C11 a_181_47# VGND 0.00261f
C12 a_27_47# VPWR 0.14545f
C13 a_27_47# VGND 0.13361f
C14 B C 0.07462f
C15 VPB A 0.0426f
C16 VPWR a_109_47# 0
C17 a_109_47# VGND 0.00123f
C18 B VPWR 0.12845f
C19 X a_27_47# 0.08704f
C20 B VGND 0.00714f
C21 a_181_47# a_27_47# 0.00401f
C22 X B 0.00111f
C23 a_27_47# a_109_47# 0.00517f
C24 a_27_47# B 0.06246f
C25 VPB C 0.0347f
C26 VPWR A 0.01846f
C27 VGND A 0.01538f
C28 VPWR VPB 0.07946f
C29 VPB VGND 0.00604f
C30 a_27_47# A 0.15687f
C31 X VPB 0.01208f
C32 a_27_47# VPB 0.05008f
C33 a_109_47# A 0
C34 VGND VNB 0.30013f
C35 X VNB 0.09228f
C36 C VNB 0.12026f
C37 A VNB 0.17412f
C38 VPWR VNB 0.27425f
C39 B VNB 0.10179f
C40 VPB VNB 0.51617f
C41 a_27_47# VNB 0.17719f
.ends

.subckt CLA VNB sky130_fd_sc_hd__and4_1_1/a_303_47# sky130_fd_sc_hd__and4_1_0/VPB
+ sky130_fd_sc_hd__xor2_1_0/VPB sky130_fd_sc_hd__and2_1_5/VPB a_187_n2185# sky130_fd_sc_hd__and4_1_0/a_27_47#
+ sky130_fd_sc_hd__or4_1_0/D sky130_fd_sc_hd__or2_1_0/a_150_297# sky130_fd_sc_hd__and2_1_5/a_59_75#
+ sky130_fd_sc_hd__and4_1_1/VGND sky130_fd_sc_hd__and3_1_0/a_109_47# sky130_fd_sc_hd__or4_1_0/VPWR
+ sky130_fd_sc_hd__and3_1_0/a_181_47# sky130_fd_sc_hd__xor2_1_0/a_285_297# sky130_fd_sc_hd__and2_1_0/B
+ sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__or4_1_0/a_109_297# sky130_fd_sc_hd__and2_1_4/VPWR
+ sky130_fd_sc_hd__and2_1_0/A sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__and3_1_0/a_27_47#
+ a_187_n2435# sky130_fd_sc_hd__and3_1_0/VPWR sky130_fd_sc_hd__and4_1_1/VPB sky130_fd_sc_hd__xor2_1_0/a_285_47#
+ a_19_n2185# sky130_fd_sc_hd__xor2_1_0/a_35_297# sky130_fd_sc_hd__and2_1_4/a_145_75#
+ sky130_fd_sc_hd__and2_1_0/a_145_75# sky130_fd_sc_hd__and4_1_1/a_27_47# a_155_n4715#
+ sky130_fd_sc_hd__or4_1_0/VGND sky130_fd_sc_hd__or4_1_0/A sky130_fd_sc_hd__and2_1_4/VGND
+ sky130_fd_sc_hd__or2_1_0/a_68_297# sky130_fd_sc_hd__and2_1_0/VPB a_195_n517# a_n63_n2185#
+ a_197_n3749# sky130_fd_sc_hd__or4_1_0/X sky130_fd_sc_hd__and4_1_0/a_109_47# a_195_n767#
+ a_197_n3999# sky130_fd_sc_hd__and2_1_5/VPWR sky130_fd_sc_hd__and3_1_0/VGND sky130_fd_sc_hd__or2_1_0/VPWR
+ sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and2_1_5/a_145_75# sky130_fd_sc_hd__and2_1_0/a_59_75#
+ sky130_fd_sc_hd__and4_1_0/VPWR a_153_n1483# a_27_n517# a_69_n4715# sky130_fd_sc_hd__or2_1_0/B
+ sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__or4_1_0/a_277_297# sky130_fd_sc_hd__and4_1_0/a_197_47#
+ sky130_fd_sc_hd__and2_1_4/VPB sky130_fd_sc_hd__xor2_1_0/a_117_297# sky130_fd_sc_hd__and3_1_0/VPB
+ sky130_fd_sc_hd__and4_1_0/a_303_47# sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and4_1_1/a_109_47#
+ sky130_fd_sc_hd__or4_1_0/VPB sky130_fd_sc_hd__or4_1_0/a_27_297# a_29_n3749# sky130_fd_sc_hd__and2_1_5/VGND
+ sky130_fd_sc_hd__or4_1_0/a_205_297# sky130_fd_sc_hd__and2_1_4/a_59_75# sky130_fd_sc_hd__or2_1_0/VGND
+ a_n53_n3749# a_n55_n517# sky130_fd_sc_hd__and4_1_1/A sky130_fd_sc_hd__xor2_1_0/B
+ sky130_fd_sc_hd__and4_1_0/VGND sky130_fd_sc_hd__xor2_1_0/A sky130_fd_sc_hd__or4_1_0/C
+ a_67_n1483# sky130_fd_sc_hd__and4_1_1/VPWR a_59_n3151# sky130_fd_sc_hd__xor2_1_0/X
+ sky130_fd_sc_hd__and4_1_1/a_197_47# VPB X B a_145_n3151# A
Xsky130_fd_sc_hd__xor2_1_3 A B A VNB VPB B X a_19_n2185# a_187_n2185# a_187_n2435#
+ a_n63_n2185# sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__and2_1_0 sky130_fd_sc_hd__and2_1_0/A sky130_fd_sc_hd__and2_1_0/B
+ sky130_fd_sc_hd__and2_1_0/A VNB sky130_fd_sc_hd__and2_1_0/VPB sky130_fd_sc_hd__and2_1_0/B
+ sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and2_1_0/a_145_75# sky130_fd_sc_hd__and2_1_0/a_59_75#
+ sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_1 A B A VNB VPB B X a_153_n1483# a_67_n1483# sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_3 A B A VNB VPB B X a_145_n3151# a_59_n3151# sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_2 A B A VNB VPB B X a_155_n4715# a_69_n4715# sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_4 X X sky130_fd_sc_hd__and2_1_4/VGND VNB sky130_fd_sc_hd__and2_1_4/VPB
+ sky130_fd_sc_hd__and2_1_4/VPWR sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__and2_1_4/a_145_75#
+ sky130_fd_sc_hd__and2_1_4/a_59_75# sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_5 X X sky130_fd_sc_hd__and2_1_5/VGND VNB sky130_fd_sc_hd__and2_1_5/VPB
+ sky130_fd_sc_hd__and2_1_5/VPWR sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and2_1_5/a_145_75#
+ sky130_fd_sc_hd__and2_1_5/a_59_75# sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__or2_1_0 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__or2_1_0/VGND
+ VNB sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__or2_1_0/VPWR sky130_fd_sc_hd__or4_1_0/A
+ sky130_fd_sc_hd__or2_1_0/a_150_297# sky130_fd_sc_hd__or2_1_0/a_68_297# sky130_fd_sc_hd__or2_1
Xsky130_fd_sc_hd__and4_1_0 X sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__xor2_1_0/X
+ X sky130_fd_sc_hd__and4_1_0/VGND VNB sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__and4_1_0/VPWR
+ sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__and4_1_0/a_109_47# sky130_fd_sc_hd__and4_1_0/a_197_47#
+ sky130_fd_sc_hd__and4_1_0/a_303_47# sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__and4_1
Xsky130_fd_sc_hd__and4_1_1 sky130_fd_sc_hd__and4_1_1/A X sky130_fd_sc_hd__and4_1_1/C
+ sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and4_1_1/VGND VNB sky130_fd_sc_hd__and4_1_1/VPB
+ sky130_fd_sc_hd__and4_1_1/VPWR sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__and4_1_1/a_109_47#
+ sky130_fd_sc_hd__and4_1_1/a_197_47# sky130_fd_sc_hd__and4_1_1/a_303_47# sky130_fd_sc_hd__and4_1_1/a_27_47#
+ sky130_fd_sc_hd__and4_1
Xsky130_fd_sc_hd__or4_1_0 sky130_fd_sc_hd__or4_1_0/A sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__or4_1_0/C
+ sky130_fd_sc_hd__or4_1_0/D sky130_fd_sc_hd__or4_1_0/VGND VNB sky130_fd_sc_hd__or4_1_0/VPB
+ sky130_fd_sc_hd__or4_1_0/VPWR sky130_fd_sc_hd__or4_1_0/X sky130_fd_sc_hd__or4_1_0/a_277_297#
+ sky130_fd_sc_hd__or4_1_0/a_205_297# sky130_fd_sc_hd__or4_1_0/a_27_297# sky130_fd_sc_hd__or4_1_0/a_109_297#
+ sky130_fd_sc_hd__or4_1
Xsky130_fd_sc_hd__and3_1_0 X X X sky130_fd_sc_hd__and3_1_0/VGND VNB sky130_fd_sc_hd__and3_1_0/VPB
+ sky130_fd_sc_hd__and3_1_0/VPWR sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__and3_1_0/a_181_47#
+ sky130_fd_sc_hd__and3_1_0/a_109_47# sky130_fd_sc_hd__and3_1_0/a_27_47# sky130_fd_sc_hd__and3_1
Xsky130_fd_sc_hd__xor2_1_0 sky130_fd_sc_hd__xor2_1_0/A sky130_fd_sc_hd__xor2_1_0/B
+ sky130_fd_sc_hd__xor2_1_0/A VNB sky130_fd_sc_hd__xor2_1_0/VPB sky130_fd_sc_hd__xor2_1_0/B
+ sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__xor2_1_0/a_117_297# sky130_fd_sc_hd__xor2_1_0/a_285_297#
+ sky130_fd_sc_hd__xor2_1_0/a_285_47# sky130_fd_sc_hd__xor2_1_0/a_35_297# sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_1 A B A VNB VPB B X a_27_n517# a_195_n517# a_195_n767# a_n55_n517#
+ sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_2 A B A VNB VPB B X a_29_n3749# a_197_n3749# a_197_n3999#
+ a_n53_n3749# sky130_fd_sc_hd__xor2_1
C0 a_n55_n517# sky130_fd_sc_hd__and4_1_0/B 0.0065f
C1 X sky130_fd_sc_hd__and3_1_0/a_181_47# 0.00275f
C2 sky130_fd_sc_hd__and3_1_0/VPWR X 0.34434f
C3 sky130_fd_sc_hd__or2_1_0/VGND sky130_fd_sc_hd__and3_1_0/a_27_47# 0
C4 X sky130_fd_sc_hd__and4_1_1/VPWR -0.00415f
C5 sky130_fd_sc_hd__and3_1_0/VPB sky130_fd_sc_hd__or2_1_0/VGND 0.00189f
C6 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and4_1_1/VPWR -0.00444f
C7 B sky130_fd_sc_hd__xor2_1_0/VPB 0
C8 sky130_fd_sc_hd__and3_1_0/a_27_47# sky130_fd_sc_hd__and3_1_0/VGND -0.00436f
C9 sky130_fd_sc_hd__and3_1_0/VPB sky130_fd_sc_hd__and3_1_0/VGND -0.00287f
C10 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and2_1_4/VPB 0
C11 a_197_n3749# A 0
C12 sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__and4_1_0/VGND 0.00246f
C13 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__or2_1_0/A 0.00329f
C14 a_67_n1483# B 0.05542f
C15 a_69_n4715# VPB 0
C16 a_n63_n2185# X 0.01073f
C17 sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__or4_1_0/C 0
C18 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__or4_1_0/VGND 0.14621f
C19 X sky130_fd_sc_hd__and4_1_0/VPWR 0.05837f
C20 sky130_fd_sc_hd__or2_1_0/a_68_297# sky130_fd_sc_hd__or4_1_0/a_27_297# 0
C21 sky130_fd_sc_hd__and3_1_0/a_27_47# sky130_fd_sc_hd__and2_1_4/a_59_75# 0
C22 sky130_fd_sc_hd__and4_1_0/VPWR sky130_fd_sc_hd__and4_1_1/C 0.01347f
C23 X sky130_fd_sc_hd__and4_1_1/VPB 0.00801f
C24 sky130_fd_sc_hd__xor2_1_0/B sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.04603f
C25 sky130_fd_sc_hd__and3_1_0/VPB sky130_fd_sc_hd__and2_1_4/a_59_75# 0
C26 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and2_1_0/A 0.03609f
C27 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and4_1_1/VPB 0.00112f
C28 sky130_fd_sc_hd__and4_1_1/a_109_47# sky130_fd_sc_hd__and4_1_1/VGND -0
C29 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and3_1_0/VGND 0
C30 X sky130_fd_sc_hd__and4_1_0/a_27_47# 0.06054f
C31 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C32 A sky130_fd_sc_hd__xor2_1_0/a_35_297# 0
C33 sky130_fd_sc_hd__and4_1_0/a_303_47# sky130_fd_sc_hd__xor2_1_0/X 0.00175f
C34 sky130_fd_sc_hd__and2_1_0/VPB sky130_fd_sc_hd__xor2_1_0/B 0.00406f
C35 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__and4_1_0/a_109_47# 0
C36 A a_187_n2435# 0.0022f
C37 sky130_fd_sc_hd__or4_1_0/a_277_297# sky130_fd_sc_hd__or4_1_0/VGND -0
C38 sky130_fd_sc_hd__or2_1_0/VGND sky130_fd_sc_hd__or2_1_0/a_150_297# -0
C39 sky130_fd_sc_hd__and3_1_0/VPWR VPB 0
C40 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__and4_1_0/VGND 0.06679f
C41 sky130_fd_sc_hd__and2_1_0/VPB A 0
C42 sky130_fd_sc_hd__and4_1_1/VPWR sky130_fd_sc_hd__and4_1_1/VGND -0.04789f
C43 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__and2_1_5/a_59_75# 0
C44 sky130_fd_sc_hd__and3_1_0/a_27_47# sky130_fd_sc_hd__and2_1_4/VPWR 0
C45 sky130_fd_sc_hd__and3_1_0/VPB sky130_fd_sc_hd__and2_1_4/VPWR 0
C46 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__or2_1_0/VPWR 0.00192f
C47 a_19_n2185# B 0.00416f
C48 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and2_1_0/B 0.01218f
C49 sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__and4_1_0/VGND -0.00404f
C50 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__or4_1_0/D 0.01853f
C51 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and2_1_4/a_59_75# 0
C52 VPB sky130_fd_sc_hd__xor2_1_0/A 0
C53 sky130_fd_sc_hd__and3_1_0/VPWR a_187_n2185# 0
C54 sky130_fd_sc_hd__xor2_1_0/a_35_297# sky130_fd_sc_hd__xor2_1_0/a_285_297# 0
C55 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and2_1_5/VPB 0.00629f
C56 a_n63_n2185# VPB 0.00419f
C57 a_n55_n517# sky130_fd_sc_hd__xor2_1_0/X 0
C58 sky130_fd_sc_hd__xor2_1_0/VPB sky130_fd_sc_hd__xor2_1_0/B 0.00802f
C59 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__or4_1_0/VPWR 0
C60 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__or4_1_0/B 0
C61 sky130_fd_sc_hd__and4_1_0/VPWR VPB 0
C62 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__and4_1_1/a_197_47# 0
C63 sky130_fd_sc_hd__or4_1_0/C B 0
C64 A sky130_fd_sc_hd__xor2_1_0/VPB 0
C65 a_27_n517# X 0
C66 B sky130_fd_sc_hd__xor2_1_0/B 0
C67 sky130_fd_sc_hd__or4_1_0/VPWR sky130_fd_sc_hd__or4_1_0/VPB -0.00543f
C68 sky130_fd_sc_hd__and4_1_1/VPB sky130_fd_sc_hd__and4_1_1/VGND -0.0052f
C69 sky130_fd_sc_hd__and3_1_0/a_109_47# sky130_fd_sc_hd__and3_1_0/VGND -0
C70 VPB sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C71 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and2_1_4/VPWR 0
C72 B A 1.17029f
C73 a_197_n3999# A 0.0022f
C74 sky130_fd_sc_hd__or2_1_0/VPWR sky130_fd_sc_hd__and4_1_0/VGND 0.00285f
C75 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__or4_1_0/a_109_297# 0
C76 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__or4_1_0/a_27_297# 0
C77 sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__and2_1_5/a_59_75# 0
C78 a_67_n1483# A 0.02856f
C79 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__or4_1_0/a_205_297# 0
C80 sky130_fd_sc_hd__and2_1_0/a_59_75# sky130_fd_sc_hd__xor2_1_0/A 0
C81 sky130_fd_sc_hd__or4_1_0/D sky130_fd_sc_hd__and4_1_0/VGND 0
C82 a_69_n4715# a_n53_n3749# 0.00144f
C83 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__or2_1_0/A 0
C84 X sky130_fd_sc_hd__and4_1_1/C 0.19117f
C85 sky130_fd_sc_hd__and4_1_0/VPWR sky130_fd_sc_hd__or4_1_0/A 0
C86 sky130_fd_sc_hd__and4_1_0/VPWR sky130_fd_sc_hd__and2_1_5/VGND 0.06986f
C87 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and2_1_0/A 0
C88 sky130_fd_sc_hd__xor2_1_0/B sky130_fd_sc_hd__xor2_1_0/a_117_297# 0.00416f
C89 X sky130_fd_sc_hd__and4_1_0/a_109_47# 0.00198f
C90 sky130_fd_sc_hd__or4_1_0/A sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C91 B sky130_fd_sc_hd__and4_1_0/VGND 0
C92 sky130_fd_sc_hd__and4_1_0/VPWR sky130_fd_sc_hd__and4_1_0/a_197_47# -0
C93 sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__and4_1_0/B 0.0108f
C94 a_67_n1483# sky130_fd_sc_hd__and4_1_0/VGND 0
C95 sky130_fd_sc_hd__or2_1_0/a_68_297# sky130_fd_sc_hd__or2_1_0/A 0.08751f
C96 sky130_fd_sc_hd__and3_1_0/VPWR sky130_fd_sc_hd__or2_1_0/B 0.04682f
C97 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.00153f
C98 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__or4_1_0/X 0.00162f
C99 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__and2_1_5/a_145_75# 0
C100 a_19_n2185# A -0
C101 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and2_1_0/VPB 0.00562f
C102 sky130_fd_sc_hd__or4_1_0/VGND sky130_fd_sc_hd__or2_1_0/a_68_297# 0
C103 sky130_fd_sc_hd__and2_1_5/a_59_75# B 0
C104 sky130_fd_sc_hd__and2_1_4/a_145_75# sky130_fd_sc_hd__and2_1_4/VPWR -0
C105 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__or2_1_0/VPB 0
C106 a_n63_n2185# a_n53_n3749# 0.00102f
C107 sky130_fd_sc_hd__or2_1_0/B a_n63_n2185# 0
C108 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and2_1_5/VPB 0.0094f
C109 X VPB 0.07236f
C110 X sky130_fd_sc_hd__and4_1_1/VGND -0.0125f
C111 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__or4_1_0/B 0.04169f
C112 sky130_fd_sc_hd__and3_1_0/VPWR sky130_fd_sc_hd__or2_1_0/VGND 0.00385f
C113 sky130_fd_sc_hd__and2_1_0/a_145_75# sky130_fd_sc_hd__and2_1_0/A 0.00152f
C114 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and4_1_1/VGND 0.19171f
C115 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__and4_1_1/a_303_47# 0
C116 A sky130_fd_sc_hd__xor2_1_0/B 0
C117 a_195_n517# X 0.01091f
C118 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__or4_1_0/VPB 0.01252f
C119 sky130_fd_sc_hd__and3_1_0/VPWR sky130_fd_sc_hd__and3_1_0/VGND -0.03312f
C120 sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C121 sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__and3_1_0/a_27_47# 0
C122 sky130_fd_sc_hd__or2_1_0/VPWR sky130_fd_sc_hd__or2_1_0/a_68_297# -0.00741f
C123 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__xor2_1_0/VPB 0
C124 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__and2_1_4/VPB 0
C125 sky130_fd_sc_hd__or4_1_0/D sky130_fd_sc_hd__or2_1_0/a_68_297# 0
C126 X a_187_n2185# 0.01155f
C127 sky130_fd_sc_hd__and4_1_0/B B 0.01591f
C128 sky130_fd_sc_hd__and4_1_1/A sky130_fd_sc_hd__and2_1_0/A 0
C129 sky130_fd_sc_hd__and4_1_0/B a_67_n1483# 0.00159f
C130 sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__and4_1_1/a_27_47# 0
C131 X sky130_fd_sc_hd__or4_1_0/A 0.00571f
C132 sky130_fd_sc_hd__and2_1_5/VPB sky130_fd_sc_hd__and4_1_1/a_27_47# 0
C133 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__or2_1_0/A 0.00515f
C134 X sky130_fd_sc_hd__and2_1_5/VGND 0.08784f
C135 X sky130_fd_sc_hd__and2_1_0/a_59_75# 0.00215f
C136 a_n63_n2185# sky130_fd_sc_hd__and3_1_0/VGND 0
C137 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and2_1_5/VGND 0.01061f
C138 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__and4_1_1/a_27_47# 0.00909f
C139 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__and4_1_0/VGND 0
C140 sky130_fd_sc_hd__and3_1_0/VPWR sky130_fd_sc_hd__and2_1_4/a_59_75# 0
C141 sky130_fd_sc_hd__xor2_1_0/B sky130_fd_sc_hd__xor2_1_0/a_285_297# 0.00746f
C142 sky130_fd_sc_hd__or4_1_0/VPB sky130_fd_sc_hd__or2_1_0/A 0
C143 X sky130_fd_sc_hd__and4_1_0/a_197_47# 0.00174f
C144 A sky130_fd_sc_hd__and4_1_0/VGND 0.00151f
C145 A sky130_fd_sc_hd__xor2_1_0/a_285_297# 0
C146 a_145_n3151# A 0.00152f
C147 sky130_fd_sc_hd__and4_1_0/a_303_47# sky130_fd_sc_hd__and4_1_0/VPWR -0
C148 sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__xor2_1_0/X 0.00937f
C149 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__and3_1_0/VGND 0
C150 a_59_n3151# a_69_n4715# 0
C151 sky130_fd_sc_hd__or2_1_0/a_150_297# sky130_fd_sc_hd__or2_1_0/A 0.00183f
C152 sky130_fd_sc_hd__and2_1_0/B sky130_fd_sc_hd__xor2_1_0/A 0.19937f
C153 sky130_fd_sc_hd__or4_1_0/VPB sky130_fd_sc_hd__or4_1_0/VGND -0.00395f
C154 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.0029f
C155 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and2_1_0/VPB 0.00261f
C156 a_n55_n517# sky130_fd_sc_hd__xor2_1_0/A 0
C157 sky130_fd_sc_hd__and4_1_1/A sky130_fd_sc_hd__and2_1_5/VPB 0
C158 sky130_fd_sc_hd__and3_1_0/a_27_47# B 0
C159 sky130_fd_sc_hd__and4_1_1/A sky130_fd_sc_hd__or4_1_0/B 0
C160 sky130_fd_sc_hd__and3_1_0/VPB B 0
C161 sky130_fd_sc_hd__and2_1_5/VPWR sky130_fd_sc_hd__and2_1_5/a_59_75# -0.00969f
C162 VPB a_187_n2185# -0
C163 a_n55_n517# a_n63_n2185# 0
C164 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__or2_1_0/VPWR 0
C165 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__and2_1_4/VGND 0.01004f
C166 X a_n53_n3749# 0.00394f
C167 sky130_fd_sc_hd__or2_1_0/B X 0.09665f
C168 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__or4_1_0/D 0
C169 sky130_fd_sc_hd__and4_1_0/VPWR sky130_fd_sc_hd__or4_1_0/VPWR 0
C170 sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__and4_1_1/C 0
C171 sky130_fd_sc_hd__and2_1_0/a_59_75# VPB 0.0016f
C172 sky130_fd_sc_hd__and2_1_5/VGND VPB 0
C173 a_195_n767# X 0
C174 sky130_fd_sc_hd__or4_1_0/VPWR sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C175 a_195_n517# sky130_fd_sc_hd__and2_1_0/a_59_75# 0
C176 X sky130_fd_sc_hd__and2_1_4/VPB 0.03834f
C177 sky130_fd_sc_hd__or2_1_0/VPWR sky130_fd_sc_hd__or2_1_0/a_150_297# -0
C178 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__xor2_1_0/B 0
C179 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__xor2_1_0/VPB 0.00903f
C180 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and2_1_5/VPWR 0.00455f
C181 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__and2_1_4/VPWR 0
C182 sky130_fd_sc_hd__and4_1_1/A sky130_fd_sc_hd__or2_1_0/A 0
C183 a_59_n3151# a_n63_n2185# 0.00144f
C184 sky130_fd_sc_hd__and2_1_5/VPWR sky130_fd_sc_hd__and4_1_1/a_197_47# 0
C185 sky130_fd_sc_hd__and4_1_0/B A 0.00988f
C186 sky130_fd_sc_hd__xor2_1_0/X B 0
C187 sky130_fd_sc_hd__xor2_1_0/A sky130_fd_sc_hd__and2_1_0/A 0.00306f
C188 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__or4_1_0/a_27_297# 0
C189 sky130_fd_sc_hd__and2_1_5/a_59_75# sky130_fd_sc_hd__and4_1_0/VGND 0
C190 sky130_fd_sc_hd__xor2_1_0/X a_67_n1483# 0
C191 sky130_fd_sc_hd__or2_1_0/VPWR sky130_fd_sc_hd__and4_1_1/a_27_47# 0
C192 X sky130_fd_sc_hd__or2_1_0/VGND 0.00322f
C193 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__or2_1_0/a_68_297# 0.00327f
C194 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__and4_1_1/a_109_47# 0
C195 sky130_fd_sc_hd__xor2_1_0/B sky130_fd_sc_hd__xor2_1_0/a_285_47# -0
C196 X sky130_fd_sc_hd__and3_1_0/VGND 0.1323f
C197 sky130_fd_sc_hd__and4_1_0/a_303_47# X 0.00226f
C198 a_69_n4715# a_197_n3749# 0
C199 sky130_fd_sc_hd__and4_1_1/A sky130_fd_sc_hd__and2_1_0/VPB 0
C200 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and4_1_0/VGND 0.04218f
C201 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__and4_1_1/VPWR 0.00963f
C202 a_n53_n3749# VPB 0.00422f
C203 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__xor2_1_0/a_285_297# 0
C204 sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__and4_1_1/VGND 0
C205 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__xor2_1_0/a_117_297# 0
C206 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__and3_1_0/a_27_47# 0
C207 sky130_fd_sc_hd__and3_1_0/VPB sky130_fd_sc_hd__or4_1_0/C 0
C208 X sky130_fd_sc_hd__and2_1_0/B 0.00148f
C209 X sky130_fd_sc_hd__and2_1_4/a_59_75# 0.06657f
C210 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__or4_1_0/X 0.00286f
C211 sky130_fd_sc_hd__and3_1_0/a_27_47# A 0.00153f
C212 sky130_fd_sc_hd__or2_1_0/a_68_297# sky130_fd_sc_hd__and4_1_0/VGND 0.00157f
C213 sky130_fd_sc_hd__and2_1_5/VPWR sky130_fd_sc_hd__and2_1_5/a_145_75# -0
C214 a_n55_n517# X 0.00926f
C215 sky130_fd_sc_hd__and4_1_0/VPWR sky130_fd_sc_hd__and2_1_5/VPB 0
C216 a_n55_n517# sky130_fd_sc_hd__and4_1_1/C 0
C217 sky130_fd_sc_hd__and4_1_0/VPWR sky130_fd_sc_hd__or4_1_0/B 0.00504f
C218 sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__and4_1_0/a_27_47# 0.00132f
C219 sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__or4_1_0/A 0
C220 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and2_1_5/a_59_75# 0.00451f
C221 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__and4_1_1/VPB 0.00459f
C222 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C223 X sky130_fd_sc_hd__and2_1_4/VPWR 0.13242f
C224 X sky130_fd_sc_hd__or4_1_0/a_27_297# 0
C225 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__xor2_1_0/B 0.03047f
C226 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__xor2_1_0/X 0
C227 a_n63_n2185# a_197_n3749# 0
C228 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and2_1_5/VPWR 0.1083f
C229 sky130_fd_sc_hd__and3_1_0/a_27_47# sky130_fd_sc_hd__and4_1_0/VGND 0
C230 sky130_fd_sc_hd__and3_1_0/VPB sky130_fd_sc_hd__and4_1_0/VGND 0.00717f
C231 sky130_fd_sc_hd__and2_1_5/VPWR sky130_fd_sc_hd__and4_1_1/a_303_47# 0
C232 X a_29_n3749# 0
C233 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__or4_1_0/VPB 0.00355f
C234 sky130_fd_sc_hd__xor2_1_0/X A 0
C235 a_59_n3151# X 0.0142f
C236 sky130_fd_sc_hd__and2_1_0/VPB sky130_fd_sc_hd__and4_1_1/VPWR 0
C237 sky130_fd_sc_hd__and4_1_0/VPWR sky130_fd_sc_hd__or2_1_0/A 0.00913f
C238 sky130_fd_sc_hd__or4_1_0/A sky130_fd_sc_hd__or2_1_0/VGND 0.01452f
C239 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__or2_1_0/a_150_297# 0
C240 X sky130_fd_sc_hd__and2_1_0/A 0.02789f
C241 VPB sky130_fd_sc_hd__and2_1_0/B 0.00134f
C242 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and2_1_0/A 0
C243 sky130_fd_sc_hd__xor2_1_0/A sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.03404f
C244 VPB sky130_fd_sc_hd__and2_1_4/a_59_75# 0
C245 a_195_n517# sky130_fd_sc_hd__and2_1_0/B 0
C246 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__and4_1_0/a_27_47# 0.00364f
C247 a_69_n4715# B 0.06183f
C248 sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__and4_1_0/VPWR -0
C249 sky130_fd_sc_hd__and2_1_0/VPB sky130_fd_sc_hd__xor2_1_0/A 0.01565f
C250 a_n55_n517# VPB 0.00367f
C251 A a_153_n1483# 0.00151f
C252 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__or2_1_0/a_68_297# 0
C253 sky130_fd_sc_hd__and2_1_5/a_59_75# sky130_fd_sc_hd__and3_1_0/a_27_47# 0
C254 sky130_fd_sc_hd__and2_1_5/VPWR sky130_fd_sc_hd__and4_1_1/a_27_47# 0
C255 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and4_1_0/VGND 0.03811f
C256 sky130_fd_sc_hd__and3_1_0/VPB sky130_fd_sc_hd__and2_1_5/a_59_75# 0
C257 a_n55_n517# a_195_n517# 0
C258 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__xor2_1_0/a_285_297# 0.0032f
C259 sky130_fd_sc_hd__or4_1_0/VGND sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C260 VPB sky130_fd_sc_hd__and2_1_4/VPWR 0
C261 sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__and2_1_4/VPB 0
C262 sky130_fd_sc_hd__and2_1_4/VGND sky130_fd_sc_hd__and3_1_0/a_27_47# 0
C263 sky130_fd_sc_hd__and2_1_0/a_59_75# sky130_fd_sc_hd__and2_1_0/B 0.05693f
C264 a_n55_n517# a_187_n2185# 0
C265 sky130_fd_sc_hd__and3_1_0/a_109_47# A 0
C266 sky130_fd_sc_hd__or2_1_0/a_150_297# sky130_fd_sc_hd__and4_1_0/VGND 0
C267 sky130_fd_sc_hd__and3_1_0/VPWR B 0.00199f
C268 X sky130_fd_sc_hd__or2_1_0/VPB 0.00576f
C269 a_59_n3151# VPB 0.00186f
C270 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__or2_1_0/VPB 0
C271 X sky130_fd_sc_hd__and2_1_5/VPB 0.03446f
C272 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and3_1_0/a_27_47# 0
C273 sky130_fd_sc_hd__and3_1_0/VPB sky130_fd_sc_hd__and4_1_0/B 0.00114f
C274 sky130_fd_sc_hd__or2_1_0/VPWR sky130_fd_sc_hd__and4_1_1/VPB 0
C275 sky130_fd_sc_hd__and2_1_5/VPB sky130_fd_sc_hd__and4_1_1/C 0.00946f
C276 a_n55_n517# sky130_fd_sc_hd__and2_1_0/a_59_75# 0
C277 a_n55_n517# sky130_fd_sc_hd__and2_1_5/VGND 0
C278 X sky130_fd_sc_hd__or4_1_0/B 0.00752f
C279 sky130_fd_sc_hd__xor2_1_0/VPB sky130_fd_sc_hd__xor2_1_0/A -0
C280 sky130_fd_sc_hd__or4_1_0/VPWR sky130_fd_sc_hd__or4_1_0/A 0.01499f
C281 sky130_fd_sc_hd__and4_1_0/VPWR sky130_fd_sc_hd__or4_1_0/D 0
C282 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__and4_1_1/C 0.00425f
C283 sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__or2_1_0/VGND 0.05365f
C284 sky130_fd_sc_hd__or2_1_0/VPWR sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C285 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and2_1_5/a_145_75# 0
C286 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and2_1_5/a_59_75# 0.03095f
C287 sky130_fd_sc_hd__and4_1_1/A sky130_fd_sc_hd__and2_1_5/VPWR 0
C288 VPB sky130_fd_sc_hd__and2_1_0/A 0.00317f
C289 B sky130_fd_sc_hd__xor2_1_0/A 0.01159f
C290 sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__and3_1_0/VGND 0.00866f
C291 sky130_fd_sc_hd__or4_1_0/D sky130_fd_sc_hd__and4_1_0/a_27_47# 0.00134f
C292 a_59_n3151# a_187_n2185# 0
C293 sky130_fd_sc_hd__and3_1_0/a_27_47# sky130_fd_sc_hd__or2_1_0/a_68_297# 0
C294 sky130_fd_sc_hd__or4_1_0/a_109_297# sky130_fd_sc_hd__or4_1_0/A 0.00226f
C295 sky130_fd_sc_hd__or4_1_0/A sky130_fd_sc_hd__or4_1_0/a_27_297# 0.11968f
C296 a_n63_n2185# B 0.04714f
C297 sky130_fd_sc_hd__and2_1_4/VPB sky130_fd_sc_hd__and3_1_0/VGND 0.00107f
C298 X a_197_n3749# 0.01127f
C299 sky130_fd_sc_hd__and4_1_0/VPWR B 0.00173f
C300 a_n63_n2185# a_67_n1483# 0.00115f
C301 B sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C302 sky130_fd_sc_hd__and4_1_0/VPWR a_67_n1483# 0
C303 X sky130_fd_sc_hd__or2_1_0/A 0.04432f
C304 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__xor2_1_0/X 0.3542f
C305 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and4_1_1/a_197_47# 0
C306 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__or2_1_0/A 0.00427f
C307 a_67_n1483# sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C308 sky130_fd_sc_hd__and2_1_0/a_59_75# sky130_fd_sc_hd__and2_1_0/A 0.0274f
C309 sky130_fd_sc_hd__xor2_1_0/A sky130_fd_sc_hd__xor2_1_0/a_117_297# -0
C310 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__and4_1_0/a_109_47# 0
C311 sky130_fd_sc_hd__and4_1_0/VPB X 0.02141f
C312 a_69_n4715# A 0.02702f
C313 X sky130_fd_sc_hd__or4_1_0/VGND 0
C314 sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__and4_1_1/VGND 0
C315 sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__and4_1_1/C 0
C316 sky130_fd_sc_hd__and3_1_0/VPB sky130_fd_sc_hd__and3_1_0/a_27_47# -0
C317 sky130_fd_sc_hd__and2_1_5/VPB sky130_fd_sc_hd__and4_1_1/VGND 0
C318 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__or2_1_0/a_68_297# 0
C319 X sky130_fd_sc_hd__xor2_1_0/a_35_297# 0
C320 sky130_fd_sc_hd__and2_1_5/VPWR sky130_fd_sc_hd__and4_1_1/a_109_47# 0
C321 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__and4_1_1/VGND 0.04642f
C322 a_n55_n517# a_195_n767# 0
C323 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__xor2_1_0/a_285_47# 0
C324 X a_187_n2435# 0
C325 sky130_fd_sc_hd__and3_1_0/VPWR sky130_fd_sc_hd__or4_1_0/C 0
C326 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and4_1_1/a_27_47# 0
C327 a_n63_n2185# a_19_n2185# -0
C328 sky130_fd_sc_hd__and3_1_0/a_181_47# A 0
C329 sky130_fd_sc_hd__and4_1_1/A sky130_fd_sc_hd__and2_1_5/a_59_75# 0
C330 sky130_fd_sc_hd__and2_1_4/VPB sky130_fd_sc_hd__and2_1_4/VPWR -0
C331 sky130_fd_sc_hd__and2_1_4/a_59_75# sky130_fd_sc_hd__and3_1_0/VGND 0
C332 a_59_n3151# a_n53_n3749# 0
C333 X sky130_fd_sc_hd__or2_1_0/VPWR 0.00738f
C334 sky130_fd_sc_hd__or4_1_0/A sky130_fd_sc_hd__or2_1_0/VPB 0.01132f
C335 a_27_n517# B 0.00416f
C336 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and2_1_0/a_145_75# 0
C337 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__or2_1_0/VPWR 0
C338 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and3_1_0/a_27_47# 0
C339 sky130_fd_sc_hd__and3_1_0/VPB sky130_fd_sc_hd__xor2_1_0/X 0
C340 sky130_fd_sc_hd__and2_1_5/VPB sky130_fd_sc_hd__and2_1_5/VGND -0.0046f
C341 X sky130_fd_sc_hd__or4_1_0/D 0
C342 sky130_fd_sc_hd__xor2_1_0/B sky130_fd_sc_hd__xor2_1_0/A 0.06504f
C343 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__or4_1_0/A 0.3049f
C344 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__and4_1_1/VGND 0.00602f
C345 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__and2_1_5/VGND 0.00369f
C346 a_59_n3151# sky130_fd_sc_hd__and2_1_4/VPB 0
C347 sky130_fd_sc_hd__or2_1_0/a_68_297# sky130_fd_sc_hd__and4_1_1/a_27_47# 0
C348 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and2_1_5/a_145_75# 0
C349 A sky130_fd_sc_hd__xor2_1_0/A 0
C350 X sky130_fd_sc_hd__xor2_1_0/VPB 0
C351 a_n63_n2185# A 0.03465f
C352 sky130_fd_sc_hd__and2_1_4/VPWR sky130_fd_sc_hd__and3_1_0/VGND 0.07231f
C353 sky130_fd_sc_hd__and4_1_1/A sky130_fd_sc_hd__and4_1_0/B 0
C354 sky130_fd_sc_hd__and3_1_0/VPWR sky130_fd_sc_hd__and4_1_0/VGND 0.123f
C355 X B 0.38254f
C356 VPB sky130_fd_sc_hd__xor2_1_0/a_35_297# 0
C357 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C358 a_195_n517# sky130_fd_sc_hd__xor2_1_0/a_35_297# 0
C359 X a_67_n1483# 0.01753f
C360 A sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C361 a_n55_n517# sky130_fd_sc_hd__and2_1_0/B 0
C362 sky130_fd_sc_hd__or4_1_0/A sky130_fd_sc_hd__or2_1_0/A 0.04854f
C363 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and4_1_1/a_303_47# 0.00135f
C364 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__or4_1_0/VPB 0
C365 sky130_fd_sc_hd__xor2_1_0/A sky130_fd_sc_hd__xor2_1_0/a_285_297# -0
C366 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__and4_1_0/a_197_47# 0
C367 sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__or2_1_0/VPB 0.00342f
C368 sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__or4_1_0/A 0
C369 sky130_fd_sc_hd__or2_1_0/VPWR sky130_fd_sc_hd__and4_1_1/VGND 0.02529f
C370 sky130_fd_sc_hd__and2_1_4/a_59_75# sky130_fd_sc_hd__and2_1_4/VPWR -0.00137f
C371 sky130_fd_sc_hd__or4_1_0/A sky130_fd_sc_hd__or4_1_0/VGND 0.06333f
C372 sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__and2_1_5/VGND 0.00281f
C373 sky130_fd_sc_hd__and4_1_0/VPWR sky130_fd_sc_hd__and4_1_0/VGND -0.03588f
C374 sky130_fd_sc_hd__and3_1_0/VPWR sky130_fd_sc_hd__and2_1_5/a_59_75# 0
C375 sky130_fd_sc_hd__and2_1_0/a_59_75# sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.00144f
C376 sky130_fd_sc_hd__and4_1_0/VGND sky130_fd_sc_hd__and4_1_0/a_27_47# -0.00307f
C377 a_59_n3151# sky130_fd_sc_hd__and2_1_4/a_59_75# 0
C378 sky130_fd_sc_hd__or4_1_0/VPWR sky130_fd_sc_hd__or4_1_0/a_109_297# -0
C379 sky130_fd_sc_hd__or4_1_0/VPWR sky130_fd_sc_hd__or4_1_0/a_27_297# -0.01391f
C380 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and4_1_1/a_27_47# 0.12778f
C381 sky130_fd_sc_hd__and2_1_0/B sky130_fd_sc_hd__and2_1_0/A 0.03965f
C382 X a_19_n2185# 0
C383 VPB B 0.08228f
C384 a_27_n517# A -0
C385 a_195_n517# B 0.00754f
C386 sky130_fd_sc_hd__or2_1_0/VGND sky130_fd_sc_hd__or2_1_0/VPB -0.00683f
C387 sky130_fd_sc_hd__or4_1_0/A sky130_fd_sc_hd__or2_1_0/VPWR 0.06282f
C388 a_67_n1483# VPB 0.00126f
C389 sky130_fd_sc_hd__and3_1_0/VPWR sky130_fd_sc_hd__and4_1_0/B 0
C390 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and4_1_1/VPWR 0
C391 sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__or2_1_0/A 0.12539f
C392 sky130_fd_sc_hd__or4_1_0/D sky130_fd_sc_hd__or4_1_0/A 0.02169f
C393 a_n55_n517# sky130_fd_sc_hd__and2_1_0/A 0
C394 a_195_n517# a_67_n1483# 0
C395 sky130_fd_sc_hd__and4_1_1/a_197_47# sky130_fd_sc_hd__and4_1_1/VPWR -0
C396 a_59_n3151# sky130_fd_sc_hd__and2_1_4/VPWR 0
C397 sky130_fd_sc_hd__and4_1_0/VPWR sky130_fd_sc_hd__and2_1_5/a_59_75# 0
C398 sky130_fd_sc_hd__and2_1_5/a_59_75# sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C399 B a_187_n2185# 0.00766f
C400 X sky130_fd_sc_hd__or4_1_0/C 0.07546f
C401 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__xor2_1_0/A 0.00331f
C402 sky130_fd_sc_hd__and2_1_0/a_59_75# sky130_fd_sc_hd__xor2_1_0/VPB 0
C403 X sky130_fd_sc_hd__and2_1_5/VPWR 0.25442f
C404 a_67_n1483# a_187_n2185# 0
C405 sky130_fd_sc_hd__and3_1_0/VPWR sky130_fd_sc_hd__or2_1_0/a_68_297# 0
C406 sky130_fd_sc_hd__and2_1_5/VPWR sky130_fd_sc_hd__and4_1_1/C 0.072f
C407 sky130_fd_sc_hd__and4_1_1/A sky130_fd_sc_hd__xor2_1_0/X 0.03531f
C408 X A 0.25089f
C409 sky130_fd_sc_hd__and2_1_0/a_59_75# B 0
C410 A sky130_fd_sc_hd__and4_1_0/a_109_47# 0
C411 sky130_fd_sc_hd__and2_1_0/a_59_75# a_67_n1483# 0
C412 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and4_1_0/VPWR 0.0319f
C413 sky130_fd_sc_hd__or2_1_0/VGND sky130_fd_sc_hd__or2_1_0/A 0.0375f
C414 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and4_1_1/VPB 0
C415 sky130_fd_sc_hd__or4_1_0/a_205_297# sky130_fd_sc_hd__or4_1_0/A 0.00121f
C416 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and4_1_0/a_27_47# 0.03791f
C417 sky130_fd_sc_hd__xor2_1_0/A sky130_fd_sc_hd__xor2_1_0/a_285_47# 0.0022f
C418 sky130_fd_sc_hd__and4_1_0/a_303_47# sky130_fd_sc_hd__or2_1_0/A 0
C419 a_n55_n517# sky130_fd_sc_hd__and2_1_5/VPB 0
C420 sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__or2_1_0/VPWR -0.00376f
C421 sky130_fd_sc_hd__and3_1_0/VPWR sky130_fd_sc_hd__and3_1_0/a_27_47# -0.00561f
C422 sky130_fd_sc_hd__and3_1_0/VPB sky130_fd_sc_hd__and3_1_0/VPWR -0.00263f
C423 sky130_fd_sc_hd__or4_1_0/VPWR sky130_fd_sc_hd__or4_1_0/B 0.18975f
C424 X sky130_fd_sc_hd__and4_1_0/VGND 0.26798f
C425 sky130_fd_sc_hd__and4_1_1/A sky130_fd_sc_hd__and4_1_1/a_27_47# 0.00637f
C426 X a_145_n3151# 0
C427 sky130_fd_sc_hd__and4_1_1/VPB sky130_fd_sc_hd__or2_1_0/a_68_297# 0
C428 sky130_fd_sc_hd__or2_1_0/a_68_297# sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C429 sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__or4_1_0/a_27_297# 0
C430 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__or4_1_0/a_27_297# 0.0078f
C431 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and4_1_1/a_109_47# 0
C432 VPB sky130_fd_sc_hd__xor2_1_0/B 0
C433 sky130_fd_sc_hd__and2_1_5/VPWR sky130_fd_sc_hd__and4_1_1/VGND 0.0025f
C434 a_195_n517# sky130_fd_sc_hd__xor2_1_0/B 0
C435 a_n53_n3749# B 0.04711f
C436 VPB A 0.05774f
C437 a_n63_n2185# sky130_fd_sc_hd__and3_1_0/a_27_47# 0
C438 sky130_fd_sc_hd__and3_1_0/VPB a_n63_n2185# 0
C439 a_195_n517# A 0
C440 sky130_fd_sc_hd__or2_1_0/VGND sky130_fd_sc_hd__or2_1_0/VPWR -0.03781f
C441 sky130_fd_sc_hd__and4_1_0/VPWR sky130_fd_sc_hd__and3_1_0/a_27_47# 0
C442 B sky130_fd_sc_hd__and2_1_4/VPB 0
C443 sky130_fd_sc_hd__and3_1_0/VPWR sky130_fd_sc_hd__xor2_1_0/X 0
C444 sky130_fd_sc_hd__or4_1_0/VPWR sky130_fd_sc_hd__or2_1_0/A 0
C445 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and4_1_1/VPWR 0.26064f
C446 X sky130_fd_sc_hd__and2_1_5/a_59_75# 0.10648f
C447 sky130_fd_sc_hd__and4_1_1/a_303_47# sky130_fd_sc_hd__and4_1_1/VPWR -0
C448 a_27_n517# sky130_fd_sc_hd__and4_1_0/B 0
C449 sky130_fd_sc_hd__and2_1_5/a_59_75# sky130_fd_sc_hd__and4_1_1/C 0.00218f
C450 sky130_fd_sc_hd__and2_1_0/B sky130_fd_sc_hd__xor2_1_0/a_35_297# 0
C451 sky130_fd_sc_hd__and3_1_0/a_27_47# sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C452 sky130_fd_sc_hd__and3_1_0/VPB sky130_fd_sc_hd__and4_1_0/a_27_47# 0.00142f
C453 A a_187_n2185# 0
C454 sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__or4_1_0/VPWR 0
C455 a_59_n3151# a_197_n3749# 0
C456 X sky130_fd_sc_hd__and2_1_4/VGND 0.06329f
C457 sky130_fd_sc_hd__and2_1_0/VPB sky130_fd_sc_hd__and2_1_0/B 0.01331f
C458 sky130_fd_sc_hd__or4_1_0/VPWR sky130_fd_sc_hd__or4_1_0/VGND -0.0364f
C459 sky130_fd_sc_hd__or4_1_0/a_109_297# sky130_fd_sc_hd__or2_1_0/A 0
C460 sky130_fd_sc_hd__or2_1_0/A sky130_fd_sc_hd__or4_1_0/a_27_297# 0.00196f
C461 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__or4_1_0/A 0.1873f
C462 sky130_fd_sc_hd__and2_1_0/a_59_75# sky130_fd_sc_hd__xor2_1_0/B 0
C463 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__xor2_1_0/A 0.03369f
C464 a_n55_n517# sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.00102f
C465 sky130_fd_sc_hd__and2_1_5/VPWR sky130_fd_sc_hd__and2_1_5/VGND -0.03541f
C466 sky130_fd_sc_hd__and2_1_5/VGND A 0
C467 sky130_fd_sc_hd__and2_1_0/a_59_75# A 0
C468 a_n55_n517# sky130_fd_sc_hd__and2_1_0/VPB 0
C469 sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__or4_1_0/a_27_297# 0
C470 sky130_fd_sc_hd__or4_1_0/a_109_297# sky130_fd_sc_hd__or4_1_0/VGND -0
C471 sky130_fd_sc_hd__or4_1_0/VGND sky130_fd_sc_hd__or4_1_0/a_27_297# -0.00274f
C472 X sky130_fd_sc_hd__and4_1_0/B 0.65102f
C473 A sky130_fd_sc_hd__and4_1_0/a_197_47# 0
C474 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and4_1_0/VPWR 0.13704f
C475 X sky130_fd_sc_hd__and4_1_1/a_197_47# 0
C476 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and4_1_1/C 0
C477 sky130_fd_sc_hd__and4_1_1/a_27_47# sky130_fd_sc_hd__and4_1_1/VPWR -0.01767f
C478 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and4_1_1/VPB 0.02121f
C479 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and4_1_1/a_197_47# 0.00243f
C480 sky130_fd_sc_hd__or4_1_0/a_277_297# sky130_fd_sc_hd__or4_1_0/A 0.00184f
C481 sky130_fd_sc_hd__and4_1_0/VPWR sky130_fd_sc_hd__or4_1_0/VPB 0
C482 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and4_1_0/a_27_47# 0.03227f
C483 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and4_1_0/a_109_47# 0.00197f
C484 sky130_fd_sc_hd__or4_1_0/VPB sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C485 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__or2_1_0/VPB 0
C486 sky130_fd_sc_hd__and2_1_0/B sky130_fd_sc_hd__xor2_1_0/VPB 0
C487 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__and2_1_5/VPB 0
C488 X sky130_fd_sc_hd__or2_1_0/a_68_297# 0.0035f
C489 sky130_fd_sc_hd__and3_1_0/VPWR sky130_fd_sc_hd__and3_1_0/a_109_47# -0
C490 a_155_n4715# B 0
C491 sky130_fd_sc_hd__or4_1_0/VPWR sky130_fd_sc_hd__or4_1_0/D -0.00384f
C492 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__or2_1_0/a_68_297# 0
C493 B sky130_fd_sc_hd__and2_1_0/B 0.00168f
C494 sky130_fd_sc_hd__and2_1_5/a_59_75# VPB 0
C495 sky130_fd_sc_hd__and2_1_5/a_59_75# sky130_fd_sc_hd__and4_1_1/VGND 0
C496 sky130_fd_sc_hd__and2_1_0/a_59_75# sky130_fd_sc_hd__xor2_1_0/a_285_297# 0
C497 sky130_fd_sc_hd__and2_1_0/A sky130_fd_sc_hd__xor2_1_0/a_35_297# 0
C498 B sky130_fd_sc_hd__and2_1_4/a_59_75# 0
C499 sky130_fd_sc_hd__or2_1_0/VPWR sky130_fd_sc_hd__or4_1_0/a_27_297# 0
C500 sky130_fd_sc_hd__and4_1_0/VGND sky130_fd_sc_hd__and4_1_0/a_197_47# -0
C501 a_67_n1483# sky130_fd_sc_hd__and2_1_0/B 0
C502 a_n55_n517# sky130_fd_sc_hd__xor2_1_0/VPB 0
C503 sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__or4_1_0/C 0.00406f
C504 sky130_fd_sc_hd__and2_1_0/VPB sky130_fd_sc_hd__and2_1_0/A 0.00109f
C505 a_n55_n517# B 0.04704f
C506 sky130_fd_sc_hd__and4_1_1/A sky130_fd_sc_hd__and4_1_1/VPWR -0.00839f
C507 a_n53_n3749# A 0.03479f
C508 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__and2_1_4/VPB 0.00887f
C509 a_n55_n517# a_67_n1483# 0.00144f
C510 sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__or2_1_0/A 0.03627f
C511 a_195_n767# A 0.0022f
C512 X sky130_fd_sc_hd__and3_1_0/a_27_47# 0.17069f
C513 sky130_fd_sc_hd__and3_1_0/VPB X 0.0389f
C514 B sky130_fd_sc_hd__and2_1_4/VPWR 0
C515 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__or2_1_0/A 0.00152f
C516 sky130_fd_sc_hd__and4_1_0/B VPB 0.01097f
C517 X sky130_fd_sc_hd__and2_1_5/a_145_75# 0.00203f
C518 sky130_fd_sc_hd__or4_1_0/VPWR sky130_fd_sc_hd__or4_1_0/a_205_297# -0
C519 sky130_fd_sc_hd__and4_1_1/a_197_47# sky130_fd_sc_hd__and4_1_1/VGND -0
C520 sky130_fd_sc_hd__and2_1_5/a_59_75# sky130_fd_sc_hd__and2_1_5/VGND -0.00121f
C521 a_195_n517# sky130_fd_sc_hd__and4_1_0/B 0.00425f
C522 sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__or4_1_0/VGND 0.00186f
C523 a_29_n3749# B 0.00416f
C524 a_59_n3151# B 0.05725f
C525 sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__or4_1_0/B 0
C526 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__or4_1_0/VGND -0.00228f
C527 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__or2_1_0/VGND 0.00393f
C528 sky130_fd_sc_hd__xor2_1_0/VPB sky130_fd_sc_hd__and2_1_0/A 0
C529 sky130_fd_sc_hd__or2_1_0/a_68_297# sky130_fd_sc_hd__and4_1_1/VGND 0
C530 a_59_n3151# a_67_n1483# 0
C531 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__and3_1_0/VGND 0
C532 sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__and4_1_0/VGND 0.00665f
C533 sky130_fd_sc_hd__and4_1_1/A sky130_fd_sc_hd__and4_1_1/VPB 0
C534 B sky130_fd_sc_hd__and2_1_0/A 0.13596f
C535 A sky130_fd_sc_hd__and3_1_0/VGND 0.00212f
C536 X sky130_fd_sc_hd__xor2_1_0/X 0.79943f
C537 sky130_fd_sc_hd__and4_1_0/VGND sky130_fd_sc_hd__and2_1_4/VPB 0
C538 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__or4_1_0/A 0
C539 a_67_n1483# sky130_fd_sc_hd__and2_1_0/A 0
C540 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and2_1_0/a_59_75# 0.01295f
C541 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and2_1_5/VGND 0.00461f
C542 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and4_1_1/C 0.1163f
C543 sky130_fd_sc_hd__and4_1_0/a_303_47# A 0
C544 sky130_fd_sc_hd__and4_1_1/a_109_47# sky130_fd_sc_hd__and4_1_1/VPWR -0
C545 X sky130_fd_sc_hd__or4_1_0/VPB 0
C546 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and4_1_1/a_303_47# 0.00124f
C547 sky130_fd_sc_hd__or2_1_0/VPB sky130_fd_sc_hd__or2_1_0/VPWR -0.00808f
C548 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and4_1_0/a_109_47# 0
C549 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and4_1_0/a_197_47# 0.00195f
C550 sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__or2_1_0/A 0.00385f
C551 sky130_fd_sc_hd__or4_1_0/D sky130_fd_sc_hd__or2_1_0/VPB 0.00363f
C552 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__or2_1_0/VPWR 0
C553 sky130_fd_sc_hd__or4_1_0/VGND sky130_fd_sc_hd__or2_1_0/A 0.00398f
C554 sky130_fd_sc_hd__and2_1_0/B sky130_fd_sc_hd__xor2_1_0/B 0.00243f
C555 X sky130_fd_sc_hd__or2_1_0/a_150_297# 0
C556 sky130_fd_sc_hd__and3_1_0/VPWR sky130_fd_sc_hd__and3_1_0/a_181_47# -0
C557 sky130_fd_sc_hd__and3_1_0/a_27_47# VPB 0
C558 a_155_n4715# A 0.00154f
C559 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__and2_1_4/a_59_75# 0.00834f
C560 sky130_fd_sc_hd__or4_1_0/A sky130_fd_sc_hd__or2_1_0/a_68_297# 0.00411f
C561 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__or4_1_0/D 0
C562 A sky130_fd_sc_hd__and2_1_0/B 0
C563 A sky130_fd_sc_hd__and2_1_4/a_59_75# 0
C564 X a_153_n1483# 0.0017f
C565 a_n55_n517# sky130_fd_sc_hd__xor2_1_0/B 0
C566 sky130_fd_sc_hd__and4_1_0/a_303_47# sky130_fd_sc_hd__and4_1_0/VGND -0
C567 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__or4_1_0/VPWR -0.00317f
C568 X sky130_fd_sc_hd__and4_1_1/a_27_47# 0.04852f
C569 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and4_1_1/a_27_47# 0.03795f
C570 sky130_fd_sc_hd__and2_1_5/VPB B 0
C571 a_n55_n517# A 0.03423f
C572 sky130_fd_sc_hd__and2_1_4/VGND sky130_fd_sc_hd__and2_1_4/VPB -0.00451f
C573 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__and2_1_4/VPWR 0.01674f
C574 sky130_fd_sc_hd__and3_1_0/VPWR a_n63_n2185# 0
C575 sky130_fd_sc_hd__or2_1_0/VPWR sky130_fd_sc_hd__or2_1_0/A 0.15486f
C576 X sky130_fd_sc_hd__and2_1_0/a_145_75# 0
C577 X sky130_fd_sc_hd__and3_1_0/a_109_47# 0.0025f
C578 sky130_fd_sc_hd__or4_1_0/A sky130_fd_sc_hd__and3_1_0/a_27_47# 0
C579 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__or4_1_0/a_109_297# 0
C580 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__or4_1_0/a_27_297# 0.03318f
C581 sky130_fd_sc_hd__and2_1_0/VPB sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.0035f
C582 sky130_fd_sc_hd__xor2_1_0/X VPB 0
C583 sky130_fd_sc_hd__or4_1_0/D sky130_fd_sc_hd__or2_1_0/A 0.00187f
C584 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and4_1_1/VGND 0.04307f
C585 sky130_fd_sc_hd__or4_1_0/X sky130_fd_sc_hd__or4_1_0/A 0.00747f
C586 sky130_fd_sc_hd__or4_1_0/VPWR sky130_fd_sc_hd__or4_1_0/a_277_297# -0
C587 sky130_fd_sc_hd__and4_1_1/a_303_47# sky130_fd_sc_hd__and4_1_1/VGND -0
C588 sky130_fd_sc_hd__and4_1_1/VPB sky130_fd_sc_hd__and4_1_1/VPWR -0.0058f
C589 sky130_fd_sc_hd__and2_1_0/B sky130_fd_sc_hd__xor2_1_0/a_285_297# 0
C590 a_195_n767# sky130_fd_sc_hd__and4_1_0/B 0
C591 sky130_fd_sc_hd__and2_1_4/a_59_75# sky130_fd_sc_hd__and4_1_0/VGND 0
C592 a_59_n3151# sky130_fd_sc_hd__or4_1_0/C 0
C593 sky130_fd_sc_hd__and3_1_0/VPWR sky130_fd_sc_hd__and4_1_0/a_27_47# 0
C594 sky130_fd_sc_hd__or2_1_0/VPWR sky130_fd_sc_hd__or4_1_0/VGND 0
C595 a_197_n3749# B 0.00778f
C596 a_29_n3749# A -0
C597 X sky130_fd_sc_hd__and2_1_4/a_145_75# 0.00133f
C598 a_59_n3151# A 0.02803f
C599 sky130_fd_sc_hd__and4_1_0/VPB sky130_fd_sc_hd__or4_1_0/D 0
C600 sky130_fd_sc_hd__or4_1_0/D sky130_fd_sc_hd__or4_1_0/VGND -0
C601 sky130_fd_sc_hd__and4_1_1/A X 0.09388f
C602 sky130_fd_sc_hd__and4_1_1/A sky130_fd_sc_hd__and4_1_1/C 0.04301f
C603 sky130_fd_sc_hd__xor2_1_0/B sky130_fd_sc_hd__and2_1_0/A 0
C604 sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__or2_1_0/a_68_297# 0.00803f
C605 B sky130_fd_sc_hd__or2_1_0/A 0
C606 A sky130_fd_sc_hd__and2_1_0/A 0.00268f
C607 sky130_fd_sc_hd__and4_1_0/VGND sky130_fd_sc_hd__and2_1_4/VPWR 0
C608 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__or4_1_0/A 0
C609 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and2_1_0/a_59_75# 0
C610 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and2_1_5/VGND 0.11264f
C611 sky130_fd_sc_hd__and4_1_0/VPB B 0
C612 sky130_fd_sc_hd__and4_1_1/a_27_47# sky130_fd_sc_hd__and4_1_1/VGND -0.014f
C613 sky130_fd_sc_hd__or4_1_0/VPB sky130_fd_sc_hd__or4_1_0/A 0.01499f
C614 sky130_fd_sc_hd__xor2_1_0/X sky130_fd_sc_hd__and4_1_0/a_197_47# 0.00123f
C615 sky130_fd_sc_hd__and4_1_0/VPWR sky130_fd_sc_hd__and4_1_0/a_27_47# -0
C616 sky130_fd_sc_hd__and4_1_0/VPB a_67_n1483# 0
C617 B sky130_fd_sc_hd__xor2_1_0/a_35_297# 0
C618 sky130_fd_sc_hd__and4_1_0/a_303_47# sky130_fd_sc_hd__and4_1_0/B 0
C619 sky130_fd_sc_hd__or4_1_0/D sky130_fd_sc_hd__or2_1_0/VPWR 0.00421f
C620 B a_187_n2435# 0
C621 sky130_fd_sc_hd__or2_1_0/B sky130_fd_sc_hd__and3_1_0/a_27_47# 0.00879f
C622 a_n55_n517# sky130_fd_sc_hd__and2_1_5/a_59_75# 0
C623 sky130_fd_sc_hd__or2_1_0/VGND sky130_fd_sc_hd__or2_1_0/a_68_297# -0.00129f
C624 sky130_fd_sc_hd__and3_1_0/VPB sky130_fd_sc_hd__or2_1_0/B 0.01095f
C625 sky130_fd_sc_hd__or4_1_0/a_205_297# sky130_fd_sc_hd__or4_1_0/VGND -0
C626 sky130_fd_sc_hd__and2_1_4/VGND sky130_fd_sc_hd__and2_1_4/a_59_75# -0
C627 sky130_fd_sc_hd__and2_1_0/VPB B 0.00364f
C628 X a_69_n4715# 0
C629 sky130_fd_sc_hd__and3_1_0/a_27_47# sky130_fd_sc_hd__and2_1_4/VPB 0
C630 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__or2_1_0/VPB 0.00444f
C631 sky130_fd_sc_hd__and4_1_0/B sky130_fd_sc_hd__and2_1_0/B 0.02591f
C632 sky130_fd_sc_hd__and2_1_5/VPB sky130_fd_sc_hd__and2_1_5/VPWR -0.00635f
C633 sky130_fd_sc_hd__or4_1_0/C sky130_fd_sc_hd__or4_1_0/B 0.00771f
C634 X sky130_fd_sc_hd__and4_1_1/a_109_47# 0
C635 sky130_fd_sc_hd__or4_1_0/A sky130_fd_sc_hd__and4_1_1/a_27_47# 0
C636 sky130_fd_sc_hd__and4_1_1/C sky130_fd_sc_hd__and4_1_1/a_109_47# 0.0023f
C637 sky130_fd_sc_hd__or4_1_0/B sky130_fd_sc_hd__and2_1_5/VPWR 0
C638 sky130_fd_sc_hd__and4_1_1/A sky130_fd_sc_hd__and4_1_1/VGND -0.007f
C639 sky130_fd_sc_hd__and2_1_4/VGND sky130_fd_sc_hd__and2_1_4/VPWR -0.02765f
C640 a_69_n4715# VNB 0.1752f
C641 a_n53_n3749# VNB 0.24712f
C642 a_59_n3151# VNB 0.17114f
C643 a_n63_n2185# VNB 0.24424f
C644 a_67_n1483# VNB 0.17003f
C645 a_n55_n517# VNB 0.24496f
C646 a_197_n3749# VNB 0.00137f
C647 a_195_n517# VNB 0.00137f
C648 sky130_fd_sc_hd__xor2_1_0/A VNB 0.45606f
C649 sky130_fd_sc_hd__xor2_1_0/B VNB 0.59565f
C650 sky130_fd_sc_hd__xor2_1_0/VPB VNB 0.69336f
C651 sky130_fd_sc_hd__xor2_1_0/a_285_297# VNB 0.00137f
C652 sky130_fd_sc_hd__xor2_1_0/a_35_297# VNB 0.25457f
C653 sky130_fd_sc_hd__and3_1_0/VGND VNB 0.30013f
C654 sky130_fd_sc_hd__or2_1_0/B VNB 0.46058f
C655 sky130_fd_sc_hd__and3_1_0/VPWR VNB 0.27425f
C656 sky130_fd_sc_hd__and3_1_0/VPB VNB 0.51617f
C657 sky130_fd_sc_hd__and3_1_0/a_27_47# VNB 0.17719f
C658 sky130_fd_sc_hd__or4_1_0/VGND VNB 0.36697f
C659 sky130_fd_sc_hd__or4_1_0/X VNB 0.08835f
C660 sky130_fd_sc_hd__or4_1_0/D VNB 0.17526f
C661 sky130_fd_sc_hd__or4_1_0/B VNB 0.799f
C662 sky130_fd_sc_hd__or4_1_0/VPWR VNB 0.28998f
C663 sky130_fd_sc_hd__or4_1_0/VPB VNB 0.60476f
C664 sky130_fd_sc_hd__or4_1_0/a_27_297# VNB 0.16291f
C665 sky130_fd_sc_hd__and4_1_1/VGND VNB 0.39291f
C666 sky130_fd_sc_hd__and4_1_1/VPWR VNB 0.33454f
C667 sky130_fd_sc_hd__and4_1_1/A VNB 0.23645f
C668 sky130_fd_sc_hd__and4_1_1/VPB VNB 0.69336f
C669 sky130_fd_sc_hd__and4_1_1/a_27_47# VNB 0.17489f
C670 sky130_fd_sc_hd__and4_1_0/VGND VNB 0.39291f
C671 sky130_fd_sc_hd__or2_1_0/A VNB 0.31965f
C672 sky130_fd_sc_hd__and4_1_0/VPWR VNB 0.33454f
C673 sky130_fd_sc_hd__xor2_1_0/X VNB 1.89098f
C674 sky130_fd_sc_hd__and4_1_0/B VNB 0.74819f
C675 sky130_fd_sc_hd__and4_1_0/VPB VNB 0.69336f
C676 sky130_fd_sc_hd__and4_1_0/a_27_47# VNB 0.17489f
C677 sky130_fd_sc_hd__or2_1_0/VGND VNB 0.32043f
C678 sky130_fd_sc_hd__or4_1_0/A VNB 0.42983f
C679 sky130_fd_sc_hd__or2_1_0/VPWR VNB 0.26856f
C680 sky130_fd_sc_hd__or2_1_0/VPB VNB 0.51617f
C681 sky130_fd_sc_hd__or2_1_0/a_68_297# VNB 0.15387f
C682 sky130_fd_sc_hd__and2_1_5/VGND VNB 0.3114f
C683 sky130_fd_sc_hd__and4_1_1/C VNB 0.33836f
C684 sky130_fd_sc_hd__and2_1_5/VPWR VNB 0.27345f
C685 sky130_fd_sc_hd__and2_1_5/VPB VNB 0.51617f
C686 sky130_fd_sc_hd__and2_1_5/a_59_75# VNB 0.17706f
C687 sky130_fd_sc_hd__and2_1_4/VGND VNB 0.3114f
C688 sky130_fd_sc_hd__or4_1_0/C VNB 1.43825f
C689 sky130_fd_sc_hd__and2_1_4/VPWR VNB 0.27345f
C690 sky130_fd_sc_hd__and2_1_4/VPB VNB 0.51617f
C691 sky130_fd_sc_hd__and2_1_4/a_59_75# VNB 0.17706f
C692 X VNB 5.38747f
C693 A VNB 2.72305f
C694 B VNB 2.14424f
C695 VPB VNB 3.62859f
C696 sky130_fd_sc_hd__and2_1_0/B VNB 0.2887f
C697 sky130_fd_sc_hd__and2_1_0/A VNB 0.39407f
C698 sky130_fd_sc_hd__and2_1_0/VPB VNB 0.51617f
C699 sky130_fd_sc_hd__and2_1_0/a_59_75# VNB 0.17706f
C700 a_187_n2185# VNB 0.00137f
.ends

.subckt sky130_fd_sc_hd__fa_1 A B CIN VGND VNB VPB VPWR COUT SUM a_1163_413# a_738_413#
+ a_1163_47# a_208_47# a_382_413# a_738_47# a_995_47# a_1091_47# a_76_199# a_1091_413#
+ a_382_47# a_208_413#
X0 a_76_199# B a_208_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X1 VGND A a_382_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_738_413# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_1091_47# CIN a_995_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 VPWR CIN a_738_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 a_382_413# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_1163_47# B a_1091_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X7 VPWR A a_382_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_995_47# a_76_199# a_738_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X9 a_382_413# CIN a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 SUM a_995_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10235 ps=0.995 w=0.65 l=0.15
X11 a_208_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.10235 ps=0.995 w=0.42 l=0.15
X12 VGND CIN a_738_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 a_76_199# B a_208_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.063 ps=0.72 w=0.42 l=0.15
X14 a_208_413# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.14785 ps=1.345 w=0.42 l=0.15
X15 a_738_413# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X16 VGND A a_1163_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10235 pd=0.995 as=0.0693 ps=0.75 w=0.42 l=0.15
X17 a_738_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X18 a_738_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06195 pd=0.715 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 a_1163_413# B a_1091_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X20 VPWR A a_1163_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14785 pd=1.345 as=0.0693 ps=0.75 w=0.42 l=0.15
X21 a_382_47# CIN a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X22 a_382_47# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X23 SUM a_995_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14785 ps=1.345 w=1 l=0.15
X24 a_995_47# a_76_199# a_738_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.06195 ps=0.715 w=0.42 l=0.15
X25 VPWR a_76_199# COUT VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14785 pd=1.345 as=0.26 ps=2.52 w=1 l=0.15
X26 a_1091_413# CIN a_995_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X27 VGND a_76_199# COUT VNB sky130_fd_pr__nfet_01v8 ad=0.10235 pd=0.995 as=0.169 ps=1.82 w=0.65 l=0.15
C0 a_995_47# VPB 0.05213f
C1 a_382_413# VPB 0.01154f
C2 a_738_47# a_1163_47# 0
C3 VPWR B 0.25287f
C4 SUM B 0.00111f
C5 a_738_413# a_1163_413# 0
C6 VPWR A 0.0705f
C7 A SUM 0.0054f
C8 a_208_47# VGND 0.00161f
C9 a_382_47# a_738_47# 0.00847f
C10 a_738_47# B 0.00556f
C11 a_1091_47# B 0
C12 A a_738_47# 0.04461f
C13 a_1091_47# A 0
C14 VGND a_1163_47# 0.00175f
C15 COUT VGND 0.05567f
C16 a_738_413# CIN 0.07973f
C17 a_382_47# VGND 0.14174f
C18 VGND B 0.0456f
C19 A VGND 0.10267f
C20 a_738_413# a_1091_413# 0
C21 a_76_199# a_995_47# 0.04882f
C22 a_76_199# VPB 0.10454f
C23 a_382_413# a_76_199# 0.03016f
C24 VPWR a_995_47# 0.21287f
C25 VPWR VPB 0.15613f
C26 SUM a_995_47# 0.1439f
C27 SUM VPB 0.01793f
C28 a_382_413# VPWR 0.15069f
C29 a_1163_413# B 0
C30 A a_1163_413# 0
C31 a_738_47# a_995_47# 0.02301f
C32 a_738_47# VPB 0
C33 a_1091_47# a_995_47# 0.00559f
C34 a_208_413# a_76_199# 0.00682f
C35 a_382_47# CIN 0.03325f
C36 a_208_413# VPWR 0
C37 CIN B 0.61202f
C38 A CIN 0.45517f
C39 a_995_47# VGND 0.19875f
C40 VGND VPB 0.00519f
C41 a_1091_413# B 0
C42 VPWR a_76_199# 0.19016f
C43 a_76_199# SUM 0
C44 a_1163_413# a_995_47# 0.00758f
C45 VPWR SUM 0.07457f
C46 a_76_199# a_738_47# 0.03622f
C47 a_1091_47# a_76_199# 0
C48 a_738_413# B 0.0177f
C49 a_738_413# A 0.01182f
C50 COUT a_208_47# 0
C51 a_995_47# CIN 0.05108f
C52 CIN VPB 0.23153f
C53 a_382_413# CIN 0.08907f
C54 a_76_199# VGND 0.41492f
C55 a_1091_47# a_738_47# 0
C56 VPWR VGND 0.04263f
C57 a_995_47# a_1091_413# 0.00487f
C58 SUM VGND 0.07127f
C59 a_208_47# A 0
C60 B a_1163_47# 0
C61 A a_1163_47# 0
C62 COUT B 0
C63 a_738_47# VGND 0.14671f
C64 COUT A 0.00345f
C65 a_1091_47# VGND 0
C66 VPWR a_1163_413# 0
C67 a_382_47# B 0.01781f
C68 a_382_47# A 0.04028f
C69 a_738_413# VPB 0.01092f
C70 a_738_413# a_995_47# 0.02283f
C71 a_382_413# a_738_413# 0.00985f
C72 A B 0.77269f
C73 a_76_199# CIN 0.21032f
C74 VPWR CIN 0.0577f
C75 a_76_199# a_1091_413# 0
C76 VPWR a_1091_413# 0
C77 a_738_47# CIN 0.04534f
C78 a_995_47# a_1163_47# 0.00792f
C79 COUT VPB 0.01094f
C80 a_738_413# a_76_199# 0.00386f
C81 a_382_47# VPB 0.00139f
C82 VGND CIN 0.06042f
C83 B VPB 0.33717f
C84 a_995_47# B 0.08206f
C85 a_382_413# B 0.03303f
C86 A a_995_47# 0.16271f
C87 A VPB 0.27513f
C88 a_382_413# A 0.01121f
C89 a_738_413# VPWR 0.14479f
C90 a_76_199# a_208_47# 0.00696f
C91 a_208_413# A 0
C92 COUT a_76_199# 0.12975f
C93 SUM a_1163_47# 0
C94 COUT VPWR 0.06663f
C95 a_382_47# a_76_199# 0.06611f
C96 a_76_199# B 0.13093f
C97 a_76_199# A 0.73176f
C98 SUM VNB 0.10031f
C99 VGND VNB 0.81236f
C100 VPWR VNB 0.66922f
C101 COUT VNB 0.09411f
C102 CIN VNB 0.32537f
C103 B VNB 0.47131f
C104 A VNB 0.49582f
C105 VPB VNB 1.49072f
C106 a_738_47# VNB 0.01584f
C107 a_382_47# VNB 0.01578f
C108 a_738_413# VNB 0.00484f
C109 a_382_413# VNB 0.00345f
C110 a_995_47# VNB 0.1359f
C111 a_76_199# VNB 0.2795f
.ends

.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X a_505_21# a_535_374# a_439_47#
+ a_218_47# a_76_199# a_218_374#
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
C0 VGND VPB 0.01345f
C1 S A0 0.03411f
C2 a_439_47# A0 0.00369f
C3 VPWR a_535_374# 0
C4 a_505_21# S 0.19751f
C5 S VPWR 0.39244f
C6 a_439_47# VPWR 0
C7 VGND X 0.05864f
C8 a_76_199# A0 0.05444f
C9 X a_218_47# 0
C10 S VPB 0.16849f
C11 A1 VGND 0.07521f
C12 VPWR a_76_199# 0.05421f
C13 a_218_374# VGND 0
C14 VPB a_76_199# 0.04809f
C15 S X 0.00823f
C16 VGND a_218_47# 0.00328f
C17 A1 S 0.08722f
C18 a_439_47# A1 0.00498f
C19 a_505_21# A0 0.03829f
C20 X a_76_199# 0.07764f
C21 VGND a_535_374# 0
C22 VPWR A0 0.00732f
C23 S VGND 0.03296f
C24 a_439_47# VGND 0.00354f
C25 a_505_21# VPWR 0.08183f
C26 a_218_374# S 0.00688f
C27 A1 a_76_199# 0.18667f
C28 VPB A0 0.1066f
C29 a_505_21# VPB 0.07806f
C30 VGND a_76_199# 0.16013f
C31 VPB VPWR 0.10994f
C32 a_218_374# a_76_199# 0.00557f
C33 a_218_47# a_76_199# 0.00783f
C34 S a_535_374# 0.00526f
C35 X VPWR 0.12783f
C36 a_535_374# a_76_199# 0
C37 A1 A0 0.2668f
C38 S a_76_199# 0.31816f
C39 a_505_21# A1 0.09927f
C40 A1 VPWR 0.01137f
C41 VGND A0 0.04323f
C42 VPB X 0.01205f
C43 a_505_21# VGND 0.12387f
C44 VGND VPWR 0.08036f
C45 A1 VPB 0.07208f
C46 a_218_374# VPWR 0.00177f
C47 a_218_47# VPWR 0
C48 VGND VNB 0.49866f
C49 A1 VNB 0.14042f
C50 A0 VNB 0.13429f
C51 S VNB 0.26814f
C52 VPWR VNB 0.41925f
C53 X VNB 0.09236f
C54 VPB VNB 0.87055f
C55 a_505_21# VNB 0.24676f
C56 a_76_199# VNB 0.13947f
.ends

.subckt tt_um_ohmy90_adders clk ena rst_n ua[0] ua[1] ua[2] ua[3] VGND ua[5] ua[6]
+ ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0]
+ uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0]
+ uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0]
+ uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0]
+ uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
Xsky130_fd_sc_hd__inv_1_4 sky130_fd_sc_hd__inv_1_4/A VGND VNB sky130_fd_sc_hd__inv_1_4/VPB
+ VGND sky130_fd_sc_hd__inv_1_5/A sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_5 sky130_fd_sc_hd__inv_1_5/A VGND VNB sky130_fd_sc_hd__inv_1_5/VPB
+ VGND sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__mux4_1_0 sky130_fd_sc_hd__inv_1_5/Y VGND VGND VGND ui_in[1] ui_in[0]
+ VGND VNB sky130_fd_sc_hd__mux4_1_0/VPB VGND ua[0] sky130_fd_sc_hd__mux4_1_0/a_1290_413#
+ sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__mux4_1_0/a_1478_413# ui_in[0]
+ sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__mux4_1_0/a_923_363#
+ sky130_fd_sc_hd__mux4_1_0/a_193_47# sky130_fd_sc_hd__mux4_1_0/a_834_97# sky130_fd_sc_hd__mux4_1_0/a_247_21#
+ sky130_fd_sc_hd__mux4_1_0/a_668_97# sky130_fd_sc_hd__mux4_1_0/a_193_413# sky130_fd_sc_hd__mux4_1_0/a_27_47#
+ sky130_fd_sc_hd__mux4_1
XCLA_0 VNB CLA_0/sky130_fd_sc_hd__and4_1_1/a_303_47# CLA_0/sky130_fd_sc_hd__and4_1_0/VPB
+ CLA_0/sky130_fd_sc_hd__xor2_1_0/VPB CLA_0/sky130_fd_sc_hd__and2_1_5/VPB CLA_0/a_187_n2185#
+ CLA_0/sky130_fd_sc_hd__and4_1_0/a_27_47# CLA_0/X CLA_0/sky130_fd_sc_hd__or2_1_0/a_150_297#
+ CLA_0/sky130_fd_sc_hd__and2_1_5/a_59_75# VGND CLA_0/sky130_fd_sc_hd__and3_1_0/a_109_47#
+ VGND CLA_0/sky130_fd_sc_hd__and3_1_0/a_181_47# CLA_0/sky130_fd_sc_hd__xor2_1_0/a_285_297#
+ VGND CLA_0/sky130_fd_sc_hd__or4_1_0/B CLA_0/sky130_fd_sc_hd__or4_1_0/a_109_297#
+ VGND VGND CLA_0/sky130_fd_sc_hd__or2_1_0/VPB CLA_0/sky130_fd_sc_hd__and3_1_0/a_27_47#
+ CLA_0/a_187_n2435# VGND CLA_0/sky130_fd_sc_hd__and4_1_1/VPB CLA_0/sky130_fd_sc_hd__xor2_1_0/a_285_47#
+ CLA_0/a_19_n2185# CLA_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# CLA_0/sky130_fd_sc_hd__and2_1_4/a_145_75#
+ CLA_0/sky130_fd_sc_hd__and2_1_0/a_145_75# CLA_0/sky130_fd_sc_hd__and4_1_1/a_27_47#
+ CLA_0/a_155_n4715# VGND CLA_0/sky130_fd_sc_hd__or4_1_0/A VGND CLA_0/sky130_fd_sc_hd__or2_1_0/a_68_297#
+ CLA_0/sky130_fd_sc_hd__and2_1_0/VPB CLA_0/a_195_n517# CLA_0/a_n63_n2185# CLA_0/a_197_n3749#
+ VGND CLA_0/sky130_fd_sc_hd__and4_1_0/a_109_47# CLA_0/a_195_n767# CLA_0/a_197_n3999#
+ VGND VGND VGND CLA_0/sky130_fd_sc_hd__and4_1_0/B CLA_0/sky130_fd_sc_hd__and2_1_5/a_145_75#
+ CLA_0/sky130_fd_sc_hd__and2_1_0/a_59_75# VGND CLA_0/a_153_n1483# CLA_0/a_27_n517#
+ CLA_0/a_69_n4715# CLA_0/sky130_fd_sc_hd__or2_1_0/B CLA_0/sky130_fd_sc_hd__or2_1_0/A
+ CLA_0/sky130_fd_sc_hd__or4_1_0/a_277_297# CLA_0/sky130_fd_sc_hd__and4_1_0/a_197_47#
+ CLA_0/sky130_fd_sc_hd__and2_1_4/VPB CLA_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# CLA_0/sky130_fd_sc_hd__and3_1_0/VPB
+ CLA_0/sky130_fd_sc_hd__and4_1_0/a_303_47# CLA_0/sky130_fd_sc_hd__and4_1_1/C CLA_0/sky130_fd_sc_hd__and4_1_1/a_109_47#
+ CLA_0/sky130_fd_sc_hd__or4_1_0/VPB CLA_0/sky130_fd_sc_hd__or4_1_0/a_27_297# CLA_0/a_29_n3749#
+ VGND CLA_0/sky130_fd_sc_hd__or4_1_0/a_205_297# CLA_0/sky130_fd_sc_hd__and2_1_4/a_59_75#
+ VGND CLA_0/a_n53_n3749# CLA_0/a_n55_n517# sky130_fd_sc_hd__inv_1_2/Y VGND VGND VGND
+ CLA_0/sky130_fd_sc_hd__or4_1_0/C CLA_0/a_67_n1483# VGND CLA_0/a_59_n3151# CLA_0/sky130_fd_sc_hd__xor2_1_0/X
+ CLA_0/sky130_fd_sc_hd__and4_1_1/a_197_47# CLA_0/VPB CLA_0/X VGND CLA_0/a_145_n3151#
+ VGND CLA
XCLA_1 VNB a_11873_15219# VPB VPB VPB a_9717_13091# a_11321_14203# VGND a_11906_13629#
+ a_11019_15169# VGND a_11019_12911# VGND a_11091_12911# a_9715_16323# VGND VGND a_12713_13987#
+ VGND VGND VPB a_11261_13361# a_9717_12841# VGND VPB a_9715_16073# a_9549_13091#
+ a_9957_16523# a_11051_11919# a_9673_15357# a_12105_15669# a_9685_10561# VGND VGND
+ VGND a_12045_13829# VPB a_9725_14759# a_9959_13291# a_9727_11527# VGND a_10895_13753#
+ a_9725_14509# a_9727_11277# VGND VGND VGND VGND a_10857_14747# a_9835_15779# VGND
+ a_9683_13793# a_9557_14759# a_9847_10983# VGND VGND a_12881_13987# a_10983_13753#
+ VPB a_9547_16323# VPB a_11089_13753# VGND a_11679_15219# VPB a_13045_14187# a_9559_11527#
+ VGND a_12809_13987# a_11213_12341# VGND a_9969_11727# a_9967_14959# VGND VGND VGND
+ VGND VGND a_9845_14215# VGND a_9837_12547# VGND a_11767_15219# VPB VGND VGND a_9675_12125#
+ VGND CLA
Xsky130_fd_sc_hd__fa_1_10 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_2079_5051# a_2343_5051#
+ a_2079_5417# a_3040_5417# a_2706_5051# a_2343_5417# a_1950_5501# a_2175_5417# a_3199_5501#
+ a_2175_5051# a_2706_5417# a_3040_5051# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_0 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_2049_1791# a_2313_1791#
+ a_2049_2157# a_3010_2157# a_2676_1791# a_2313_2157# a_1920_2241# a_2145_2157# a_3169_2241#
+ a_2145_1791# a_2676_2157# a_3010_1791# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_11 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_3949_5047# a_4213_5047#
+ a_3949_5413# a_4910_5413# a_4576_5047# a_4213_5413# a_3820_5497# a_4045_5413# a_5069_5497#
+ a_4045_5047# a_4576_5413# a_4910_5047# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_1 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_3919_1787# a_4183_1787#
+ a_3919_2153# a_4880_2153# a_4546_1787# a_4183_2153# a_3790_2237# a_4015_2153# a_5039_2237#
+ a_4015_1787# a_4546_2153# a_4880_1787# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_12 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_11331_5467#
+ a_11595_5467# a_11331_5833# a_12292_5833# a_11958_5467# a_11595_5833# a_11202_5917#
+ a_11427_5833# a_12451_5917# a_11427_5467# a_11958_5833# a_12292_5467# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_3 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_7605_1779# a_7869_1779#
+ a_7605_2145# a_8566_2145# a_8232_1779# a_7869_2145# a_7476_2229# a_7701_2145# a_8725_2229#
+ a_7701_1779# a_8232_2145# a_8566_1779# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_2 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_5735_1783# a_5999_1783#
+ a_5735_2149# a_6696_2149# a_6362_1783# a_5999_2149# a_5606_2233# a_5831_2149# a_6855_2233#
+ a_5831_1783# a_6362_2149# a_6696_1783# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_4 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_14975_1765# a_15239_1765#
+ a_14975_2131# a_15936_2131# a_15602_1765# a_15239_2131# a_14846_2215# a_15071_2131#
+ a_16095_2215# a_15071_1765# a_15602_2131# a_15936_1765# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_13 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_9461_5471# a_9725_5471#
+ a_9461_5837# a_10422_5837# a_10088_5471# a_9725_5837# a_9332_5921# a_9557_5837#
+ a_9695_5921# a_9557_5471# a_10088_5837# a_10422_5471# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_15 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_15017_5459#
+ a_15281_5459# a_15017_5825# a_15978_5825# a_15644_5459# a_15281_5825# a_14888_5909#
+ a_15113_5825# a_16137_5909# a_15113_5459# a_15644_5825# a_15978_5459# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_14 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_13147_5463#
+ a_13411_5463# a_13147_5829# a_14108_5829# a_13774_5463# a_13411_5829# a_13018_5913#
+ a_13243_5829# a_14267_5913# a_13243_5463# a_13774_5829# a_14108_5463# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_5 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_13105_1769# a_13369_1769#
+ a_13105_2135# a_14066_2135# a_13732_1769# a_13369_2135# a_12976_2219# a_13201_2135#
+ a_14225_2219# a_13201_1769# a_13732_2135# a_14066_1769# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_16 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_11359_4593#
+ a_11623_4593# a_11359_4959# a_12320_4959# a_11986_4593# a_11623_4959# a_11230_5043#
+ a_11455_4959# a_12479_5043# a_11455_4593# a_11986_4959# a_12320_4593# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_6 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_9419_1777# a_9683_1777#
+ a_9419_2143# a_10380_2143# a_10046_1777# a_9683_2143# a_9290_2227# a_9515_2143#
+ a_9653_2227# a_9515_1777# a_10046_2143# a_10380_1777# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_7 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_11289_1773# a_11553_1773#
+ a_11289_2139# a_12250_2139# a_11916_1773# a_11553_2139# a_11160_2223# a_11385_2139#
+ a_12409_2223# a_11385_1773# a_11916_2139# a_12250_1773# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_17 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_9489_4597# a_9753_4597#
+ a_9489_4963# a_10450_4963# a_10116_4597# a_9753_4963# a_9360_5047# a_9585_4963#
+ a_9723_5047# a_9585_4597# a_10116_4963# a_10450_4597# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__mux2_1_0 VGND VGND VGND VGND VNB sky130_fd_sc_hd__mux2_1_0/VPB VGND
+ VGND sky130_fd_sc_hd__mux2_1_0/a_505_21# sky130_fd_sc_hd__mux2_1_0/a_535_374# sky130_fd_sc_hd__mux2_1_0/a_439_47#
+ sky130_fd_sc_hd__mux2_1_0/a_218_47# sky130_fd_sc_hd__mux2_1_0/a_76_199# sky130_fd_sc_hd__mux2_1_0/a_218_374#
+ sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__fa_1_18 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_13175_4589#
+ a_13439_4589# a_13175_4955# a_14136_4955# a_13802_4589# a_13439_4955# a_13046_5039#
+ a_13271_4955# a_14295_5039# a_13271_4589# a_13802_4955# a_14136_4589# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__inv_1_1 VGND VGND VNB VPB VGND VGND sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__inv_1_0 VGND VGND VNB sky130_fd_sc_hd__inv_1_0/VPB VGND VGND sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__fa_1_8 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_7635_5039# a_7899_5039#
+ a_7635_5405# a_8596_5405# a_8262_5039# a_7899_5405# a_7506_5489# a_7731_5405# a_8755_5489#
+ a_7731_5039# a_8262_5405# a_8596_5039# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__inv_1_2 VGND VGND VNB sky130_fd_sc_hd__inv_1_2/VPB VGND sky130_fd_sc_hd__inv_1_2/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__fa_1_19 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_15045_4585#
+ a_15309_4585# a_15045_4951# a_16006_4951# a_15672_4585# a_15309_4951# a_14916_5035#
+ a_15141_4951# a_16165_5035# a_15141_4585# a_15672_4951# a_16006_4585# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__fa_1_9 VGND VGND VGND VGND VNB VPB VGND VGND SUM a_5765_5043# a_6029_5043#
+ a_5765_5409# a_6726_5409# a_6392_5043# a_6029_5409# a_5636_5493# a_5861_5409# a_6885_5493#
+ a_5861_5043# a_6392_5409# a_6726_5043# sky130_fd_sc_hd__fa_1
Xsky130_fd_sc_hd__inv_1_3 sky130_fd_sc_hd__inv_1_5/Y VGND VNB sky130_fd_sc_hd__inv_1_3/VPB
+ VGND sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__inv_1
C0 a_4546_1787# VGND 0.02548f
C1 VPB a_3790_2237# 0
C2 a_15045_4951# VGND 0
C3 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__mux4_1_0/a_193_47# 0
C4 sky130_fd_sc_hd__inv_1_0/VPB VGND 0.05044f
C5 a_16095_2215# VPB -0
C6 ua[5] a_11160_2223# 0
C7 CLA_0/sky130_fd_sc_hd__or2_1_0/A VGND 0.13949f
C8 a_6855_2233# VGND 0.09158f
C9 a_6696_2149# VGND 0
C10 a_13147_5463# VGND 0
C11 sky130_fd_sc_hd__mux4_1_0/a_757_363# ui_in[0] -0
C12 CLA_0/sky130_fd_sc_hd__or4_1_0/B CLA_0/X 0.07386f
C13 CLA_0/sky130_fd_sc_hd__and4_1_1/a_109_47# VGND 0
C14 VGND a_10046_2143# 0.00692f
C15 a_7899_5405# VGND 0.01507f
C16 a_13732_2135# VGND 0.00689f
C17 a_9653_2227# a_10046_2143# 0
C18 CLA_0/VPB VGND 0.17645f
C19 ua[4] a_14975_1765# 0
C20 a_11160_2223# VPB 0
C21 a_14916_5035# a_14888_5909# 0
C22 a_14888_5909# a_16137_5909# -0.00146f
C23 a_12881_13987# a_13045_14187# -0
C24 CLA_0/a_195_n517# CLA_0/X -0
C25 a_9673_15357# VGND 0.0031f
C26 a_14888_5909# VPB 0
C27 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0
C28 a_7605_1779# VGND 0
C29 a_8725_2229# VGND 0.08985f
C30 a_3169_2241# a_3790_2237# 0.00446f
C31 CLA_0/sky130_fd_sc_hd__and2_1_5/VPB CLA_0/X -0
C32 CLA_0/a_197_n3999# VGND 0.00312f
C33 sky130_fd_sc_hd__mux4_1_0/a_193_47# VGND 0
C34 a_9845_14215# a_9837_12547# -0
C35 CLA_0/sky130_fd_sc_hd__or4_1_0/a_205_297# CLA_0/X 0
C36 sky130_fd_sc_hd__mux4_1_0/a_668_97# VGND 0.01571f
C37 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__inv_1_5/A 0.05599f
C38 SUM a_6885_5493# -0
C39 a_7605_2145# VGND 0
C40 a_14267_5913# VGND 0.13481f
C41 a_9845_14215# VGND 0.05008f
C42 a_11202_5917# a_11427_5833# -0
C43 VGND a_11427_5467# 0
C44 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_0/a_193_413# -0
C45 CLA_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# CLA_0/sky130_fd_sc_hd__and4_1_0/B -0
C46 CLA_0/sky130_fd_sc_hd__and2_1_5/VPB CLA_0/sky130_fd_sc_hd__and4_1_1/C -0
C47 uo_out[6] uo_out[5] 0.03102f
C48 a_14975_1765# VGND 0
C49 a_9685_10561# VGND 0.00186f
C50 a_8596_5039# VGND 0
C51 a_15239_1765# VGND 0.01595f
C52 a_5861_5043# VGND 0
C53 a_13802_4955# VGND 0.00794f
C54 sky130_fd_sc_hd__inv_1_2/Y VGND 1.61762f
C55 CLA_0/X CLA_0/sky130_fd_sc_hd__or2_1_0/VPB 0
C56 SUM a_5069_5497# -0
C57 a_9835_15779# VPB 0
C58 a_8566_1779# VGND 0
C59 SUM a_9332_5921# 0
C60 a_11230_5043# a_11455_4593# -0
C61 sky130_fd_sc_hd__mux4_1_0/a_1478_413# VGND 0.00234f
C62 SUM ua[5] 0
C63 CLA_0/a_29_n3749# VGND 0.00521f
C64 a_9360_5047# VGND 0.10061f
C65 a_16137_5909# SUM -0
C66 CLA_0/sky130_fd_sc_hd__and2_1_4/a_145_75# VGND 0.00112f
C67 a_11160_2223# a_11289_2139# 0
C68 a_5069_5497# a_3820_5497# -0.00146f
C69 a_9957_16523# a_9967_14959# -0
C70 CLA_0/sky130_fd_sc_hd__xor2_1_0/VPB CLA_0/sky130_fd_sc_hd__and4_1_0/B -0
C71 VGND a_11359_4959# 0
C72 a_15309_4585# VGND 0.0153f
C73 a_10088_5471# VGND 0.02811f
C74 SUM VPB 0.03448f
C75 CLA_0/a_n53_n3749# VGND 0.06201f
C76 ui_in[1] sky130_fd_sc_hd__mux4_1_0/a_1290_413# 0.02507f
C77 ui_in[7] ui_in[6] 0.03102f
C78 uio_out[3] uio_out[2] 0.03102f
C79 uio_in[4] uio_in[3] 0.03102f
C80 a_11019_12911# VGND 0.00147f
C81 a_4880_1787# VGND 0
C82 VPB a_3820_5497# 0
C83 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__mux4_1_0/a_27_413# 0.05016f
C84 a_2676_2157# VGND 0.01205f
C85 a_11261_13361# a_9959_13291# -0
C86 CLA_0/a_n63_n2185# CLA_0/X -0.00179f
C87 uio_oe[5] uio_oe[4] 0.03102f
C88 a_14108_5829# VGND 0
C89 CLA_0/sky130_fd_sc_hd__or4_1_0/a_27_297# CLA_0/X 0.02052f
C90 a_7731_5405# VGND 0.00117f
C91 sky130_fd_sc_hd__inv_1_2/Y CLA_0/sky130_fd_sc_hd__or2_1_0/A 0
C92 VGND a_9683_2143# 0.01374f
C93 a_9653_2227# a_9683_2143# -0
C94 a_13369_2135# VGND 0.01323f
C95 VGND a_3790_2237# 0.10989f
C96 SUM a_3169_2241# -0
C97 a_16095_2215# VGND 0.08521f
C98 a_9969_11727# VPB 0
C99 a_12320_4593# VGND 0
C100 CLA_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0
C101 CLA_0/a_n55_n517# VGND 0.06497f
C102 sky130_fd_sc_hd__inv_1_3/VPB sky130_fd_sc_hd__inv_1_5/Y 0.02733f
C103 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__mux4_1_0/a_27_47# 0.00682f
C104 a_6885_5493# a_7506_5489# 0.00446f
C105 CLA_0/a_69_n4715# VGND 0.03311f
C106 ui_in[0] sky130_fd_sc_hd__mux4_1_0/VPB 0.01835f
C107 a_11160_2223# VGND 0.10935f
C108 a_9653_2227# a_11160_2223# 0.00446f
C109 CLA_0/a_67_n1483# VGND 0.04655f
C110 a_9557_5471# a_9332_5921# -0
C111 sky130_fd_sc_hd__mux4_1_0/a_27_413# VGND -0
C112 a_8725_2229# a_8566_1779# -0
C113 a_14888_5909# VGND 0.12814f
C114 CLA_0/sky130_fd_sc_hd__and4_1_0/VPB CLA_0/sky130_fd_sc_hd__or4_1_0/C -0
C115 a_15936_2131# VGND 0
C116 a_8262_5039# VGND 0.02727f
C117 a_11202_5917# a_9695_5921# 0.00446f
C118 a_9332_5921# a_7506_5489# 0
C119 CLA_0/a_197_n3749# VGND 0.02436f
C120 a_13439_4955# VGND 0.00817f
C121 CLA_0/sky130_fd_sc_hd__and3_1_0/VPB CLA_0/X -0.00135f
C122 a_5765_5043# VGND 0
C123 CLA_0/sky130_fd_sc_hd__or4_1_0/C CLA_0/sky130_fd_sc_hd__and2_1_4/VPB 0
C124 a_11202_5917# a_11595_5467# 0
C125 SUM a_12479_5043# -0
C126 a_11230_5043# a_11359_4593# -0
C127 CLA_0/sky130_fd_sc_hd__and4_1_0/B CLA_0/X -0.02121f
C128 a_5606_2233# a_5039_2237# 0.00492f
C129 VGND a_2175_5051# 0
C130 a_14888_5909# a_15113_5825# -0
C131 sky130_fd_sc_hd__inv_1_3/VPB VGND 0.0254f
C132 sky130_fd_sc_hd__inv_1_5/Y ui_in[0] 0.0136f
C133 VPB a_7506_5489# 0
C134 a_4576_5047# VGND 0.0254f
C135 sky130_fd_sc_hd__mux4_1_0/a_27_47# VGND 0.01764f
C136 a_10088_5837# a_9695_5921# 0
C137 CLA_0/X CLA_0/sky130_fd_sc_hd__or4_1_0/A 0.13855f
C138 a_15141_4585# VGND 0
C139 CLA_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# CLA_0/sky130_fd_sc_hd__and4_1_0/B -0
C140 a_9725_5471# VGND 0.01857f
C141 uio_oe[0] uio_out[7] 0.03102f
C142 a_9957_16523# a_9725_14759# -0
C143 a_9835_15779# VGND 0.05453f
C144 a_9957_16523# VPB 0
C145 a_5606_2233# a_5999_1783# 0
C146 a_11091_12911# VGND 0
C147 ua[0] ui_in[1] 0.36102f
C148 rst_n clk 0.03102f
C149 CLA_0/X CLA_0/sky130_fd_sc_hd__and4_1_0/a_109_47# -0
C150 a_4015_2153# VGND 0.00111f
C151 a_9959_13291# VPB -0
C152 a_13045_14187# a_12713_13987# 0
C153 sky130_fd_sc_hd__mux4_1_0/VPB sky130_fd_sc_hd__mux4_1_0/a_247_21# -0
C154 SUM VGND 1.55293f
C155 a_9559_11527# VGND 0.00521f
C156 SUM a_9653_2227# -0
C157 VGND a_9515_2143# 0.0011f
C158 a_7635_5405# VGND 0
C159 a_13201_2135# VGND 0.0011f
C160 ui_in[0] VGND 0.31308f
C161 a_8755_5489# a_9695_5921# 0
C162 a_9683_13793# VGND 0.00278f
C163 CLA_0/sky130_fd_sc_hd__and4_1_1/a_27_47# CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0.00235f
C164 VGND a_3820_5497# 0.10969f
C165 VGND a_12250_1773# 0
C166 a_11986_4593# VGND 0.0272f
C167 CLA_0/sky130_fd_sc_hd__or4_1_0/B CLA_0/sky130_fd_sc_hd__or4_1_0/A -0
C168 a_16165_5035# a_15672_4951# 0
C169 CLA_0/sky130_fd_sc_hd__and4_1_0/B CLA_0/a_195_n517# -0
C170 ui_in[1] sky130_fd_sc_hd__mux4_1_0/a_750_97# 0.19133f
C171 a_4183_2153# a_5039_2237# -0
C172 a_9547_16323# VGND 0.00465f
C173 a_13018_5913# a_13243_5829# -0
C174 CLA_0/sky130_fd_sc_hd__and4_1_0/VPB VGND 0.02374f
C175 CLA_0/sky130_fd_sc_hd__and3_1_0/a_27_47# CLA_0/X -0.00174f
C176 a_11202_5917# a_11331_5833# 0
C177 CLA_0/sky130_fd_sc_hd__and2_1_5/VPB CLA_0/sky130_fd_sc_hd__and4_1_0/B -0
C178 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.017f
C179 CLA_0/sky130_fd_sc_hd__or4_1_0/C CLA_0/sky130_fd_sc_hd__or2_1_0/a_68_297# -0
C180 a_14888_5909# a_14267_5913# 0.00446f
C181 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__inv_1_4/VPB 0.00994f
C182 CLA_0/sky130_fd_sc_hd__and2_1_4/VPB VGND 0.02145f
C183 a_9969_11727# VGND 0.06157f
C184 CLA_0/X CLA_0/sky130_fd_sc_hd__xor2_1_0/X 0.01329f
C185 VPB a_14225_2219# 0
C186 VGND CLA_0/sky130_fd_sc_hd__and2_1_0/a_145_75# 0.0031f
C187 uo_out[5] uo_out[4] 0.03102f
C188 a_9723_5047# a_9695_5921# 0.00177f
C189 a_15602_2131# VGND 0.00957f
C190 CLA_0/sky130_fd_sc_hd__or4_1_0/VPB CLA_0/X 0.01615f
C191 a_7899_5039# VGND 0.02189f
C192 a_11331_5467# VGND 0
C193 a_9835_15779# a_9673_15357# 0
C194 SUM a_6855_2233# -0
C195 CLA_0/sky130_fd_sc_hd__and3_1_0/a_109_47# CLA_0/X -0
C196 sky130_fd_sc_hd__mux4_1_0/a_834_97# VGND 0.01458f
C197 a_13271_4955# VGND 0.00115f
C198 CLA_0/sky130_fd_sc_hd__xor2_1_0/X CLA_0/sky130_fd_sc_hd__and2_1_0/VPB -0
C199 CLA_0/sky130_fd_sc_hd__and4_1_1/C CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0.00251f
C200 CLA_0/sky130_fd_sc_hd__or4_1_0/a_277_297# VGND 0
C201 a_9290_2227# VPB 0
C202 uo_out[0] uio_in[7] 0.03102f
C203 a_3169_2241# a_2676_1791# 0
C204 CLA_0/sky130_fd_sc_hd__and4_1_0/a_303_47# VGND 0.00141f
C205 a_13045_14187# VPB 0
C206 a_6362_2149# VGND 0.00706f
C207 a_4910_5413# VGND 0
C208 a_11230_5043# a_11202_5917# 0
C209 a_2145_2157# VGND 0.00147f
C210 CLA_0/X a_9967_14959# 0
C211 a_9360_5047# a_8262_5039# 0
C212 ua[0] sky130_fd_sc_hd__mux4_1_0/a_1290_413# 0.00198f
C213 CLA_0/sky130_fd_sc_hd__or2_1_0/VPB CLA_0/sky130_fd_sc_hd__or4_1_0/A -0
C214 a_9725_5837# a_9695_5921# -0
C215 a_9717_12841# VGND 0.00364f
C216 a_9835_15779# a_9845_14215# -0
C217 a_15045_4585# VGND 0
C218 ui_in[1] sky130_fd_sc_hd__mux4_1_0/a_923_363# 0.00109f
C219 VGND sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.05556f
C220 a_9557_5471# VGND 0
C221 sky130_fd_sc_hd__inv_1_4/VPB VGND 0.02147f
C222 SUM a_8725_2229# -0
C223 rst_n ui_in[0] 0.03102f
C224 CLA_0/a_27_n517# VGND 0.00521f
C225 ui_in[6] ui_in[5] 0.03102f
C226 a_15978_5459# VGND 0
C227 a_5606_2233# a_5831_1783# -0
C228 CLA_0/sky130_fd_sc_hd__or4_1_0/B CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0
C229 uio_in[3] uio_in[2] 0.03102f
C230 VGND a_7506_5489# 0.11f
C231 CLA_0/sky130_fd_sc_hd__and4_1_0/a_197_47# VGND 0.00146f
C232 a_14267_5913# SUM -0
C233 a_4576_5413# a_5069_5497# 0
C234 a_13774_5829# VGND 0.00916f
C235 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__mux4_1_0/a_193_413# 0.01304f
C236 sky130_fd_sc_hd__mux4_1_0/a_668_97# ui_in[0] 0
C237 uio_oe[4] uio_oe[3] 0.03102f
C238 a_9957_16523# VGND 0.06504f
C239 VGND a_9419_2143# 0
C240 a_5606_2233# VPB 0
C241 CLA_0/sky130_fd_sc_hd__and2_1_5/VPB CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0
C242 CLA_0/X a_9717_13091# 0
C243 a_13045_14187# a_11321_14203# -0
C244 sky130_fd_sc_hd__mux4_1_0/a_757_363# ui_in[1] 0.03011f
C245 a_9959_13291# VGND 0.0634f
C246 a_10116_4963# a_8755_5489# 0
C247 VGND a_11916_1773# 0.02553f
C248 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__inv_1_5/VPB 0.02677f
C249 VGND CLA_0/sky130_fd_sc_hd__or2_1_0/a_68_297# 0.03248f
C250 CLA_0/sky130_fd_sc_hd__or4_1_0/a_27_297# CLA_0/sky130_fd_sc_hd__or4_1_0/A -0
C251 a_11623_4593# VGND 0.01618f
C252 a_16165_5035# a_15309_4951# -0
C253 ui_in[0] sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.02886f
C254 a_9715_16323# VGND 0.01931f
C255 a_13105_2135# VGND 0
C256 sky130_fd_sc_hd__inv_1_2/Y CLA_0/sky130_fd_sc_hd__and4_1_0/VPB 0
C257 a_2676_1791# VGND 0.03005f
C258 VGND sky130_fd_sc_hd__mux4_1_0/a_193_413# 0.004f
C259 CLA_0/X a_9847_10983# 0
C260 a_15239_2131# VGND 0.00994f
C261 a_7731_5039# VGND 0
C262 a_10116_4963# a_9723_5047# 0
C263 a_14916_5035# a_16165_5035# -0.00146f
C264 CLA_0/sky130_fd_sc_hd__and2_1_4/a_59_75# VGND 0.02988f
C265 a_16165_5035# a_16137_5909# 0.00177f
C266 VGND a_9549_13091# 0.00548f
C267 a_14225_2219# a_12976_2219# -0.00146f
C268 a_13175_4955# VGND 0
C269 VGND sky130_fd_sc_hd__mux2_1_0/a_76_199# 0.06911f
C270 a_16165_5035# VPB 0.00166f
C271 a_11230_5043# a_9723_5047# 0.00446f
C272 sky130_fd_sc_hd__inv_1_5/VPB VGND 0.02281f
C273 CLA_0/sky130_fd_sc_hd__and4_1_0/a_27_47# CLA_0/X -0.00351f
C274 VGND a_14225_2219# 0.09101f
C275 a_5999_2149# VGND 0.01281f
C276 a_11202_5917# a_12451_5917# -0.00146f
C277 a_2343_5417# VGND 0.01943f
C278 a_9360_5047# a_7899_5039# 0
C279 a_16095_2215# SUM -0
C280 a_9723_5047# a_8755_5489# 0
C281 CLA_0/sky130_fd_sc_hd__or2_1_0/A CLA_0/sky130_fd_sc_hd__or2_1_0/a_68_297# 0
C282 a_6726_5409# VGND 0
C283 a_9461_5471# VGND 0
C284 CLA_0/X VPB 0.00952f
C285 CLA_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# VGND 0.06112f
C286 a_12809_13987# VGND 0
C287 uio_out[7] uio_out[6] 0.03102f
C288 a_9290_2227# VGND 0.1057f
C289 a_9290_2227# a_9653_2227# -0.00146f
C290 a_10380_1777# VGND 0
C291 a_15644_5459# VGND 0.03671f
C292 a_13045_14187# VGND 0.04146f
C293 a_5606_2233# a_5735_1783# -0
C294 CLA_0/sky130_fd_sc_hd__or4_1_0/a_27_297# CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0
C295 CLA_0/sky130_fd_sc_hd__or4_1_0/C CLA_0/sky130_fd_sc_hd__or2_1_0/a_150_297# -0
C296 CLA_0/a_195_n767# VGND 0.00409f
C297 a_12105_15669# a_12045_13829# 0
C298 clk ena 0.03102f
C299 a_14888_5909# SUM 0
C300 a_13411_5829# VGND 0.0127f
C301 CLA_0/sky130_fd_sc_hd__and4_1_0/B CLA_0/sky130_fd_sc_hd__and4_1_0/a_109_47# -0
C302 a_16165_5035# a_15281_5825# 0
C303 VGND sky130_fd_sc_hd__mux2_1_0/VPB 0.06241f
C304 a_1920_2241# VPB 0
C305 CLA_0/X CLA_0/a_187_n2185# -0
C306 a_9360_5047# a_7506_5489# 0
C307 a_9959_13291# a_9845_14215# -0
C308 CLA_0/X a_9727_11527# 0
C309 ua[0] sky130_fd_sc_hd__mux4_1_0/a_750_97# 0
C310 CLA_0/sky130_fd_sc_hd__xor2_1_0/VPB VGND 0.02286f
C311 a_12292_5467# VGND 0
C312 a_16095_2215# a_15602_2131# 0
C313 CLA_0/sky130_fd_sc_hd__or4_1_0/C CLA_0/X 0.30643f
C314 a_11051_11919# VGND 0.00122f
C315 a_9753_4963# a_8755_5489# 0
C316 VPB a_12045_13829# 0
C317 VGND a_11553_1773# 0.02225f
C318 a_11455_4593# VGND 0
C319 a_11230_5043# a_12451_5917# 0
C320 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__inv_1_5/Y 0.10217f
C321 CLA_0/sky130_fd_sc_hd__or4_1_0/B VPB 0
C322 a_9332_5921# a_9695_5921# -0.00146f
C323 a_9715_16073# VGND 0.00347f
C324 a_14846_2215# VPB 0
C325 CLA_0/sky130_fd_sc_hd__and2_1_0/a_59_75# CLA_0/sky130_fd_sc_hd__and4_1_0/B -0
C326 a_9723_5047# a_9725_5837# 0
C327 a_5606_2233# VGND 0.10652f
C328 ui_in[0] sky130_fd_sc_hd__mux4_1_0/a_27_47# 0
C329 CLA_0/a_59_n3151# VGND 0.04734f
C330 a_4576_5413# VGND 0.00699f
C331 CLA_0/sky130_fd_sc_hd__and4_1_1/C CLA_0/sky130_fd_sc_hd__and4_1_1/VPB -0
C332 VGND a_10450_4597# 0
C333 VPB a_9695_5921# 0
C334 ui_in[1] sky130_fd_sc_hd__mux4_1_0/VPB 0.03979f
C335 a_2706_5051# a_3199_5501# 0
C336 uo_out[4] uo_out[3] 0.03102f
C337 a_15071_2131# VGND 0.00115f
C338 CLA_0/sky130_fd_sc_hd__and4_1_0/B CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0.0092f
C339 a_3169_2241# a_1920_2241# -0.00146f
C340 a_3199_5501# a_1950_5501# -0.00146f
C341 a_7635_5039# VGND 0
C342 a_9753_4963# a_9723_5047# -0
C343 CLA_0/X a_9675_12125# 0
C344 VGND sky130_fd_sc_hd__mux2_1_0/a_505_21# 0.1379f
C345 a_11427_5833# VGND 0.00157f
C346 a_7869_2145# VGND 0.01407f
C347 CLA_0/sky130_fd_sc_hd__or4_1_0/A CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0
C348 CLA_0/sky130_fd_sc_hd__or4_1_0/C CLA_0/sky130_fd_sc_hd__or4_1_0/B -0
C349 VPB a_3199_5501# 0
C350 a_9290_2227# a_8725_2229# 0.00511f
C351 CLA_0/sky130_fd_sc_hd__or4_1_0/VPB CLA_0/sky130_fd_sc_hd__or4_1_0/A -0.00133f
C352 a_11202_5917# a_11595_5833# -0
C353 sky130_fd_sc_hd__inv_1_4/A VGND 0.21173f
C354 a_5831_2149# VGND 0.0011f
C355 CLA_0/sky130_fd_sc_hd__and4_1_1/VPB CLA_0/sky130_fd_sc_hd__or4_1_0/B 0
C356 a_6392_5409# VGND 0.00697f
C357 VGND a_2706_5417# 0.00894f
C358 VGND CLA_0/sky130_fd_sc_hd__or2_1_0/a_150_297# 0
C359 a_12105_15669# a_11679_15219# 0
C360 CLA_0/sky130_fd_sc_hd__and4_1_1/a_27_47# VGND 0.03923f
C361 CLA_0/X a_9725_14509# 0
C362 a_13411_5463# a_14295_5039# 0
C363 a_5636_5493# a_6885_5493# -0.00146f
C364 a_10422_5837# VGND 0.00106f
C365 a_16165_5035# VGND 0.09749f
C366 CLA_0/sky130_fd_sc_hd__or4_1_0/a_109_297# CLA_0/X 0
C367 sky130_fd_sc_hd__inv_1_5/Y ui_in[1] 0.02018f
C368 a_10046_1777# VGND 0.02569f
C369 a_5606_2233# a_6855_2233# -0.00146f
C370 a_15281_5459# VGND 0.01642f
C371 sky130_fd_sc_hd__inv_1_2/Y CLA_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0
C372 ui_in[5] ui_in[4] 0.03102f
C373 uio_in[2] uio_in[1] 0.03102f
C374 uo_out[0] uo_out[1] 0.03102f
C375 a_14916_5035# a_14295_5039# 0.00446f
C376 a_4183_2153# VGND 0.01342f
C377 a_2343_5051# VGND 0.02053f
C378 CLA_0/sky130_fd_sc_hd__and4_1_1/a_303_47# CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0
C379 ui_in[1] ui_in[2] 0.03102f
C380 a_5636_5493# a_5069_5497# 0.00492f
C381 CLA_0/X a_9837_12547# 0.00128f
C382 a_13243_5829# VGND 0.00141f
C383 VPB a_14295_5039# 0.00228f
C384 CLA_0/X VGND 4.39357f
C385 CLA_0/sky130_fd_sc_hd__or2_1_0/B CLA_0/X 0
C386 a_11202_5917# VPB 0
C387 CLA_0/sky130_fd_sc_hd__and2_1_0/a_59_75# CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0
C388 a_11873_15219# a_12105_15669# -0
C389 a_13018_5913# a_12451_5917# 0.00492f
C390 CLA_0/X a_9727_11277# 0
C391 CLA_0/sky130_fd_sc_hd__or4_1_0/C CLA_0/sky130_fd_sc_hd__or2_1_0/VPB -0.00129f
C392 VGND CLA_0/sky130_fd_sc_hd__and2_1_0/VPB 0.03875f
C393 CLA_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# VGND 0.0196f
C394 CLA_0/sky130_fd_sc_hd__and4_1_1/C VGND 0.15806f
C395 a_14846_2215# ua[4] 0
C396 sky130_fd_sc_hd__mux4_1_0/a_834_97# ui_in[0] 0.00187f
C397 a_16095_2215# a_15239_2131# -0
C398 a_5636_5493# VPB 0
C399 a_13046_5039# a_14295_5039# -0.00146f
C400 VGND a_11385_1773# 0
C401 VGND a_14136_4589# 0
C402 sky130_fd_sc_hd__inv_1_2/Y CLA_0/sky130_fd_sc_hd__xor2_1_0/VPB 0
C403 a_11359_4593# VGND 0
C404 ui_in[1] VGND 0.50076f
C405 CLA_0/sky130_fd_sc_hd__or4_1_0/a_27_297# VPB 0
C406 a_8566_2145# VGND 0
C407 a_1920_2241# VGND 0.08933f
C408 a_3919_1787# VGND 0
C409 CLA_0/sky130_fd_sc_hd__or4_1_0/VPB CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0
C410 a_12479_5043# a_11595_5467# 0
C411 uio_out[1] uio_out[0] 0.03102f
C412 VGND a_12045_13829# 0.03188f
C413 ui_in[0] sky130_fd_sc_hd__mux4_1_0/a_247_21# -0
C414 VGND a_10116_4597# 0.02905f
C415 CLA_0/sky130_fd_sc_hd__or4_1_0/B VGND 0.23274f
C416 a_14846_2215# VGND 0.10989f
C417 a_8596_5405# a_8755_5489# -0
C418 a_8755_5489# a_9332_5921# 0
C419 CLA_0/X CLA_0/sky130_fd_sc_hd__or2_1_0/A 0
C420 a_4880_2153# VGND 0
C421 VGND sky130_fd_sc_hd__mux2_1_0/a_218_374# 0.00282f
C422 CLA_0/sky130_fd_sc_hd__and2_1_5/a_59_75# CLA_0/sky130_fd_sc_hd__and4_1_0/B -0
C423 CLA_0/a_195_n517# VGND 0.02568f
C424 a_11230_5043# VPB 0.00157f
C425 a_15017_5825# VGND 0
C426 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__mux4_1_0/a_1290_413# 0
C427 CLA_0/sky130_fd_sc_hd__or4_1_0/C CLA_0/sky130_fd_sc_hd__or4_1_0/a_27_297# 0
C428 CLA_0/VPB CLA_0/X 0.00689f
C429 a_15113_5459# VGND 0
C430 VGND a_9695_5921# 0.1627f
C431 a_5735_2149# VGND 0
C432 VPB a_8755_5489# 0
C433 a_10450_4963# VGND 0
C434 a_14066_1769# VGND 0
C435 a_2079_5051# VGND 0
C436 a_7476_2229# VPB 0
C437 CLA_0/sky130_fd_sc_hd__and2_1_5/VPB VGND 0.02314f
C438 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__inv_1_5/A 0.10823f
C439 a_6029_5409# VGND 0.01545f
C440 a_11595_5467# VGND 0.01604f
C441 VPB a_11213_12341# 0
C442 CLA_0/sky130_fd_sc_hd__or4_1_0/a_205_297# VGND 0
C443 uio_out[6] uio_out[5] 0.03102f
C444 uio_in[7] uio_in[6] 0.03102f
C445 a_9683_1777# VGND 0.01793f
C446 VGND a_3199_5501# 0.13369f
C447 sky130_fd_sc_hd__inv_1_2/Y CLA_0/sky130_fd_sc_hd__and4_1_1/a_27_47# 0.00861f
C448 VGND a_12250_2139# 0
C449 a_5069_5497# a_4213_5413# 0
C450 a_4546_2153# a_5039_2237# 0
C451 CLA_0/X a_9845_14215# 0.00124f
C452 VPB CLA_0/sky130_fd_sc_hd__or4_1_0/A 0
C453 a_6696_1783# VGND 0
C454 a_13147_5829# VGND 0
C455 CLA_0/sky130_fd_sc_hd__or2_1_0/VPB VGND 0.02525f
C456 a_7701_2145# VGND 0.0011f
C457 a_9723_5047# VPB 0.00228f
C458 CLA_0/sky130_fd_sc_hd__xor2_1_0/X CLA_0/sky130_fd_sc_hd__and4_1_1/a_197_47# -0
C459 sky130_fd_sc_hd__mux4_1_0/a_1290_413# VGND 0
C460 a_11160_2223# a_11553_1773# 0
C461 sky130_fd_sc_hd__inv_1_2/Y CLA_0/X 0.11818f
C462 a_8725_2229# a_8566_2145# -0
C463 CLA_0/sky130_fd_sc_hd__and3_1_0/VPB CLA_0/sky130_fd_sc_hd__or4_1_0/C -0
C464 a_9969_11727# a_9959_13291# -0
C465 ui_in[1] sky130_fd_sc_hd__mux4_1_0/a_668_97# 0.00464f
C466 sky130_fd_sc_hd__inv_1_5/A VGND 0.23315f
C467 a_11906_13629# VGND 0
C468 SUM a_14225_2219# -0
C469 VGND a_11289_1773# 0
C470 a_14295_5039# VGND 0.09988f
C471 VGND a_13802_4589# 0.02742f
C472 sky130_fd_sc_hd__inv_1_2/Y CLA_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0
C473 sky130_fd_sc_hd__inv_1_2/Y CLA_0/sky130_fd_sc_hd__and4_1_1/C 0.05432f
C474 VGND a_11679_15219# 0
C475 a_12320_4959# VGND 0
C476 CLA_0/X CLA_0/sky130_fd_sc_hd__and2_1_4/a_145_75# 0
C477 a_11202_5917# VGND 0.12857f
C478 VGND a_4045_5047# 0
C479 CLA_0/X CLA_0/a_n53_n3749# -0
C480 ua[0] sky130_fd_sc_hd__mux4_1_0/VPB 0.0095f
C481 CLA_0/sky130_fd_sc_hd__or4_1_0/C CLA_0/sky130_fd_sc_hd__or4_1_0/A -0.01788f
C482 CLA_0/sky130_fd_sc_hd__and2_1_5/a_59_75# CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0
C483 a_5636_5493# VGND 0.10644f
C484 CLA_0/sky130_fd_sc_hd__and4_1_0/B CLA_0/sky130_fd_sc_hd__and2_1_5/a_145_75# -0
C485 ui_in[1] sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.02448f
C486 CLA_0/a_n63_n2185# VGND 0.06519f
C487 VGND a_9753_4597# 0.02355f
C488 a_11230_5043# a_12479_5043# -0.00146f
C489 a_6029_5043# a_5636_5493# 0
C490 a_11331_5833# VGND 0
C491 uo_out[3] uo_out[2] 0.03102f
C492 CLA_0/sky130_fd_sc_hd__or4_1_0/a_27_297# VGND 0.0245f
C493 CLA_0/sky130_fd_sc_hd__and4_1_0/a_27_47# CLA_0/sky130_fd_sc_hd__xor2_1_0/X 0
C494 a_2313_1791# VGND 0.017f
C495 CLA_0/sky130_fd_sc_hd__or2_1_0/A CLA_0/sky130_fd_sc_hd__or2_1_0/VPB 0
C496 a_10088_5837# VGND 0.01153f
C497 a_13018_5913# VPB 0
C498 VPB a_5039_2237# 0
C499 sky130_fd_sc_hd__inv_1_2/Y CLA_0/sky130_fd_sc_hd__or4_1_0/B 0.002f
C500 VGND sky130_fd_sc_hd__mux2_1_0/a_535_374# 0.00127f
C501 a_11873_15219# VGND 0
C502 a_12451_5917# VPB 0.00104f
C503 VPB a_4183_1787# 0
C504 a_15017_5459# VGND 0
C505 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_0/VPB -0.00138f
C506 a_10116_4963# VGND 0.00727f
C507 a_13018_5913# a_13046_5039# 0
C508 a_13732_1769# VGND 0.02573f
C509 a_11767_15219# VGND 0.00137f
C510 a_12881_13987# VGND 0
C511 a_12409_2223# VPB 0
C512 a_5861_5409# VGND 0.00112f
C513 CLA_0/a_n55_n517# CLA_0/X -0
C514 a_11230_5043# VGND 0.11872f
C515 a_9515_1777# VGND 0
C516 VGND a_11916_2139# 0.00693f
C517 CLA_0/X CLA_0/a_69_n4715# 0.02088f
C518 a_16006_4951# VGND 0
C519 sky130_fd_sc_hd__inv_1_3/VPB sky130_fd_sc_hd__inv_1_4/A 0.00851f
C520 ua[6] VPB 0
C521 a_9360_5047# a_9695_5921# 0
C522 ui_in[4] ui_in[3] 0.03102f
C523 uio_in[1] uio_in[0] 0.03102f
C524 VPB a_9967_14959# 0
C525 VGND a_8755_5489# 0.10016f
C526 a_7476_2229# VGND 0.10915f
C527 CLA_0/sky130_fd_sc_hd__and3_1_0/VPB VGND 0.01956f
C528 CLA_0/sky130_fd_sc_hd__and3_1_0/VPB CLA_0/sky130_fd_sc_hd__or2_1_0/B -0
C529 a_6362_1783# VGND 0.02618f
C530 a_9837_12547# a_11213_12341# 0
C531 a_11958_5467# VGND 0.02766f
C532 a_14108_5463# VGND 0
C533 CLA_0/sky130_fd_sc_hd__or4_1_0/C CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0
C534 VGND a_11213_12341# 0.02974f
C535 a_11261_13361# VPB -0
C536 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__mux4_1_0/a_750_97# 0
C537 CLA_0/sky130_fd_sc_hd__or4_1_0/VPB CLA_0/sky130_fd_sc_hd__or4_1_0/C -0
C538 CLA_0/sky130_fd_sc_hd__and4_1_0/B VGND 0.77402f
C539 VGND a_4910_5047# 0
C540 CLA_0/a_197_n3749# CLA_0/X -0
C541 a_4015_1787# VGND 0
C542 CLA_0/sky130_fd_sc_hd__and4_1_1/VPB CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0.00242f
C543 ua[0] VGND 0.02135f
C544 a_9557_5837# a_9332_5921# -0
C545 a_14267_5913# a_14295_5039# 0.00177f
C546 ui_in[1] sky130_fd_sc_hd__mux4_1_0/a_27_413# 0.00288f
C547 CLA_0/sky130_fd_sc_hd__or4_1_0/A VGND 0.19457f
C548 a_14846_2215# a_16095_2215# -0.00146f
C549 VGND a_13439_4589# 0.01451f
C550 CLA_0/sky130_fd_sc_hd__xor2_1_0/a_285_47# VGND 0.00347f
C551 a_9723_5047# VGND 0.10765f
C552 a_11202_5917# a_11427_5467# 0
C553 a_4213_5413# VGND 0.01304f
C554 a_13018_5913# a_13243_5463# -0
C555 VGND a_2313_2157# 0.01589f
C556 a_16165_5035# SUM -0
C557 CLA_0/a_145_n3151# VGND 0.00275f
C558 a_16137_5909# a_15644_5825# 0
C559 CLA_0/sky130_fd_sc_hd__and4_1_0/a_109_47# VGND 0.00188f
C560 uio_out[0] uo_out[7] 0.03102f
C561 CLA_0/sky130_fd_sc_hd__or4_1_0/a_27_297# a_9845_14215# 0
C562 VGND a_9585_4597# 0
C563 a_12451_5917# a_12479_5043# 0.00177f
C564 sky130_fd_sc_hd__mux4_1_0/a_750_97# VGND 0.07286f
C565 a_7476_2229# a_6855_2233# 0.00446f
C566 a_5861_5043# a_5636_5493# -0
C567 a_11958_5833# VGND 0.01066f
C568 a_2145_1791# VGND 0
C569 uio_oe[2] uio_oe[1] 0.03102f
C570 a_3010_1791# VGND 0
C571 a_9725_5837# VGND 0.0198f
C572 CLA_0/X a_9559_11527# 0
C573 a_11261_13361# a_11321_14203# -0
C574 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__mux4_1_0/a_923_363# 0
C575 CLA_0/sky130_fd_sc_hd__and4_1_1/a_303_47# VGND 0.00102f
C576 VGND sky130_fd_sc_hd__mux2_1_0/a_218_47# 0.00146f
C577 a_10983_13753# VGND 0.00146f
C578 a_6885_5493# VPB 0
C579 a_14888_5909# a_15113_5459# -0
C580 VPB a_9847_10983# 0
C581 a_15978_5825# VGND 0
C582 CLA_0/sky130_fd_sc_hd__or4_1_0/a_109_297# CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0
C583 CLA_0/sky130_fd_sc_hd__and2_1_0/a_59_75# VGND 0.0542f
C584 CLA_0/X a_9683_13793# 0
C585 CLA_0/VPB CLA_0/sky130_fd_sc_hd__and4_1_0/B -0.00101f
C586 a_13369_1769# VGND 0.01786f
C587 a_9753_4963# VGND 0.00858f
C588 CLA_0/sky130_fd_sc_hd__and3_1_0/a_181_47# VGND 0
C589 a_13018_5913# VGND 0.12456f
C590 CLA_0/sky130_fd_sc_hd__and3_1_0/a_27_47# VGND 0.0328f
C591 a_5765_5409# VGND 0
C592 a_12105_15669# VPB -0
C593 a_8725_2229# a_7476_2229# -0.00146f
C594 VGND a_5039_2237# 0.08712f
C595 a_10895_13753# a_11321_14203# 0
C596 a_2049_2157# VGND 0
C597 a_5069_5497# VPB 0
C598 a_11089_13753# a_11321_14203# -0
C599 uio_out[5] uio_out[4] 0.03102f
C600 a_12409_2223# a_12976_2219# 0.00492f
C601 VPB a_9332_5921# 0
C602 a_12451_5917# VGND 0.11482f
C603 CLA_0/sky130_fd_sc_hd__and4_1_0/VPB CLA_0/X 0
C604 CLA_0/sky130_fd_sc_hd__xor2_1_0/X VGND 0.58975f
C605 uio_in[6] uio_in[5] 0.03102f
C606 a_14916_5035# a_16137_5909# 0
C607 VGND a_4183_1787# 0.01988f
C608 a_9419_1777# VGND 0
C609 VGND a_11553_2139# 0.01554f
C610 VPB a_1950_5501# 0
C611 a_15672_4951# VGND 0.00791f
C612 ua[5] VPB 0
C613 ui_in[1] ui_in[0] 5.44909f
C614 CLA_0/sky130_fd_sc_hd__or4_1_0/VPB VGND 0.01897f
C615 a_14916_5035# VPB 0.00157f
C616 a_12292_5833# VGND 0
C617 a_16137_5909# VPB 0
C618 CLA_0/a_19_n2185# VGND 0.00521f
C619 CLA_0/X CLA_0/sky130_fd_sc_hd__and2_1_4/VPB 0
C620 sky130_fd_sc_hd__mux4_1_0/a_757_363# sky130_fd_sc_hd__inv_1_5/Y 0
C621 a_8596_5039# a_8755_5489# 0
C622 a_12409_2223# VGND 0.08623f
C623 CLA_0/X a_9969_11727# 0.00232f
C624 CLA_0/sky130_fd_sc_hd__and3_1_0/a_109_47# VGND 0.00165f
C625 sky130_fd_sc_hd__mux4_1_0/a_923_363# VGND 0
C626 uio_oe[7] uio_oe[6] 0.03102f
C627 a_5999_1783# VGND 0.01636f
C628 a_13774_5463# VGND 0.02696f
C629 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__inv_1_4/VPB 0.01175f
C630 a_13201_1769# VGND 0
C631 ua[6] VGND 0
C632 a_9845_14215# CLA_0/sky130_fd_sc_hd__or4_1_0/A 0
C633 a_9967_14959# VGND 0.06763f
C634 a_9360_5047# a_8755_5489# 0
C635 CLA_0/sky130_fd_sc_hd__or4_1_0/a_277_297# CLA_0/X 0
C636 a_11230_5043# a_11359_4959# -0
C637 sky130_fd_sc_hd__inv_1_2/Y CLA_0/sky130_fd_sc_hd__and4_1_0/B 0
C638 VPB a_4213_5047# 0
C639 SUM a_9695_5921# -0
C640 a_9557_14759# VGND 0.00521f
C641 a_13046_5039# VPB 0.00168f
C642 CLA_0/sky130_fd_sc_hd__and4_1_0/a_303_47# CLA_0/X 0
C643 a_13045_14187# a_12809_13987# -0
C644 CLA_0/sky130_fd_sc_hd__and4_1_0/a_27_47# CLA_0/sky130_fd_sc_hd__or4_1_0/C -0
C645 a_10088_5471# a_8755_5489# 0
C646 VGND a_13271_4589# 0
C647 a_11261_13361# VGND 0.03105f
C648 ua[7] VPB 0
C649 CLA_0/X a_9717_12841# 0
C650 ua[0] sky130_fd_sc_hd__mux4_1_0/a_1478_413# 0.00699f
C651 sky130_fd_sc_hd__mux4_1_0/a_834_97# ui_in[1] 0.00243f
C652 sky130_fd_sc_hd__inv_1_3/VPB sky130_fd_sc_hd__inv_1_5/A 0
C653 SUM a_3199_5501# -0
C654 sky130_fd_sc_hd__mux4_1_0/a_757_363# VGND 0.00676f
C655 a_16137_5909# a_15281_5825# -0
C656 a_12479_5043# a_11595_5833# 0
C657 a_3169_2241# VPB 0
C658 CLA_0/sky130_fd_sc_hd__and4_1_1/a_109_47# CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0
C659 a_9360_5047# a_9723_5047# -0.00146f
C660 VGND a_9489_4597# 0
C661 uo_out[2] uo_out[1] 0.03102f
C662 a_10895_13753# VGND 0.00156f
C663 a_6726_5043# VGND 0
C664 a_11089_13753# VGND 0.00141f
C665 a_2049_1791# VGND 0
C666 a_9557_5837# VGND 0.00172f
C667 VPB a_11321_14203# 0
C668 a_11019_15169# VPB -0
C669 a_5999_2149# a_5606_2233# -0
C670 a_4546_2153# VGND 0.00698f
C671 a_3820_5497# a_3199_5501# 0.00446f
C672 a_12713_13987# VGND 0
C673 ui_in[1] sky130_fd_sc_hd__mux4_1_0/a_247_21# 0.09466f
C674 VGND sky130_fd_sc_hd__mux2_1_0/a_439_47# 0.00227f
C675 VGND a_9717_13091# 0.03032f
C676 a_8232_2145# VGND 0.00694f
C677 CLA_0/sky130_fd_sc_hd__and4_1_1/a_197_47# VGND 0.00153f
C678 uio_out[2] uio_out[1] 0.03102f
C679 VGND a_3919_2153# 0
C680 a_8262_5405# a_9332_5921# 0
C681 a_15644_5825# VGND 0.01798f
C682 ui_in[0] sky130_fd_sc_hd__mux4_1_0/a_1290_413# 0.13587f
C683 a_14267_5913# a_13018_5913# -0.00146f
C684 a_9585_4963# VGND 0.00111f
C685 VGND a_11986_4959# 0.00753f
C686 CLA_0/X a_9959_13291# 0.00237f
C687 SUM a_14295_5039# -0
C688 CLA_0/X CLA_0/sky130_fd_sc_hd__or2_1_0/a_68_297# 0
C689 sky130_fd_sc_hd__inv_1_2/Y CLA_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 0
C690 a_8232_1779# VGND 0.02546f
C691 a_11595_5833# VGND 0.01174f
C692 SUM a_11202_5917# 0
C693 a_9837_12547# a_9847_10983# -0
C694 CLA_0/a_n55_n517# CLA_0/sky130_fd_sc_hd__and4_1_0/B -0
C695 a_6885_5493# VGND 0.0915f
C696 sky130_fd_sc_hd__inv_1_4/A sky130_fd_sc_hd__inv_1_5/VPB 0
C697 a_12479_5043# VPB 0.00242f
C698 CLA_0/sky130_fd_sc_hd__or4_1_0/VPB a_9845_14215# 0
C699 VGND a_11385_2139# 0.0011f
C700 a_15309_4951# VGND 0.00787f
C701 VGND a_9847_10983# 0.05412f
C702 ui_in[3] ui_in[2] 0.03102f
C703 a_16165_5035# sky130_fd_sc_hd__mux2_1_0/a_76_199# 0
C704 sky130_fd_sc_hd__inv_1_2/Y CLA_0/sky130_fd_sc_hd__xor2_1_0/X 0.23966f
C705 CLA_0/sky130_fd_sc_hd__and2_1_5/a_59_75# VGND 0.02473f
C706 a_8262_5039# a_8755_5489# 0
C707 a_12105_15669# VGND 0.04564f
C708 a_5831_1783# VGND 0
C709 a_13411_5463# VGND 0.01368f
C710 a_5069_5497# VGND 0.08677f
C711 a_8596_5405# VGND 0
C712 a_13046_5039# a_12479_5043# 0.00492f
C713 CLA_0/a_187_n2435# VGND 0.00364f
C714 a_11019_15169# a_11321_14203# -0
C715 a_13105_1769# VGND 0
C716 a_2706_5051# VGND 0.02639f
C717 VGND a_9332_5921# 0.11077f
C718 CLA_0/X a_9549_13091# 0
C719 CLA_0/X CLA_0/sky130_fd_sc_hd__and2_1_4/a_59_75# -0
C720 VGND a_1950_5501# 0.08905f
C721 CLA_0/sky130_fd_sc_hd__and4_1_0/a_27_47# VGND 0.0546f
C722 VPB a_12976_2219# 0
C723 ua[5] VGND 0.00178f
C724 a_14975_2131# VGND 0
C725 sky130_fd_sc_hd__mux2_1_0/a_505_21# sky130_fd_sc_hd__mux2_1_0/VPB -0
C726 a_14916_5035# VGND 0.12124f
C727 a_16137_5909# VGND 0.12087f
C728 sky130_fd_sc_hd__inv_1_2/VPB VGND 0.03516f
C729 VPB a_9837_12547# 0
C730 ui_in[1] sky130_fd_sc_hd__mux4_1_0/a_193_413# 0.00324f
C731 a_9725_14759# VGND 0.02439f
C732 sky130_fd_sc_hd__inv_1_5/Y sky130_fd_sc_hd__mux4_1_0/VPB 0.02307f
C733 VPB VGND 2.02615f
C734 a_9725_5471# a_8755_5489# 0
C735 a_9653_2227# VPB 0
C736 VGND a_13175_4589# 0
C737 CLA_0/a_155_n4715# VGND 0.00186f
C738 sky130_fd_sc_hd__mux4_1_0/a_1290_413# sky130_fd_sc_hd__mux4_1_0/a_247_21# -0.00452f
C739 a_10857_14747# VGND 0.00195f
C740 ui_in[7] uio_in[0] 0.03102f
C741 a_16165_5035# sky130_fd_sc_hd__mux2_1_0/VPB 0.00175f
C742 sky130_fd_sc_hd__mux4_1_0/a_27_413# sky130_fd_sc_hd__mux4_1_0/a_750_97# -0
C743 VGND a_4213_5047# 0.0194f
C744 a_3790_2237# a_5039_2237# -0.00146f
C745 a_13046_5039# VGND 0.11794f
C746 uo_out[7] uo_out[6] 0.03102f
C747 SUM a_8755_5489# -0
C748 ua[7] VGND 0
C749 a_15936_1765# VGND 0
C750 sky130_fd_sc_hd__inv_1_5/A sky130_fd_sc_hd__inv_1_4/VPB 0.00953f
C751 a_6392_5043# VGND 0.02568f
C752 CLA_0/a_187_n2185# VGND 0.02415f
C753 a_3040_5417# VGND 0
C754 a_9845_14215# a_9717_13091# -0
C755 a_9461_5837# VGND 0.00106f
C756 a_3010_2157# VGND 0
C757 a_5831_2149# a_5606_2233# -0
C758 a_9725_5471# a_9723_5047# 0
C759 a_9727_11527# VGND 0.02361f
C760 a_4045_5413# VGND 0.00111f
C761 CLA_0/sky130_fd_sc_hd__or4_1_0/C VGND 0.39841f
C762 CLA_0/sky130_fd_sc_hd__or4_1_0/C CLA_0/sky130_fd_sc_hd__or2_1_0/B -0.00108f
C763 a_8232_1779# a_8725_2229# 0
C764 a_3169_2241# VGND 0.13397f
C765 a_7899_5405# a_9332_5921# 0
C766 sky130_fd_sc_hd__mux4_1_0/VPB VGND 0.02744f
C767 a_15281_5825# VGND 0.01246f
C768 CLA_0/sky130_fd_sc_hd__and4_1_1/VPB VGND 0.01711f
C769 a_11160_2223# a_11553_2139# -0
C770 a_14846_2215# a_14225_2219# 0.00446f
C771 a_9489_4963# VGND 0
C772 a_16006_4585# VGND 0
C773 a_11019_15169# VGND 0.02409f
C774 VGND a_11623_4959# 0.00844f
C775 VGND a_11321_14203# 0.05088f
C776 a_6855_2233# VPB 0
C777 ua[0] ui_in[0] 0.53168f
C778 SUM a_9723_5047# -0
C779 CLA_0/sky130_fd_sc_hd__and2_1_5/a_145_75# VGND 0.00202f
C780 a_7869_1779# VGND 0.02049f
C781 a_11160_2223# a_12409_2223# -0.00146f
C782 uio_out[4] uio_out[3] 0.03102f
C783 uio_in[5] uio_in[4] 0.03102f
C784 VGND a_11289_2139# 0
C785 a_15141_4951# VGND 0.00124f
C786 CLA_0/sky130_fd_sc_hd__and4_1_0/VPB CLA_0/sky130_fd_sc_hd__and4_1_0/B -0
C787 a_16165_5035# sky130_fd_sc_hd__mux2_1_0/a_505_21# 0
C788 CLA_0/X CLA_0/a_59_n3151# -0
C789 a_9675_12125# VGND 0.00275f
C790 VGND CLA_0/a_153_n1483# 0.00278f
C791 uio_oe[6] uio_oe[5] 0.03102f
C792 a_5735_1783# VGND 0
C793 a_13243_5463# VGND 0
C794 sky130_fd_sc_hd__inv_1_5/Y VGND 1.32539f
C795 VGND a_10380_2143# 0
C796 a_8262_5405# VGND 0.00798f
C797 a_8725_2229# VPB 0
C798 a_14066_2135# VGND 0
C799 a_3040_5051# VGND 0
C800 a_12479_5043# VGND 0.09961f
C801 ua[4] a_15071_1765# 0
C802 ua[4] VGND 0.0019f
C803 sky130_fd_sc_hd__mux4_1_0/a_750_97# ui_in[0] 0.01723f
C804 CLA_0/sky130_fd_sc_hd__or4_1_0/C CLA_0/sky130_fd_sc_hd__or2_1_0/A -0
C805 uio_oe[3] uio_oe[2] 0.03102f
C806 a_14267_5913# VPB 0
C807 VPB a_9845_14215# 0
C808 a_9725_14509# VGND 0.00409f
C809 a_16165_5035# a_15281_5459# 0
C810 sky130_fd_sc_hd__inv_1_2/Y sky130_fd_sc_hd__inv_1_2/VPB 0.00969f
C811 CLA_0/sky130_fd_sc_hd__or4_1_0/a_109_297# VGND 0
C812 a_9360_5047# a_9332_5921# 0
C813 a_13018_5913# SUM 0
C814 SUM a_5039_2237# -0
C815 CLA_0/X CLA_0/sky130_fd_sc_hd__or2_1_0/a_150_297# -0
C816 VGND a_12976_2219# 0.10623f
C817 sky130_fd_sc_hd__inv_1_5/A sky130_fd_sc_hd__inv_1_5/VPB 0.01139f
C818 a_14267_5913# a_13046_5039# 0
C819 a_8755_5489# a_7506_5489# -0.00146f
C820 SUM a_12451_5917# -0
C821 VGND a_9837_12547# 0.04734f
C822 a_15071_1765# VGND 0
C823 a_9360_5047# VPB 0.0017f
C824 CLA_0/sky130_fd_sc_hd__or2_1_0/B VGND 0.12155f
C825 a_9653_2227# VGND 0.09125f
C826 SUM a_12409_2223# -0
C827 a_15602_1765# VGND 0.02574f
C828 a_6029_5043# VGND 0.01991f
C829 a_14136_4955# VGND 0
C830 CLA_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# VGND 0.00465f
C831 a_2175_5417# VGND 0.00147f
C832 a_5735_2149# a_5606_2233# -0
C833 a_7701_1779# VGND 0
C834 a_9727_11277# VGND 0.00312f
C835 a_11230_5043# a_11623_4593# 0
C836 a_3949_5413# VGND 0
C837 a_15113_5825# VGND 0.00139f
C838 CLA_0/sky130_fd_sc_hd__and4_1_0/VPB CLA_0/sky130_fd_sc_hd__xor2_1_0/X -0
C839 a_9845_14215# a_11321_14203# -0
C840 CLA_0/sky130_fd_sc_hd__and4_1_1/C CLA_0/X -0.00844f
C841 a_11160_2223# a_11385_2139# -0
C842 a_13411_5829# a_14295_5039# 0
C843 a_15672_4585# VGND 0.02903f
C844 VGND a_11455_4959# 0.00139f
C845 a_10422_5471# VGND 0
C846 sky130_fd_sc_hd__mux4_1_0/a_750_97# sky130_fd_sc_hd__mux4_1_0/a_247_21# -0
C847 sky130_fd_sc_hd__inv_1_2/Y CLA_0/sky130_fd_sc_hd__and4_1_1/VPB 0.00632f
C848 uio_oe[1] uio_oe[0] 0.03102f
C849 a_2079_5417# VGND 0
C850 a_3949_5047# VGND 0
C851 ua[1] VNB 0.14696f
C852 ua[2] VNB 0.14696f
C853 ua[3] VNB 0.14696f
C854 ua[4] VNB 0.14465f
C855 ua[5] VNB 0.14471f
C856 ua[6] VNB 0.14538f
C857 ua[7] VNB 0.1455f
C858 ena VNB 0.07038f
C859 clk VNB 0.04288f
C860 rst_n VNB 0.04288f
C861 ui_in[2] VNB 0.04288f
C862 ui_in[3] VNB 0.04288f
C863 ui_in[4] VNB 0.04288f
C864 ui_in[5] VNB 0.04288f
C865 ui_in[6] VNB 0.04288f
C866 ui_in[7] VNB 0.04288f
C867 uio_in[0] VNB 0.04288f
C868 uio_in[1] VNB 0.04288f
C869 uio_in[2] VNB 0.04288f
C870 uio_in[3] VNB 0.04288f
C871 uio_in[4] VNB 0.04288f
C872 uio_in[5] VNB 0.04288f
C873 uio_in[6] VNB 0.04288f
C874 uio_in[7] VNB 0.04288f
C875 uo_out[0] VNB 0.04288f
C876 uo_out[1] VNB 0.04288f
C877 uo_out[2] VNB 0.04288f
C878 uo_out[3] VNB 0.04288f
C879 uo_out[4] VNB 0.04288f
C880 uo_out[5] VNB 0.04288f
C881 uo_out[6] VNB 0.04288f
C882 uo_out[7] VNB 0.04288f
C883 uio_out[0] VNB 0.04288f
C884 uio_out[1] VNB 0.04288f
C885 uio_out[2] VNB 0.04288f
C886 uio_out[3] VNB 0.04288f
C887 uio_out[4] VNB 0.04288f
C888 uio_out[5] VNB 0.04288f
C889 uio_out[6] VNB 0.04288f
C890 uio_out[7] VNB 0.04288f
C891 uio_oe[0] VNB 0.04288f
C892 uio_oe[1] VNB 0.04288f
C893 uio_oe[2] VNB 0.04288f
C894 uio_oe[3] VNB 0.04288f
C895 uio_oe[4] VNB 0.04288f
C896 uio_oe[5] VNB 0.04288f
C897 uio_oe[6] VNB 0.04288f
C898 uio_oe[7] VNB 0.07038f
C899 a_16095_2215# VNB 0.27343f
C900 a_14846_2215# VNB 0.13081f
C901 a_12976_2219# VNB 0.13025f
C902 a_14225_2219# VNB 0.26543f
C903 a_12409_2223# VNB 0.26466f
C904 a_11160_2223# VNB 0.13081f
C905 a_9653_2227# VNB 0.26543f
C906 a_9290_2227# VNB 0.13016f
C907 a_7476_2229# VNB 0.13081f
C908 a_8725_2229# VNB 0.26452f
C909 a_6855_2233# VNB 0.26543f
C910 a_5606_2233# VNB 0.13025f
C911 a_5039_2237# VNB 0.26466f
C912 a_3790_2237# VNB 0.13081f
C913 a_1920_2241# VNB 0.1359f
C914 a_3169_2241# VNB 0.26543f
C915 a_16165_5035# VNB 0.26397f
C916 a_14916_5035# VNB 0.12906f
C917 a_13046_5039# VNB 0.12849f
C918 a_14295_5039# VNB 0.26214f
C919 a_12479_5043# VNB 0.26136f
C920 a_11230_5043# VNB 0.12906f
C921 a_9723_5047# VNB 0.26214f
C922 a_9360_5047# VNB 0.13349f
C923 a_16137_5909# VNB 0.27134f
C924 a_14888_5909# VNB 0.12984f
C925 a_14267_5913# VNB 0.26335f
C926 a_13018_5913# VNB 0.12928f
C927 a_12451_5917# VNB 0.26257f
C928 a_11202_5917# VNB 0.12984f
C929 a_9695_5921# VNB 0.26335f
C930 a_9332_5921# VNB 0.13493f
C931 a_7506_5489# VNB 0.13081f
C932 a_8755_5489# VNB 0.27172f
C933 a_5636_5493# VNB 0.13025f
C934 a_6885_5493# VNB 0.26543f
C935 a_5069_5497# VNB 0.26466f
C936 a_3820_5497# VNB 0.13081f
C937 a_3199_5501# VNB 0.26543f
C938 a_1950_5501# VNB 0.1359f
C939 a_11213_12341# VNB 0.17706f
C940 a_11261_13361# VNB 0.17719f
C941 a_12045_13829# VNB 0.15387f
C942 a_11321_14203# VNB 0.17489f
C943 a_13045_14187# VNB 0.16291f
C944 a_11019_15169# VNB 0.17706f
C945 a_12105_15669# VNB 0.17489f
C946 a_9835_15779# VNB 0.17706f
C947 a_9957_16523# VNB 0.25457f
C948 sky130_fd_sc_hd__inv_1_4/A VNB 0.40476f
C949 sky130_fd_sc_hd__inv_1_3/VPB VNB 0.33898f
C950 a_6029_5409# VNB 0.01584f
C951 a_6392_5409# VNB 0.01578f
C952 a_6029_5043# VNB 0.00484f
C953 a_6392_5043# VNB 0.00345f
C954 a_15309_4951# VNB 0.01584f
C955 a_15672_4951# VNB 0.01578f
C956 a_15309_4585# VNB 0.00484f
C957 a_15672_4585# VNB 0.00345f
C958 sky130_fd_sc_hd__inv_1_2/VPB VNB 0.33898f
C959 a_7899_5405# VNB 0.01584f
C960 a_8262_5405# VNB 0.01578f
C961 a_7899_5039# VNB 0.00484f
C962 a_8262_5039# VNB 0.00345f
C963 sky130_fd_sc_hd__inv_1_0/VPB VNB 0.33898f
C964 a_13439_4955# VNB 0.01584f
C965 a_13802_4955# VNB 0.01578f
C966 a_13439_4589# VNB 0.00484f
C967 a_13802_4589# VNB 0.00345f
C968 sky130_fd_sc_hd__mux2_1_0/VPB VNB 0.87055f
C969 sky130_fd_sc_hd__mux2_1_0/a_505_21# VNB 0.24676f
C970 sky130_fd_sc_hd__mux2_1_0/a_76_199# VNB 0.13947f
C971 a_9753_4963# VNB 0.01584f
C972 a_10116_4963# VNB 0.01578f
C973 a_9753_4597# VNB 0.00484f
C974 a_10116_4597# VNB 0.00345f
C975 a_11553_2139# VNB 0.01584f
C976 a_11916_2139# VNB 0.01578f
C977 a_11553_1773# VNB 0.00484f
C978 a_11916_1773# VNB 0.00345f
C979 a_9683_2143# VNB 0.01584f
C980 a_10046_2143# VNB 0.01578f
C981 a_9683_1777# VNB 0.00484f
C982 a_10046_1777# VNB 0.00345f
C983 a_11623_4959# VNB 0.01584f
C984 a_11986_4959# VNB 0.01578f
C985 a_11623_4593# VNB 0.00484f
C986 a_11986_4593# VNB 0.00345f
C987 a_13369_2135# VNB 0.01584f
C988 a_13732_2135# VNB 0.01578f
C989 a_13369_1769# VNB 0.00484f
C990 a_13732_1769# VNB 0.00345f
C991 a_13411_5829# VNB 0.01584f
C992 a_13774_5829# VNB 0.01578f
C993 a_13411_5463# VNB 0.00484f
C994 a_13774_5463# VNB 0.00345f
C995 a_15281_5825# VNB 0.01584f
C996 a_15644_5825# VNB 0.01578f
C997 a_15281_5459# VNB 0.00484f
C998 a_15644_5459# VNB 0.00345f
C999 a_9725_5837# VNB 0.01584f
C1000 a_10088_5837# VNB 0.01578f
C1001 a_9725_5471# VNB 0.00484f
C1002 a_10088_5471# VNB 0.00345f
C1003 a_15239_2131# VNB 0.01584f
C1004 a_15602_2131# VNB 0.01578f
C1005 a_15239_1765# VNB 0.00484f
C1006 a_15602_1765# VNB 0.00345f
C1007 a_5999_2149# VNB 0.01584f
C1008 a_6362_2149# VNB 0.01578f
C1009 a_5999_1783# VNB 0.00484f
C1010 a_6362_1783# VNB 0.00345f
C1011 a_7869_2145# VNB 0.01584f
C1012 a_8232_2145# VNB 0.01578f
C1013 a_7869_1779# VNB 0.00484f
C1014 a_8232_1779# VNB 0.00345f
C1015 a_11595_5833# VNB 0.01584f
C1016 a_11958_5833# VNB 0.01578f
C1017 a_11595_5467# VNB 0.00484f
C1018 a_11958_5467# VNB 0.00345f
C1019 a_4183_2153# VNB 0.01584f
C1020 a_4546_2153# VNB 0.01578f
C1021 a_4183_1787# VNB 0.00484f
C1022 a_4546_1787# VNB 0.00345f
C1023 a_4213_5413# VNB 0.01584f
C1024 a_4576_5413# VNB 0.01578f
C1025 a_4213_5047# VNB 0.00484f
C1026 a_4576_5047# VNB 0.00345f
C1027 SUM VNB 1.43445f
C1028 VPB VNB 39.04759f
C1029 a_2313_2157# VNB 0.01584f
C1030 a_2676_2157# VNB 0.01578f
C1031 a_2313_1791# VNB 0.00484f
C1032 a_2676_1791# VNB 0.00345f
C1033 a_2343_5417# VNB 0.01584f
C1034 a_2706_5417# VNB 0.01578f
C1035 a_2343_5051# VNB 0.00484f
C1036 a_2706_5051# VNB 0.00345f
C1037 a_9847_10983# VNB 0.1752f
C1038 a_9969_11727# VNB 0.24712f
C1039 a_9837_12547# VNB 0.17114f
C1040 a_9959_13291# VNB 0.24424f
C1041 a_9845_14215# VNB 0.16601f
C1042 a_9967_14959# VNB 0.24496f
C1043 a_9727_11527# VNB 0.00137f
C1044 a_9725_14759# VNB 0.00137f
C1045 a_9715_16323# VNB 0.00137f
C1046 VGND VNB 0.20612p
C1047 a_9717_13091# VNB 0.00137f
C1048 CLA_0/a_69_n4715# VNB 0.1752f
C1049 CLA_0/a_n53_n3749# VNB 0.24712f
C1050 CLA_0/a_59_n3151# VNB 0.17114f
C1051 CLA_0/a_n63_n2185# VNB 0.24424f
C1052 CLA_0/a_67_n1483# VNB 0.17003f
C1053 CLA_0/a_n55_n517# VNB 0.24496f
C1054 CLA_0/a_197_n3749# VNB 0.00137f
C1055 CLA_0/a_195_n517# VNB 0.00137f
C1056 CLA_0/sky130_fd_sc_hd__xor2_1_0/VPB VNB 0.69336f
C1057 CLA_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# VNB 0.00137f
C1058 CLA_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# VNB 0.25457f
C1059 CLA_0/sky130_fd_sc_hd__or2_1_0/B VNB 0.46058f
C1060 CLA_0/sky130_fd_sc_hd__and3_1_0/VPB VNB 0.51617f
C1061 CLA_0/sky130_fd_sc_hd__and3_1_0/a_27_47# VNB 0.17719f
C1062 CLA_0/sky130_fd_sc_hd__or4_1_0/B VNB 0.799f
C1063 CLA_0/sky130_fd_sc_hd__or4_1_0/VPB VNB 0.60476f
C1064 CLA_0/sky130_fd_sc_hd__or4_1_0/a_27_297# VNB 0.16291f
C1065 sky130_fd_sc_hd__inv_1_2/Y VNB 2.47775f
C1066 CLA_0/sky130_fd_sc_hd__and4_1_1/VPB VNB 0.69336f
C1067 CLA_0/sky130_fd_sc_hd__and4_1_1/a_27_47# VNB 0.17489f
C1068 CLA_0/sky130_fd_sc_hd__or2_1_0/A VNB 0.31965f
C1069 CLA_0/sky130_fd_sc_hd__xor2_1_0/X VNB 1.89098f
C1070 CLA_0/sky130_fd_sc_hd__and4_1_0/B VNB 0.74819f
C1071 CLA_0/sky130_fd_sc_hd__and4_1_0/VPB VNB 0.69336f
C1072 CLA_0/sky130_fd_sc_hd__and4_1_0/a_27_47# VNB 0.17489f
C1073 CLA_0/sky130_fd_sc_hd__or4_1_0/A VNB 0.42983f
C1074 CLA_0/sky130_fd_sc_hd__or2_1_0/VPB VNB 0.51617f
C1075 CLA_0/sky130_fd_sc_hd__or2_1_0/a_68_297# VNB 0.15387f
C1076 CLA_0/sky130_fd_sc_hd__and4_1_1/C VNB 0.33836f
C1077 CLA_0/sky130_fd_sc_hd__and2_1_5/VPB VNB 0.51617f
C1078 CLA_0/sky130_fd_sc_hd__and2_1_5/a_59_75# VNB 0.17706f
C1079 CLA_0/sky130_fd_sc_hd__or4_1_0/C VNB 1.43825f
C1080 CLA_0/sky130_fd_sc_hd__and2_1_4/VPB VNB 0.51617f
C1081 CLA_0/sky130_fd_sc_hd__and2_1_4/a_59_75# VNB 0.17706f
C1082 CLA_0/X VNB 7.24455f
C1083 CLA_0/VPB VNB 3.62859f
C1084 CLA_0/sky130_fd_sc_hd__and2_1_0/VPB VNB 0.51617f
C1085 CLA_0/sky130_fd_sc_hd__and2_1_0/a_59_75# VNB 0.17706f
C1086 CLA_0/a_187_n2185# VNB 0.00137f
C1087 ua[0] VNB 9.60658f
C1088 ui_in[0] VNB 8.82066f
C1089 ui_in[1] VNB 8.40071f
C1090 sky130_fd_sc_hd__inv_1_5/Y VNB 3.59173f
C1091 sky130_fd_sc_hd__mux4_1_0/VPB VNB 1.9337f
C1092 sky130_fd_sc_hd__mux4_1_0/a_834_97# VNB 0.02499f
C1093 sky130_fd_sc_hd__mux4_1_0/a_668_97# VNB 0.02039f
C1094 sky130_fd_sc_hd__mux4_1_0/a_27_47# VNB 0.04207f
C1095 sky130_fd_sc_hd__mux4_1_0/a_1478_413# VNB 0.16413f
C1096 sky130_fd_sc_hd__mux4_1_0/a_1290_413# VNB 0.2199f
C1097 sky130_fd_sc_hd__mux4_1_0/a_750_97# VNB 0.04192f
C1098 sky130_fd_sc_hd__mux4_1_0/a_757_363# VNB 0.00666f
C1099 sky130_fd_sc_hd__mux4_1_0/a_247_21# VNB 0.34344f
C1100 sky130_fd_sc_hd__mux4_1_0/a_193_413# VNB 0.00373f
C1101 sky130_fd_sc_hd__mux4_1_0/a_27_413# VNB 0.02865f
C1102 sky130_fd_sc_hd__inv_1_5/VPB VNB 0.33898f
C1103 sky130_fd_sc_hd__inv_1_5/A VNB 0.45825f
C1104 sky130_fd_sc_hd__inv_1_4/VPB VNB 0.33898f
.ends

