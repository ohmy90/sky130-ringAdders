* NGSPICE file created from tt_um_ohmy90_flat_adders.ext - technology: sky130A

.subckt tt_um_ohmy90_flat_adders clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5]
+ ua[6] ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7]
+ uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
+ uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
+ uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
+ VDPWR VGND
X0 VDPWR VGND a_12281_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X1 VDPWR a_9703_16093# a_11501_15239# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X2 a_24234_14385# ui_in[0] a_24152_14385# VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.10855 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X3 VGND a_9381_11547# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr d=10010,284
X4 a_16793_4785# a_15711_4547# a_17210_4895# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X5 VDPWR VGND a_16539_5473# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X6 a_16679_4895# VDPWR a_16583_4895# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X7 a_4711_15373# VGND a_4625_15373# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X8 a_5174_5409# VDPWR a_4423_5299# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X9 a_18625_4938# a_17733_4529# a_18553_4938# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=7728,268
X10 VGND VGND a_9369_16343# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X11 VDPWR VGND a_2313_1791# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X12 a_12533_5715# a_11411_5471# a_12950_5825# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X13 a_14545_5467# a_14491_5723# a_14152_5441# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X14 a_1950_5025# a_2217_5025# a_2175_5051# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X15 a_12419_5825# VDPWR a_12323_5825# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X16 VDPWR a_12194_5433# a_12142_5459# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X17 a_16033_2159# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X18 a_17236_5839# VDPWR a_16485_5729# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X19 a_4513_14775# VDPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X20 a_6129_12927# a_4913_13781# a_6057_12927# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=1764,126
X21 VGND VGND a_16297_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X22 VGND a_9381_11547# a_9631_11547# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=3.156 pd=47.08 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X23 a_7113_13395# a_6862_13645# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4010,197 d=6760,364
X24 a_12323_5459# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X25 a_11255_13773# a_10717_13773# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X26 VDPWR VGND a_7032_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X27 a_11501_15239# a_8193_13753# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X28 a_4383_2153# a_4329_2043# a_3990_1761# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X29 a_14281_5833# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X30 VDPWR VGND a_4587_13107# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X31 a_9631_11297# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X32 a_8169_1793# VDPWR a_8073_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X33 a_14771_4803# a_13709_4553# a_15188_4547# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X34 a_22274_16171# a_21506_16181# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X35 a_2175_5417# VDPWR a_2079_5417# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X36 a_6089_11935# VGND a_6003_11935# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X37 VDPWR VDPWR a_14596_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X38 VGND a_11888_1767# a_11836_1793# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X39 a_10289_2159# a_10235_2049# a_9896_1767# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X40 a_12697_14007# a_9781_10553# a_12615_14007# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2772,150
X41 VDPWR VGND a_4597_11543# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X42 a_7221_1787# a_6281_2043# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X43 VDPWR VDPWR a_9491_15377# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X44 VDPWR VDPWR a_6792_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X45 VDPWR VDPWR a_14825_4547# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X46 a_12644_2159# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X47 VDPWR VDPWR a_16660_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X48 VDPWR VDPWR a_16847_4529# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X49 a_9629_14779# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X50 a_10525_5837# a_10471_5727# a_10132_5445# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X51 VDPWR VGND a_14233_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X52 a_5942_1761# a_5269_1787# a_6167_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X53 sky130_fd_sc_hd__mux4_1_0.A3 a_18625_4938# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=6334,279 d=10400,504
X54 VDPWR VDPWR a_10289_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X55 VGND a_1920_1765# a_1868_1791# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X56 a_8038_5023# a_7315_5043# a_8263_5049# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X57 VDPWR sky130_fd_sc_hd__mux4_1_0.A1 a_6629_15387# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X58 a_7126_5409# VDPWR a_6375_5299# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X59 VDPWR VDPWR a_4753_16339# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X60 VGND VGND a_5174_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X61 a_12769_4809# a_11439_4597# a_13186_4553# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X62 VDPWR VDPWR a_4746_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X63 VDPWR VDPWR a_8431_5049# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X64 a_4903_15345# a_4625_15373# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X65 VDPWR VDPWR a_4763_14775# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X66 VDPWR VDPWR a_12823_4553# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X67 a_13520_4919# VDPWR a_12769_4809# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X68 a_4913_13781# a_4635_13809# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X69 VGND VDPWR a_17210_4895# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X70 a_10160_4571# VDPWR a_10385_4963# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X71 a_4084_5017# a_3229_5051# a_4309_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X72 VGND VGND a_14930_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X73 a_16847_4895# a_15711_4547# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X74 a_4723_10577# VGND a_4637_10577# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X75 a_15431_5467# a_14491_5723# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X76 a_4587_13107# VDPWR a_4505_13107# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X77 VGND VGND a_9381_11547# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X78 a_16146_5447# a_15431_5467# a_16371_5839# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X79 a_14377_5467# VDPWR a_14281_5467# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X80 a_2079_5051# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X81 a_16902_5839# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X82 a_9223_1793# a_8283_2049# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X83 VGND VDPWR a_16539_5839# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X84 a_4597_11543# VDPWR a_4515_11543# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X85 a_9491_15377# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X86 a_6944_13645# a_6329_12927# a_6862_13645# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X87 a_10132_5445# VGND a_10357_5471# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X88 VGND a_13840_1767# a_13788_1793# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X89 a_8700_1793# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X90 a_4635_13809# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X91 a_2706_5417# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X92 VDPWR VGND a_2343_5051# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X93 VGND a_4513_14775# a_4847_14525# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X94 a_10986_2159# VDPWR a_10235_2049# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X95 a_4215_2153# VDPWR a_4119_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X96 VGND a_11979_13399# a_12615_14007# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2268,138 d=4075,198
X97 VGND VGND a_12978_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X98 a_9779_13785# a_9501_13813# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X99 a_10888_5471# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X100 a_18625_4938# a_17425_5473# a_18625_5265# VGND sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=3990,179
X101 VGND a_4503_16339# a_4837_16089# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X102 a_8337_1793# a_7221_1787# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X103 VGND VGND a_7126_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X104 VDPWR VDPWR a_10525_5471# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X105 a_14825_4547# a_13709_4553# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X106 a_8377_5305# a_7315_5043# a_8794_5415# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X107 VDPWR VDPWR a_9503_10581# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X108 VDPWR a_8038_5023# a_7986_5049# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X109 a_11888_1767# a_11175_1793# a_12113_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X110 VGND sky130_fd_sc_hd__mux4_1_0.A1 a_23511_14335# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X111 VGND a_3990_1761# a_3938_1787# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X112 a_9371_13111# VDPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X113 VDPWR VDPWR a_6698_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X114 a_6805_15235# a_4847_14525# a_6717_15235# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X115 a_9705_12861# VDPWR a_9621_12861# VGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X116 VGND VGND a_13520_4919# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X117 VDPWR VGND a_10289_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X118 a_8167_5049# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X119 a_1920_1765# a_2187_1765# a_2145_2157# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X120 a_5269_1787# a_4329_2043# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X121 VDPWR VDPWR a_13186_4553# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X122 a_16486_16197# VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X123 a_23677_14701# ui_in[0] ui_in[1] VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.36 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=4316,272
X124 a_4905_12113# a_4627_12141# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X125 a_12823_4553# a_11439_4597# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X126 a_4915_10549# a_4637_10577# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X127 a_6087_14735# a_5809_14763# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X128 a_12793_14007# a_11147_11911# a_12697_14007# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X129 VGND VDPWR a_2313_2157# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X130 VGND a_14152_5441# a_14100_5467# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X131 VDPWR VGND a_17236_5473# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X132 a_7749_14003# a_7173_15235# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X133 VGND a_9317_5049# a_18371_4938# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=5796,222
X134 a_4213_5409# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X135 a_10121_1793# VDPWR a_10025_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X136 a_4383_1787# a_3199_1791# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X137 a_10289_4963# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X138 VDPWR VGND a_3010_1791# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X139 a_14432_4521# a_13709_4553# a_14657_4913# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X140 a_12615_14007# a_12039_15239# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X141 a_12227_2049# a_11175_1793# a_12644_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X142 VDPWR a_7944_1767# a_7892_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X143 a_4763_14525# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X144 a_16275_5839# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X145 a_17425_5473# a_16485_5729# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X146 a_24962_14701# ui_in[1] a_24234_14385# VGND sky130_fd_pr__nfet_01v8 ad=0.15102 pd=1.285 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=6041,257
X147 VGND VGND a_16994_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X148 VDPWR a_10132_5445# a_10080_5471# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X149 VGND VGND a_16539_5839# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X150 a_15188_4913# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X151 VGND VDPWR a_12587_5825# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X152 a_2259_2047# a_2187_1765# a_2676_1791# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X153 a_4746_2153# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X154 VGND VGND a_10553_4963# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X155 a_9503_10581# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X156 a_9781_10553# a_9503_10581# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X157 a_8337_2159# a_8283_2049# a_7944_1767# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X158 a_1950_5025# a_2217_5025# a_2175_5417# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X159 a_14179_2049# a_13167_1793# a_14596_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X160 a_10261_5471# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X161 a_10652_2159# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X162 a_15904_1767# a_15119_1793# a_16129_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X163 a_12865_14007# a_12039_15239# a_12793_14007# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X164 VDPWR VGND a_9461_14779# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X165 a_7749_14003# a_4915_10549# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=4368,272 d=2772,150
X166 VDPWR VGND a_10525_5471# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X167 VGND VDPWR a_14233_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X168 VDPWR a_9317_5049# a_18839_4938# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=6334,279
X169 a_3040_5051# VDPWR a_2289_5307# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X170 a_5895_14763# VGND a_5809_14763# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X171 a_8431_5415# a_7315_5043# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X172 VGND VDPWR a_4711_15373# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X173 VGND a_6281_11907# a_7749_14003# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2772,150 d=2268,138
X174 a_10499_4853# VDPWR a_10916_4597# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X175 a_6335_1787# a_5269_1787# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X176 VDPWR a_9896_1767# a_9844_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X177 VGND VDPWR a_6792_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X178 VGND VDPWR a_2676_2157# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X179 VGND VGND a_4513_14775# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X180 a_10717_13773# a_9703_16093# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X181 a_11810_13649# a_11195_12931# a_11728_13649# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X182 VGND VGND a_12281_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X183 a_16847_4529# a_16793_4785# a_16454_4503# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X184 a_16243_2049# a_15119_1793# a_16660_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X185 a_10025_1793# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X186 VGND VGND a_2313_2157# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X187 a_8193_13753# a_7749_14003# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5930,268 d=10800,508
X188 a_14152_5441# a_14419_5441# a_14377_5467# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X189 ua[0] a_24962_14701# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X190 a_4755_13107# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X191 a_12769_4809# a_11439_4597# a_13186_4919# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X192 VGND VDPWR a_9587_13813# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X193 a_9128_5049# VDPWR a_8377_5305# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X194 a_5933_13769# VGND a_5851_13769# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
X195 a_7032_2153# VDPWR a_6281_2043# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X196 VGND a_7113_13395# a_7749_14003# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2268,138 d=4075,198
X197 VGND a_9371_13111# a_9705_12861# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X198 a_10869_11939# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X199 VDPWR VDPWR a_12644_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X200 a_4765_11543# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X201 VGND VGND a_16847_4895# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X202 a_21506_16181# a_20384_16179# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X203 a_14561_4913# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X204 VGND VDPWR a_12823_4919# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X205 VDPWR VDPWR a_4840_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X206 VGND VGND a_12587_5825# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X207 a_3990_1761# a_3199_1791# a_4215_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X208 a_4503_16339# VDPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X209 VGND VGND a_14825_4913# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X210 VDPWR VDPWR a_16902_5473# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X211 a_8169_2159# VDPWR a_8073_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X212 VDPWR VGND a_3040_5051# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X213 VDPWR a_11255_13773# a_11810_13649# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5830,267
X214 a_2079_5417# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X215 a_3229_5051# a_2289_5307# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X216 VGND VDPWR a_14596_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X217 VGND sky130_fd_sc_hd__mux4_1_0.A3 a_2217_5025# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X218 VGND VDPWR a_4383_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X219 VGND VDPWR a_16660_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X220 a_11250_4963# VDPWR a_10499_4853# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X221 a_10132_5445# VGND a_10357_5837# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X222 a_2289_5307# a_2217_5025# a_2706_5051# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X223 ui_in[1] a_23731_14309# a_23677_14335# VGND sky130_fd_pr__nfet_01v8 ad=0.09322 pd=1.07 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3409,185
X224 a_6389_13769# a_5851_13769# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X225 VGND VGND a_14233_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X226 VDPWR a_4903_15345# a_5851_13769# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X227 VGND VGND a_2343_5417# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X228 VGND VDPWR a_10289_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X229 VDPWR VDPWR a_2343_5051# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X230 a_9451_16343# VDPWR a_9369_16343# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X231 a_10888_5837# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X232 a_9379_14779# VDPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X233 VGND VDPWR a_4723_10577# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X234 VGND VDPWR a_10525_5837# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X235 VDPWR VGND a_10986_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X236 VDPWR VDPWR a_9619_16343# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X237 a_4625_15373# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X238 a_10675_14767# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X239 a_9713_14529# VDPWR a_9629_14529# VGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X240 a_11222_5471# VDPWR a_10471_5727# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X241 a_19510_16177# a_18742_16187# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X242 a_9587_13813# VGND a_9501_13813# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X243 VGND VDPWR a_14908_5833# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X244 a_10553_4597# VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X245 a_14491_5723# a_14419_5441# a_14908_5833# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X246 VDPWR VGND a_9128_5049# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X247 a_9769_15349# a_9491_15377# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X248 VDPWR a_11979_13399# a_12865_14007# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=5930,268
X249 a_11175_1793# a_10235_2049# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X250 a_16793_4785# a_15711_4547# a_17210_4529# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X251 a_17733_4529# a_16793_4785# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X252 VGND a_10160_4571# a_10108_4597# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X253 a_24774_14701# ui_in[1] VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X254 a_16679_4529# VDPWR a_16583_4529# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X255 a_14657_4547# VDPWR a_14561_4547# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X256 a_9896_1767# a_9223_1793# a_10121_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X257 a_18742_16187# a_18128_16189# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X258 VDPWR VDPWR a_4635_13809# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X259 a_9317_5049# a_8377_5305# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X260 a_8431_5415# a_8377_5305# a_8038_5023# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X261 a_6281_2043# a_5269_1787# a_6698_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X262 a_6375_5299# a_5363_5043# a_6792_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X263 VGND VDPWR a_13186_4919# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X264 a_9705_12861# a_9371_13111# a_9621_13111# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X265 a_13167_1793# a_12227_2049# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X266 a_12823_4919# a_11439_4597# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X267 VDPWR sky130_fd_sc_hd__mux4_1_0.A1 a_23511_14701# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X268 a_11979_13399# a_11728_13649# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5830,267 d=13600,536
X269 a_6335_1787# a_6281_2043# a_5942_1761# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X270 VDPWR sky130_fd_sc_hd__mux4_1_0.A2 a_2187_1765# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X271 a_13709_4553# a_12769_4809# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X272 VDPWR a_22274_16171# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr d=10400,504
X273 ui_in[1] a_24774_14701# a_24962_14701# VGND sky130_fd_pr__nfet_01v8 ad=0.09322 pd=1.07 as=0.15102 ps=1.285 w=0.42 l=0.15
**devattr s=6041,257 d=4368,272
X274 a_6057_12927# VGND a_5975_12927# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X275 a_8700_2159# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X276 VGND VDPWR a_6335_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X277 VGND VGND a_17236_5839# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X278 a_3199_1791# a_2259_2047# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X279 VGND VGND a_11250_4963# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X280 a_23677_14335# VDPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X281 VDPWR VGND a_14545_5467# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X282 VGND VGND a_9371_13111# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X283 VDPWR a_9771_12117# a_10869_11939# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X284 a_4119_2153# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X285 a_12655_4553# VDPWR a_12559_4553# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X286 VGND a_6389_13769# a_6862_13645# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4010,197
X287 a_18625_5265# a_18371_4938# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=5796,222 d=2772,150
X288 a_12281_1793# a_11175_1793# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X289 a_8337_2159# a_7221_1787# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X290 a_17544_4895# VDPWR a_16793_4785# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X291 a_4477_5043# a_3229_5051# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X292 a_9619_16343# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X293 a_9629_14529# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X294 VDPWR VGND a_11222_5471# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X295 a_2313_1791# a_2187_1765# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X296 a_5975_12927# a_4913_13781# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0805 pd=0.94333 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2646,147
X297 a_13284_5825# VDPWR a_12533_5715# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X298 VGND VGND a_4383_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X299 a_10916_4963# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X300 VDPWR VDPWR a_2706_5051# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X301 a_15522_4913# VDPWR a_14771_4803# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X302 VGND VDPWR a_10553_4963# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X303 VGND a_4837_16089# a_6911_15235# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X304 VGND VGND a_10289_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X305 a_11195_12931# a_10841_12931# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5689,267 d=10400,504
X306 a_10261_5837# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X307 a_11411_5471# a_10471_5727# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X308 a_9463_11547# VDPWR a_9381_11547# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X309 VGND VGND a_10525_5837# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X310 a_4847_14525# VDPWR a_4763_14525# VGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X311 VDPWR VDPWR a_9631_11547# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X312 a_9034_1793# VDPWR a_8283_2049# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X313 VGND a_14432_4521# a_14380_4547# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X314 a_15119_1793# a_14179_2049# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X315 VGND a_16454_4503# a_16402_4529# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X316 a_3040_5417# VDPWR a_2289_5307# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X317 VDPWR VDPWR a_12950_5459# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X318 a_14545_5833# a_14419_5441# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X319 sky130_fd_sc_hd__mux4_1_0.A2 a_16243_2049# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X320 VDPWR VDPWR a_17210_4529# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X321 VDPWR VDPWR a_15188_4547# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X322 a_4713_12141# VGND a_4627_12141# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X323 a_12587_5459# a_11411_5471# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X324 a_10121_2159# VDPWR a_10025_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X325 a_16847_4529# a_15711_4547# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X326 VGND a_6036_5017# a_5984_5043# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X327 a_6792_5043# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X328 VGND VGND a_3010_2157# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X329 a_12227_2049# a_11175_1793# a_12644_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X330 a_6717_15235# a_6629_15387# a_6635_15235# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
X331 a_8263_5415# VDPWR a_8167_5415# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X332 VDPWR VDPWR a_10652_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X333 a_4837_16089# a_4503_16339# a_4753_16339# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X334 a_14233_1793# a_13167_1793# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X335 a_6071_2153# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X336 a_6429_5043# a_5363_5043# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X337 VGND VGND a_17544_4895# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X338 VDPWR VDPWR a_8794_5049# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X339 a_16297_1793# a_15119_1793# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X340 a_6167_1787# VDPWR a_6071_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X341 a_2259_2047# a_2187_1765# a_2676_2157# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X342 VGND a_12430_4527# a_12378_4553# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X343 VGND a_9379_14779# a_9713_14529# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X344 a_10553_4597# a_10499_4853# a_10160_4571# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X345 a_4753_16089# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X346 VDPWR VGND a_5975_12927# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0805 ps=0.94333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X347 VGND VGND a_6335_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X348 VGND a_4839_12857# a_5895_14763# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X349 VGND VGND a_13284_5825# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X350 VGND VGND a_15522_4913# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X351 VDPWR VGND a_8431_5049# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X352 a_12039_15239# a_11501_15239# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X353 a_16454_4503# a_15711_4547# a_16679_4895# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X354 a_18128_16189# a_17254_16187# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X355 a_9771_12117# a_9493_12145# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X356 a_17210_4895# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X357 VDPWR VDPWR a_9493_12145# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X358 VGND VDPWR a_4840_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X359 VGND VDPWR a_10916_4963# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X360 a_12194_5433# a_11411_5471# a_12419_5825# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X361 a_15242_5467# VDPWR a_14491_5723# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X362 sky130_fd_sc_hd__mux4_1_0.A1 a_12615_14007# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4075,198 d=7020,368
X363 a_12950_5825# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X364 VGND sky130_fd_sc_hd__mux4_1_0.A1 a_6629_15387# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X365 VGND VDPWR a_16902_5839# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X366 VGND VGND a_3040_5417# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X367 VGND a_4505_13107# a_4839_12857# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X368 a_10953_14739# a_10675_14767# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X369 VDPWR VDPWR a_4755_13107# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X370 a_4477_5043# a_4423_5299# a_4084_5017# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X371 a_4905_12113# a_4627_12141# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X372 a_2289_5307# a_2217_5025# a_2706_5417# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X373 a_7944_1767# a_7221_1787# a_8169_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X374 a_5080_2153# VDPWR a_4329_2043# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X375 VDPWR sky130_fd_sc_hd__mux4_1_0.A3 a_24407_14651# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.09013 ps=0.995 w=0.42 l=0.15
**devattr s=3605,199 d=2268,138
X376 VDPWR VDPWR a_4765_11543# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X377 VDPWR VDPWR a_10888_5471# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X378 VDPWR a_15904_1767# a_15852_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X379 a_16539_5473# a_16485_5729# a_16146_5447# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X380 a_10471_5727# VGND a_10888_5471# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X381 a_16243_2049# a_15119_1793# a_16660_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X382 VDPWR VDPWR a_8337_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X383 a_13969_1793# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X384 a_10025_2159# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X385 VGND VGND a_4503_16339# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X386 VGND VDPWR a_2343_5417# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X387 a_8794_5415# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X388 a_7221_1787# a_6281_2043# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X389 a_9621_13111# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X390 a_11222_5837# VDPWR a_10471_5727# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X391 VGND VDPWR a_12644_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X392 a_6698_1787# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X393 a_20384_16179# a_19510_16177# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X394 sky130_fd_sc_hd__mux4_1_0.A3 a_18625_4938# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4514,209 d=6760,364
X395 a_9493_12145# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X396 a_17254_16187# a_16486_16197# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X397 VGND VDPWR a_9577_15377# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X398 a_6862_13645# a_6329_12927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X399 a_12587_5459# a_12533_5715# a_12194_5433# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X400 a_10385_4597# VDPWR a_10289_4597# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X401 a_14825_4547# a_14771_4803# a_14432_4521# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X402 VDPWR VGND a_15242_5467# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X403 a_5851_13769# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X404 a_4721_13809# VGND a_4635_13809# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X405 a_6375_5299# a_5363_5043# a_6792_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X406 a_14545_5833# a_14491_5723# a_14152_5441# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X407 VDPWR VGND a_9451_16343# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X408 VDPWR a_4847_14525# a_6635_15235# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X409 VGND VGND a_9379_14779# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X410 VDPWR a_9705_12861# a_10675_14767# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X411 a_16583_4895# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X412 VDPWR VDPWR a_4625_15373# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X413 a_6429_5043# a_6375_5299# a_6036_5017# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X414 a_15431_5467# a_14491_5723# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X415 a_16297_1793# a_16243_2049# a_15904_1767# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X416 a_14233_1793# a_14179_2049# a_13840_1767# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X417 VGND VGND a_5080_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X418 a_7113_13395# a_6862_13645# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5830,267 d=13600,536
X419 a_12323_5825# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X420 a_12978_1793# VDPWR a_12227_2049# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X421 a_14908_5467# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X422 a_12655_4919# VDPWR a_12559_4919# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X423 VDPWR VDPWR a_14545_5467# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X424 a_12823_4553# a_12769_4809# a_12430_4527# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X425 VGND VGND a_10986_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X426 a_14771_4803# a_13709_4553# a_15188_4913# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X427 a_9631_11547# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X428 a_4477_5409# a_3229_5051# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X429 a_4329_2043# a_3199_1791# a_4746_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X430 a_11255_13773# a_10717_13773# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X431 a_5363_5043# a_4423_5299# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X432 a_4423_5299# a_3229_5051# a_4840_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X433 a_24774_14701# ui_in[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X434 a_4309_5043# VDPWR a_4213_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X435 VGND VGND a_11222_5837# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X436 a_23677_14701# VDPWR VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.36 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X437 a_8073_1793# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X438 a_4383_1787# a_4329_2043# a_3990_1761# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X439 VGND VDPWR a_14825_4913# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X440 a_16485_5729# a_15431_5467# a_16902_5473# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X441 VGND VGND a_4505_13107# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X442 VGND VDPWR a_2706_5417# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X443 a_9896_1767# a_9223_1793# a_10121_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X444 VDPWR a_5942_1761# a_5890_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X445 VGND a_9317_5049# a_18846_5265# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=4514,209
X446 a_9577_15377# VGND a_9491_15377# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X447 a_10993_13773# a_9703_16093# a_10887_13773# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X448 VDPWR VGND a_8337_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X449 ua[0] a_24962_14701# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X450 a_2145_1791# VDPWR a_2049_1791# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X451 a_8038_5023# a_7315_5043# a_8263_5415# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X452 a_10525_5471# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X453 a_5809_14763# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X454 VGND VDPWR a_8431_5415# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X455 VDPWR VGND a_16847_4529# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X456 a_5942_1761# a_5269_1787# a_6167_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X457 VDPWR a_4837_16089# a_6635_15235# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X458 a_13473_5459# a_12533_5715# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X459 a_12533_5715# a_11411_5471# a_12950_5459# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X460 VGND VGND a_7032_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X461 a_15711_4547# a_14771_4803# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X462 a_12559_4553# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X463 a_6792_5409# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X464 a_12419_5459# VDPWR a_12323_5459# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X465 a_12281_2159# a_11175_1793# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X466 a_14377_5833# VDPWR a_14281_5833# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X467 VDPWR a_14152_5441# a_14100_5467# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X468 a_10235_2049# a_9223_1793# a_10652_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X469 a_14930_1793# VDPWR a_14179_2049# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X470 a_16994_1793# VDPWR a_16243_2049# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X471 VDPWR VGND a_9463_11547# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X472 a_6429_5409# a_5363_5043# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X473 a_7315_5043# a_6375_5299# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X474 a_2313_2157# a_2187_1765# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X475 VDPWR VDPWR a_9501_13813# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X476 a_14065_1793# VDPWR a_13969_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X477 a_16129_1793# VDPWR a_16033_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X478 a_22274_16171# a_21506_16181# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X479 a_4505_13107# VDPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X480 a_14281_5467# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X481 VGND a_7944_1767# a_7892_1793# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X482 a_6635_15235# a_6629_15387# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X483 VGND VDPWR a_4713_12141# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X484 a_6261_5043# VDPWR a_6165_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X485 VGND VGND a_4515_11543# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X486 VGND a_4084_5017# a_4032_5043# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X487 a_4840_5043# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X488 VGND a_16146_5447# a_16094_5473# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X489 a_9034_2159# VDPWR a_8283_2049# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X490 a_9769_15349# a_9491_15377# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X491 VGND VDPWR a_4746_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X492 a_14825_4913# a_13709_4553# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X493 a_2676_1791# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X494 a_11671_15239# a_9713_14529# a_11583_15239# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X495 a_9779_13785# a_9501_13813# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X496 a_4215_1787# VDPWR a_4119_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X497 a_11195_12931# a_10841_12931# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=5266,228 d=6760,364
X498 a_4837_16089# VDPWR a_4753_16089# VGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X499 a_16539_5473# a_15431_5467# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X500 a_4913_13781# a_4635_13809# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X501 VDPWR a_4839_12857# a_5975_12927# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0805 ps=0.94333 w=0.42 l=0.15
**devattr s=2646,147 d=5689,267
X502 a_6329_12927# a_5975_12927# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5689,267 d=10400,504
X503 VGND a_1950_5025# a_1898_5051# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X504 a_8167_5415# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X505 VGND VDPWR a_10652_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X506 a_4477_5409# a_4423_5299# a_4084_5017# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X507 a_14233_2159# a_13167_1793# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X508 VGND VDPWR a_10888_5837# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X509 a_16539_5839# a_16485_5729# a_16146_5447# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X510 a_11439_4597# a_10499_4853# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X511 a_24234_14385# ui_in[0] a_24241_14651# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1274 pd=1.16667 as=0.10855 ps=1.36 w=0.42 l=0.15
**devattr s=4316,272 d=2268,138
X512 a_16297_2159# a_15119_1793# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X513 a_6281_11907# a_6003_11935# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X514 a_10955_11939# VGND a_10869_11939# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X515 a_10471_5727# VGND a_10888_5837# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X516 VGND a_12194_5433# a_12142_5459# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X517 a_18553_4938# a_18371_4938# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X518 a_10160_4571# VDPWR a_10385_4597# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X519 VDPWR a_4905_12113# a_6003_11935# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X520 a_9501_13813# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X521 a_4847_14525# a_4513_14775# a_4763_14775# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X522 a_11147_11911# a_10869_11939# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X523 VGND a_9896_1767# a_9844_1793# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X524 a_4515_11543# VDPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X525 VDPWR VGND a_10841_12931# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0805 ps=0.94333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X526 a_17544_4529# VDPWR a_16793_4785# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X527 VDPWR a_11888_1767# a_11836_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X528 a_14596_1793# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X529 a_16660_1793# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X530 a_24241_14651# sky130_fd_sc_hd__mux4_1_0.A2 VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.36 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X531 a_12017_1793# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X532 VGND VDPWR a_6698_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X533 a_9453_13111# VDPWR a_9371_13111# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X534 a_6021_13769# a_4903_15345# a_5933_13769# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X535 VDPWR a_1920_1765# a_1868_1791# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X536 a_11501_15239# a_10953_14739# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X537 VGND sky130_fd_sc_hd__mux4_1_0.A3 a_24152_14385# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.10855 ps=1.36 w=0.42 l=0.15
**devattr s=4316,272 d=2268,138
X538 a_6127_13769# a_4837_16089# a_6021_13769# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X539 VDPWR VDPWR a_9621_13111# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X540 a_4627_12141# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X541 a_8377_5305# a_7315_5043# a_8794_5049# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X542 a_9713_14529# a_9379_14779# a_9629_14779# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X543 a_6429_5409# a_6375_5299# a_6036_5017# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X544 a_7944_1767# a_7221_1787# a_8169_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X545 a_10887_13773# a_9769_15349# a_10799_13773# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X546 a_4746_1787# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X547 a_10761_14767# VGND a_10675_14767# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X548 a_4637_10577# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X549 VDPWR sky130_fd_sc_hd__mux4_1_0.A3 a_2217_5025# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X550 VDPWR VDPWR a_12281_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X551 VGND VDPWR a_8337_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X552 a_13969_2159# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X553 VGND ui_in[0] a_23731_14309# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X554 a_6003_11935# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X555 VDPWR VDPWR a_4477_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X556 VDPWR VGND a_9034_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X557 a_12823_4919# a_12769_4809# a_12430_4527# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X558 a_7831_14003# a_4915_10549# a_7749_14003# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2772,150
X559 a_16486_16197# VDPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X560 VGND VDPWR a_4721_13809# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X561 a_4423_5299# a_3229_5051# a_4840_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X562 a_4383_2153# a_3199_1791# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X563 a_10499_4853# VDPWR a_10916_4963# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X564 a_4309_5409# VDPWR a_4213_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X565 a_16485_5729# a_15431_5467# a_16902_5839# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X566 a_9223_1793# a_8283_2049# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X567 VDPWR VGND a_17544_4529# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X568 a_12281_1793# a_12227_2049# a_11888_1767# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X569 a_2343_5051# a_2217_5025# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X570 a_7927_14003# a_6281_11907# a_7831_14003# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X571 a_10289_4597# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X572 a_7173_15235# a_6635_15235# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X573 a_12039_15239# a_11501_15239# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X574 a_10525_5837# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X575 VDPWR a_13840_1767# a_13788_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X576 a_8283_2049# a_7221_1787# a_8700_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X577 a_14432_4521# a_13709_4553# a_14657_4547# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X578 a_24234_14385# a_24774_14701# a_24962_14701# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1274 pd=1.16667 as=0.09209 ps=0.99 w=0.42 l=0.15
**devattr s=3683,198 d=10752,424
X579 a_14152_5441# a_14419_5441# a_14377_5833# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X580 a_2313_1791# a_2259_2047# a_1920_1765# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X581 a_17733_4529# a_16793_4785# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X582 a_9771_12117# a_9493_12145# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X583 VGND a_9771_12117# a_10955_11939# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X584 a_16454_4503# a_15711_4547# a_16679_4529# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X585 a_9128_5415# VDPWR a_8377_5305# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X586 a_11777_15239# a_10953_14739# a_11671_15239# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X587 a_17210_4529# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X588 a_15188_4547# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X589 VDPWR a_9705_12861# a_10717_13773# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X590 a_10357_5471# VDPWR a_10261_5471# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X591 VDPWR VDPWR a_12587_5459# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X592 a_11175_1793# a_10235_2049# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X593 VDPWR VGND a_10553_4597# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X594 a_9781_10553# a_9503_10581# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X595 a_14233_2159# a_14179_2049# a_13840_1767# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X596 a_16297_2159# a_16243_2049# a_15904_1767# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X597 a_13840_1767# a_13167_1793# a_14065_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X598 a_8193_13753# a_7749_14003# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4075,198 d=7020,368
X599 a_4755_12857# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X600 a_12978_2159# VDPWR a_12227_2049# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X601 VGND a_4515_11543# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr d=10010,284
X602 a_6036_5017# a_5363_5043# a_6261_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X603 VDPWR a_9705_12861# a_10841_12931# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0805 ps=0.94333 w=0.42 l=0.15
**devattr s=2646,147 d=5689,267
X604 a_13709_4553# a_12769_4809# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X605 a_12559_4919# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X606 VDPWR a_3990_1761# a_3938_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X607 a_4585_16339# VDPWR a_4503_16339# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X608 a_12430_4527# a_11439_4597# a_12655_4553# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X609 a_10953_14739# a_10675_14767# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X610 VDPWR a_7113_13395# a_7999_14003# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=5930,268
X611 VGND a_8038_5023# a_7986_5049# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X612 VDPWR VDPWR a_6429_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X613 a_7032_1787# VDPWR a_6281_2043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X614 VDPWR VDPWR a_16297_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X615 a_10289_1793# a_9223_1793# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X616 VDPWR a_4839_12857# a_5809_14763# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X617 a_6335_2153# a_5269_1787# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X618 a_4595_14775# VDPWR a_4513_14775# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X619 a_7999_14003# a_7173_15235# a_7927_14003# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X620 a_5269_1787# a_4329_2043# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X621 a_8073_2159# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X622 a_13186_4553# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X623 a_3990_1761# a_3199_1791# a_4215_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X624 a_8431_5049# a_7315_5043# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X625 VGND VGND a_8337_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X626 a_18846_5265# a_17733_4529# a_18625_4938# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
**devattr s=3990,179 d=2772,150
X627 a_6261_5409# VDPWR a_6165_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X628 a_2049_1791# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X629 a_2145_2157# VDPWR a_2049_2157# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X630 a_4840_5409# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X631 VDPWR VGND a_4477_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X632 VDPWR VDPWR a_4383_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X633 a_6389_13769# a_5851_13769# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X634 a_4839_12857# a_4505_13107# a_4755_13107# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X635 VGND VDPWR a_16847_4895# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X636 a_10553_4963# VDPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X637 a_19510_16177# a_18742_16187# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X638 VGND a_4839_12857# a_6127_13769# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X639 VDPWR a_9769_15349# a_10717_13773# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X640 VGND VGND a_9128_5415# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X641 a_16539_5839# a_15431_5467# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X642 a_12113_1793# VDPWR a_12017_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X643 a_3010_1791# VDPWR a_2259_2047# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X644 VGND a_9705_12861# a_10993_13773# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X645 VDPWR a_16454_4503# a_16402_4529# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X646 VDPWR a_14432_4521# a_14380_4547# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X647 a_14657_4913# VDPWR a_14561_4913# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X648 a_17425_5473# a_16485_5729# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X649 a_23511_14335# ui_in[0] ui_in[1] VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.09322 ps=1.07 w=0.42 l=0.15
**devattr s=3409,185 d=4368,272
X650 VDPWR VDPWR a_8700_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X651 a_4765_11293# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X652 VGND a_10132_5445# a_10080_5471# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X653 a_21506_16181# a_20384_16179# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X654 a_14930_2159# VDPWR a_14179_2049# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X655 a_16994_2159# VDPWR a_16243_2049# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X656 a_10235_2049# a_9223_1793# a_10652_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X657 a_16583_4529# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X658 a_14561_4547# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X659 a_16371_5473# VDPWR a_16275_5473# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X660 a_4903_15345# a_4625_15373# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X661 VDPWR a_6036_5017# a_5984_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X662 VDPWR VGND a_12587_5459# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X663 a_14065_2159# VDPWR a_13969_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X664 a_16129_2159# VDPWR a_16033_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X665 VDPWR VGND a_14825_4547# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X666 VGND a_11255_13773# a_11728_13649# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4010,197
X667 a_6165_5043# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X668 VGND VGND a_14545_5833# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X669 a_2343_5051# a_2289_5307# a_1950_5025# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X670 a_16033_1793# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X671 a_6281_2043# a_5269_1787# a_6698_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X672 VDPWR a_12430_4527# a_12378_4553# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X673 VDPWR VGND a_6429_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X674 VDPWR a_6389_13769# a_6944_13645# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5830,267
X675 VDPWR VGND a_16297_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X676 a_11250_4597# VDPWR a_10499_4853# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X677 VDPWR VDPWR a_6335_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X678 a_24407_14651# a_23731_14309# a_24234_14385# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.09013 pd=0.995 as=0.1274 ps=1.16667 w=0.42 l=0.15
**devattr s=2268,138 d=3605,199
X679 VGND a_4839_12857# a_6129_12927# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5266,228
X680 a_2676_2157# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X681 a_4119_1787# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X682 a_9369_16343# VDPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X683 VGND a_9703_16093# a_11777_15239# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X684 VDPWR VGND a_12823_4553# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X685 a_9703_16093# VDPWR a_9619_16093# VGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X686 VGND a_9705_12861# a_10995_12931# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5266,228
X687 a_10289_1793# a_10235_2049# a_9896_1767# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X688 VDPWR VDPWR a_14908_5467# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X689 a_10841_12931# a_9779_13785# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0805 pd=0.94333 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2646,147
X690 VDPWR VGND a_4383_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X691 a_14491_5723# a_14419_5441# a_14908_5467# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X692 a_12644_1793# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X693 VDPWR a_9317_5049# a_18371_4938# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2772,150
X694 a_18742_16187# a_18128_16189# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X695 a_6335_2153# a_6281_2043# a_5942_1761# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X696 VGND VDPWR a_9579_12145# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X697 a_6329_12927# a_5975_12927# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=5266,228 d=6760,364
X698 VGND VDPWR a_4477_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X699 VGND VDPWR a_12950_5825# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X700 a_5174_5043# VDPWR a_4423_5299# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X701 VGND VDPWR a_15188_4913# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X702 a_8431_5049# a_8377_5305# a_8038_5023# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X703 a_11583_15239# a_8193_13753# a_11501_15239# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
X704 a_11728_13649# a_11195_12931# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X705 a_12587_5825# a_11411_5471# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X706 VGND VDPWR a_9589_10581# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X707 a_17236_5473# VDPWR a_16485_5729# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X708 VDPWR a_22274_16171# VGND VGND sky130_fd_pr__nfet_01v8 ad=9.689 pd=135.58 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X709 a_11979_13399# a_11728_13649# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4010,197 d=6760,364
X710 VDPWR VGND a_9453_13111# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X711 a_24318_14385# sky130_fd_sc_hd__mux4_1_0.A2 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10858 pd=1.36 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X712 a_10717_13773# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X713 a_10923_12931# VGND a_10841_12931# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X714 a_14596_2159# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X715 VGND a_15904_1767# a_15852_1793# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X716 a_16660_2159# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X717 VDPWR VDPWR a_4627_12141# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X718 a_6281_11907# a_6003_11935# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X719 VGND a_9705_12861# a_10761_14767# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X720 a_4915_10549# a_4637_10577# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X721 a_2343_5417# a_2217_5025# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X722 VGND VDPWR a_8794_5415# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X723 VDPWR VGND a_11250_4597# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X724 a_24318_14385# a_23731_14309# a_24234_14385# VGND sky130_fd_pr__nfet_01v8 ad=0.10858 pd=1.36 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=4318,272
X725 a_12615_14007# a_9781_10553# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=4368,272 d=2772,150
X726 a_11147_11911# a_10869_11939# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X727 a_3229_5051# a_2289_5307# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X728 a_6087_14735# a_5809_14763# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X729 VDPWR VDPWR a_4637_10577# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X730 a_10553_4963# a_10499_4853# a_10160_4571# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X731 a_12017_2159# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X732 VDPWR VGND a_14930_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X733 a_4753_16339# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X734 a_9619_16093# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X735 VGND VGND a_8431_5415# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X736 a_2175_5051# VDPWR a_2079_5051# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X737 a_6071_1787# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X738 a_4763_14775# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X739 a_10357_5837# VDPWR a_10261_5837# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X740 a_13284_5459# VDPWR a_12533_5715# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X741 a_10916_4597# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X742 VDPWR VGND a_6335_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X743 a_15522_4547# VDPWR a_14771_4803# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X744 a_18128_16189# a_17254_16187# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X745 a_10525_5471# a_10471_5727# a_10132_5445# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X746 VDPWR VDPWR a_10553_4597# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X747 VGND VDPWR a_12281_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X748 a_6036_5017# a_5363_5043# a_6261_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X749 a_15242_5833# VDPWR a_14491_5723# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X750 a_10995_12931# a_9779_13785# a_10923_12931# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=1764,126
X751 a_9579_12145# VGND a_9493_12145# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X752 a_9381_11547# VDPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X753 a_10986_1793# VDPWR a_10235_2049# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X754 VDPWR VGND a_12978_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X755 VGND VGND a_9034_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X756 a_12430_4527# a_11439_4597# a_12655_4919# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X757 VGND VDPWR a_6429_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X758 a_7126_5043# VDPWR a_6375_5299# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X759 VGND VDPWR a_9631_11297# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X760 a_9589_10581# VGND a_9503_10581# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X761 VDPWR VGND a_5174_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X762 a_13167_1793# a_12227_2049# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X763 a_13186_4919# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X764 a_9317_5049# a_8377_5305# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X765 a_14545_5467# a_14419_5441# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X766 a_12281_2159# a_12227_2049# a_11888_1767# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X767 a_11888_1767# a_11175_1793# a_12113_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X768 a_13520_4553# VDPWR a_12769_4809# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X769 a_10799_13773# VGND a_10717_13773# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
X770 a_5363_5043# a_4423_5299# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X771 a_6167_2153# VDPWR a_6071_2153# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X772 a_4839_12857# VDPWR a_4755_12857# VGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X773 a_4084_5017# a_3229_5051# a_4309_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X774 a_8283_2049# a_7221_1787# a_8700_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X775 a_3199_1791# a_2259_2047# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X776 VGND VGND a_4477_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X777 a_2313_2157# a_2259_2047# a_1920_1765# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X778 a_8263_5049# VDPWR a_8167_5049# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X779 VDPWR ui_in[0] a_23731_14309# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.1083 ps=1.36 w=0.42 l=0.15
**devattr s=4332,272 d=4316,272
X780 a_1920_1765# a_2187_1765# a_2145_1791# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X781 VDPWR VGND a_4585_16339# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X782 a_5080_1787# VDPWR a_4329_2043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X783 a_16146_5447# a_15431_5467# a_16371_5473# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X784 VGND a_9369_16343# a_9703_16093# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X785 a_16902_5473# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X786 VDPWR VGND a_4595_14775# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X787 a_13840_1767# a_13167_1793# a_14065_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X788 VDPWR VDPWR a_16539_5473# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X789 VGND a_5942_1761# a_5890_1787# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X790 a_16847_4895# a_16793_4785# a_16454_4503# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X791 VDPWR VGND a_13284_5459# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X792 VDPWR VDPWR a_2313_1791# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X793 a_9621_12861# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X794 VDPWR VGND a_15522_4547# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X795 a_2706_5051# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X796 a_12587_5825# a_12533_5715# a_12194_5433# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X797 VDPWR a_10160_4571# a_10108_4597# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X798 a_10385_4963# VDPWR a_10289_4963# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X799 a_17254_16187# a_16486_16197# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X800 VDPWR a_9713_14529# a_11501_15239# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X801 VGND VGND a_15242_5833# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X802 a_14825_4913# a_14771_4803# a_14432_4521# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X803 sky130_fd_sc_hd__mux4_1_0.A1 a_12615_14007# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5930,268 d=10800,508
X804 a_6635_15235# a_6087_14735# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X805 VGND VDPWR a_16297_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X806 a_9703_16093# a_9369_16343# a_9619_16343# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X807 a_13473_5459# a_12533_5715# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X808 a_16371_5839# VDPWR a_16275_5839# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X809 a_10289_2159# a_9223_1793# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X810 ui_in[1] a_23731_14309# a_23511_14701# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X811 a_18839_4938# a_17425_5473# a_18625_4938# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
**devattr s=7728,268 d=3066,157
X812 a_15711_4547# a_14771_4803# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X813 VDPWR VDPWR a_10916_4597# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X814 VDPWR VGND a_7126_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X815 a_12194_5433# a_11411_5471# a_12419_5459# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X816 VDPWR VGND a_16994_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X817 a_12950_5459# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X818 a_11411_5471# a_10471_5727# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X819 a_15119_1793# a_14179_2049# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X820 a_24962_14701# ui_in[1] ui_in[1] VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.09209 pd=0.99 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=3683,198
X821 a_8337_1793# a_8283_2049# a_7944_1767# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X822 a_6165_5409# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X823 a_7315_5043# a_6375_5299# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X824 a_14908_5833# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X825 a_2049_2157# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X826 a_2343_5417# a_2289_5307# a_1950_5025# VGND sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X827 sky130_fd_sc_hd__mux4_1_0.A2 a_16243_2049# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20731 ps=2.00287 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X828 VDPWR VGND a_13520_4553# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X829 VGND a_11147_11911# a_12615_14007# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2772,150 d=2268,138
X830 VGND VDPWR a_14545_5833# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X831 a_10652_1793# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X832 a_14179_2049# a_13167_1793# a_14596_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X833 VGND sky130_fd_sc_hd__mux4_1_0.A2 a_2187_1765# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X834 VGND VGND a_6429_5409# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X835 a_15904_1767# a_15119_1793# a_16129_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X836 a_11439_4597# a_10499_4853# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X837 VGND VDPWR a_4765_11293# VGND sky130_fd_pr__nfet_01v8 ad=0.13063 pd=1.32737 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X838 VDPWR a_4084_5017# a_4032_5043# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X839 VDPWR VDPWR a_14233_1793# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X840 VDPWR VGND a_5080_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X841 a_6698_2153# VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.08441 ps=0.85768 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X842 a_12113_2159# VDPWR a_12017_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X843 a_3010_2157# VDPWR a_2259_2047# VGND sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X844 VGND VGND a_12823_4919# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X845 a_8794_5049# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X846 a_7173_15235# a_6635_15235# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X847 VDPWR a_16146_5447# a_16094_5473# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X848 a_5851_13769# a_4837_16089# VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X849 VGND a_4515_11543# a_4765_11543# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=3.156 pd=47.08 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X850 VGND a_4905_12113# a_6089_11935# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X851 VGND VDPWR a_8700_2159# VGND sky130_fd_pr__nfet_01v8 ad=0.08441 pd=0.85768 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X852 a_4213_5043# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X853 a_4329_2043# a_3199_1791# a_4746_1787# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X854 a_9461_14779# VDPWR a_9379_14779# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X855 a_20384_16179# a_19510_16177# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13063 ps=1.32737 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X856 a_6911_15235# a_6087_14735# a_6805_15235# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X857 VDPWR a_4839_12857# a_5851_13769# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X858 a_16275_5473# VGND VDPWR VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08707 ps=0.84121 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X859 VDPWR VDPWR a_9629_14779# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X860 VDPWR a_1950_5025# a_1898_5051# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.20731 pd=2.00287 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X861 VDPWR VDPWR a_2676_1791# VDPWR sky130_fd_pr__pfet_01v8_hvt ad=0.08707 pd=0.84121 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
C0 a_10499_4853# a_11439_4597# 0.14008f
C1 a_14491_5723# a_14377_5833# 0
C2 a_24774_14701# sky130_fd_sc_hd__mux4_1_0.A3 0
C3 VDPWR a_10652_2159# 0.02101f
C4 a_2259_2047# a_2676_2157# 0.06611f
C5 a_14491_5723# a_14545_5833# 0.03622f
C6 a_10953_14739# a_11728_13649# 0
C7 a_12378_4553# a_12559_4919# 0
C8 a_15431_5467# a_14491_5723# 0.13739f
C9 a_11411_5471# sky130_fd_sc_hd__mux4_1_0.A3 0.00685f
C10 a_9317_5049# a_9128_5415# 0
C11 a_16146_5447# a_16539_5473# 0.02283f
C12 a_11501_15239# a_11728_13649# 0
C13 a_9501_13813# a_8193_13753# 0.00137f
C14 VDPWR a_8794_5415# 0.02123f
C15 a_12378_4553# a_11439_4597# 0.04873f
C16 a_15119_1793# a_16660_2159# 0.03325f
C17 a_3010_2157# a_2259_2047# 0.00696f
C18 a_11255_13773# a_11979_13399# 0.0615f
C19 a_10953_14739# a_10675_14767# 0.1109f
C20 a_11810_13649# a_9705_12861# 0
C21 a_6792_5409# a_6375_5299# 0.06611f
C22 a_16146_5447# a_15711_4547# 0
C23 a_9705_12861# a_10799_13773# 0
C24 sky130_fd_sc_hd__mux4_1_0.A2 ua[0] 0
C25 a_18742_16187# a_18128_16189# 0.10376f
C26 a_10499_4853# a_11411_5471# 0
C27 a_9705_12861# a_10923_12931# 0.00148f
C28 VDPWR a_1950_5025# 0.36083f
C29 a_16486_16197# sky130_fd_sc_hd__mux4_1_0.A1 0
C30 VDPWR a_10357_5837# 0
C31 a_14233_1793# a_14179_2049# 0.00386f
C32 a_9491_15377# a_9379_14779# 0
C33 a_11728_13649# a_9703_16093# 0
C34 a_14377_5467# a_14545_5467# 0
C35 a_13840_1767# a_14065_1793# 0.00487f
C36 a_11255_13773# a_10717_13773# 0.07901f
C37 VDPWR a_9369_16343# 0.5106f
C38 a_6635_15235# a_6087_14735# 0.08698f
C39 a_10235_2049# a_11836_1793# 0
C40 VDPWR a_7113_13395# 0.50533f
C41 a_14179_2049# a_14930_2159# 0.00696f
C42 a_9781_10553# a_11728_13649# 0
C43 a_14281_5833# a_14545_5833# 0
C44 VDPWR a_12419_5825# 0
C45 a_10675_14767# a_9703_16093# 0.03093f
C46 a_6129_12927# a_4913_13781# 0
C47 a_4635_13809# a_4513_14775# 0.00144f
C48 a_4839_12857# a_6862_13645# 0.00327f
C49 a_7986_5049# sky130_fd_sc_hd__mux4_1_0.A3 0.00121f
C50 a_16539_5839# a_16485_5729# 0.03622f
C51 VDPWR a_12793_14007# 0
C52 VDPWR a_5975_12927# 0.22891f
C53 a_13167_1793# a_14065_1793# 0
C54 a_8169_1793# a_8283_2049# 0
C55 a_6087_14735# a_7173_15235# 0.00407f
C56 a_10235_2049# a_10652_2159# 0.06611f
C57 sky130_fd_sc_hd__mux4_1_0.A2 a_9844_1793# 0.00121f
C58 a_13840_1767# a_14065_2159# 0.00559f
C59 a_13473_5459# a_13284_5825# 0
C60 a_4625_15373# a_4753_16339# 0
C61 a_9317_5049# a_17210_4895# 0
C62 VDPWR a_16371_5839# 0
C63 a_6036_5017# a_6165_5409# 0.00792f
C64 a_4505_13107# a_6329_12927# 0
C65 a_11147_11911# a_9781_10553# 0.43338f
C66 a_15904_1767# a_16129_2159# 0.00559f
C67 VDPWR a_12615_14007# 0.13215f
C68 a_18625_4938# sky130_fd_sc_hd__mux4_1_0.A3 0.10138f
C69 a_16902_5473# a_15431_5467# 0.08907f
C70 a_14596_1793# a_13167_1793# 0.08907f
C71 a_9779_13785# a_10993_13773# 0
C72 a_2145_2157# a_2187_1765# 0
C73 a_10357_5471# a_10471_5727# 0
C74 a_4913_13781# a_6087_14735# 0
C75 a_14377_5467# a_14152_5441# 0.00487f
C76 a_14377_5467# a_13473_5459# 0
C77 a_6429_5043# a_6036_5017# 0.02283f
C78 a_12587_5825# a_11439_4597# 0
C79 a_4903_15345# a_4847_14525# 0.15227f
C80 a_4505_13107# a_4635_13809# 0.00115f
C81 VDPWR a_14491_5723# 0.45311f
C82 a_4477_5409# a_4084_5017# 0.02301f
C83 a_4840_5409# a_3229_5051# 0.03325f
C84 a_8700_2159# a_8283_2049# 0.06611f
C85 sky130_fd_sc_hd__mux4_1_0.A2 a_16297_2159# 0.00107f
C86 a_7892_1793# a_6281_2043# 0
C87 a_4903_15345# a_4763_14525# 0
C88 sky130_fd_sc_hd__mux4_1_0.A2 a_9223_1793# 0.00282f
C89 a_12587_5459# sky130_fd_sc_hd__mux4_1_0.A3 0
C90 a_4839_12857# a_7749_14003# 0
C91 a_1868_1791# VDPWR 0.14821f
C92 sky130_fd_sc_hd__mux4_1_0.A2 a_5942_1761# 0
C93 uio_out[7] uio_out[6] 0.03102f
C94 a_2259_2047# a_1920_1765# 0.04737f
C95 a_16454_4503# a_9317_5049# 0
C96 a_14380_4547# a_14561_4913# 0
C97 a_3199_1791# a_2187_1765# 0.00472f
C98 a_5942_1761# a_6071_1787# 0.00758f
C99 a_16902_5839# a_16485_5729# 0.06611f
C100 VDPWR a_4905_12113# 0.4562f
C101 a_11583_15239# a_12039_15239# 0
C102 a_15711_4547# a_16539_5473# 0
C103 a_11411_5471# a_12587_5825# 0.04534f
C104 VDPWR a_12950_5825# 0.01932f
C105 a_5363_5043# a_4840_5043# 0
C106 a_16243_2049# a_15904_1767# 0.04737f
C107 a_11255_13773# a_8193_13753# 0
C108 a_6167_2153# a_6281_2043# 0
C109 a_9491_15377# a_9369_16343# 0.00144f
C110 a_8337_1793# a_8073_1793# 0
C111 a_16793_4785# a_16847_4895# 0.03622f
C112 VDPWR a_8431_5415# 0.00982f
C113 VDPWR a_14281_5833# 0
C114 a_8169_1793# a_7944_1767# 0.00487f
C115 VDPWR a_2079_5051# 0.00123f
C116 sky130_fd_sc_hd__mux4_1_0.A2 a_8073_1793# 0
C117 a_23511_14335# sky130_fd_sc_hd__mux4_1_0.A1 0.04403f
C118 a_16146_5447# a_16454_4503# 0
C119 a_4503_16339# a_4753_16339# 0.02504f
C120 a_11255_13773# a_10993_13773# 0
C121 VDPWR a_13186_4919# 0.02137f
C122 a_14771_4803# a_15188_4547# 0.03016f
C123 a_9493_12145# a_9501_13813# 0
C124 a_12323_5825# a_12142_5459# 0
C125 a_14545_5467# a_14491_5723# 0.00386f
C126 uio_in[7] uio_in[6] 0.03102f
C127 a_6429_5043# a_6165_5043# 0
C128 a_9705_12861# a_9379_14779# 0.00442f
C129 a_5363_5043# a_4423_5299# 0.13739f
C130 a_6389_13769# a_4915_10549# 0.00248f
C131 a_10499_4853# sky130_fd_sc_hd__mux4_1_0.A3 0
C132 a_5851_13769# a_5809_14763# 0
C133 ui_in[1] a_23511_14335# 0.08552f
C134 a_4915_10549# a_4837_16089# 0.01618f
C135 a_16902_5473# VDPWR 0.21501f
C136 a_12950_5459# a_11439_4597# 0
C137 a_9501_13813# a_9769_15349# 0.00159f
C138 VDPWR a_10995_12931# 0
C139 a_6335_2153# a_5269_1787# 0.04534f
C140 VDPWR a_10869_11939# 0.22337f
C141 a_4903_15345# a_4595_14775# 0
C142 a_10888_5471# a_11411_5471# 0
C143 a_12378_4553# sky130_fd_sc_hd__mux4_1_0.A3 0
C144 a_14771_4803# a_15431_5467# 0
C145 a_5363_5043# a_6429_5409# 0.04534f
C146 a_10953_14739# a_11583_15239# 0.00232f
C147 a_12769_4809# a_12533_5715# 0
C148 a_9705_12861# a_9587_13813# 0
C149 a_16902_5473# a_17425_5473# 0
C150 a_12769_4809# a_13186_4553# 0.03016f
C151 VDPWR a_10841_12931# 0.22889f
C152 VDPWR a_8263_5049# 0
C153 a_11501_15239# a_11583_15239# 0.00578f
C154 a_16243_2049# a_16129_2159# 0
C155 a_4625_15373# a_4635_13809# 0
C156 sky130_fd_sc_hd__mux4_1_0.A2 a_14233_1793# 0
C157 VDPWR a_10261_5837# 0
C158 VDPWR a_12142_5459# 0.14245f
C159 ui_in[0] a_23731_14309# 0.48785f
C160 a_12378_4553# a_10499_4853# 0
C161 a_12823_4553# a_13186_4553# 0.00985f
C162 VDPWR a_15522_4913# 0
C163 a_9621_13111# a_9501_13813# 0
C164 VDPWR a_9371_13111# 0.51474f
C165 a_11411_5471# a_12950_5459# 0.08907f
C166 VDPWR a_8169_1793# 0
C167 ui_in[0] a_24318_14385# 0.00255f
C168 sky130_fd_sc_hd__mux4_1_0.A2 a_14930_2159# 0
C169 a_6635_15235# a_7173_15235# 0.08446f
C170 a_6911_15235# VDPWR 0
C171 ui_in[5] ui_in[6] 0.03102f
C172 a_5269_1787# a_6335_1787# 0.08312f
C173 a_13473_5459# a_14491_5723# 0
C174 VDPWR a_10955_11939# 0
C175 a_4723_10577# a_4637_10577# 0.00658f
C176 a_14491_5723# a_14152_5441# 0.04737f
C177 a_14908_5467# a_15431_5467# 0
C178 a_4847_14525# a_4513_14775# 0.1679f
C179 a_4840_5409# a_2217_5025# 0
C180 a_11583_15239# a_9703_16093# 0
C181 a_4513_14775# a_4763_14525# 0.00723f
C182 a_4839_12857# a_6127_13769# 0.00253f
C183 sky130_fd_sc_hd__mux4_1_0.A1 a_18128_16189# 0
C184 a_6129_12927# a_5975_12927# 0.00401f
C185 a_15711_4547# a_17210_4895# 0.03325f
C186 a_11836_1793# a_11888_1767# 0.1439f
C187 a_9779_13785# a_9769_15349# 0.11595f
C188 a_6429_5043# a_6375_5299# 0.00386f
C189 a_18553_4938# a_17733_4529# 0.00143f
C190 VDPWR a_9381_11547# 0.50586f
C191 VDPWR a_7126_5043# 0
C192 VDPWR a_18846_5265# 0
C193 a_22274_16171# sky130_fd_sc_hd__mux4_1_0.A1 0
C194 a_10121_1793# a_10289_1793# 0
C195 VDPWR a_10025_1793# 0.00118f
C196 a_8337_2159# a_8073_2159# 0
C197 a_15119_1793# a_16660_1793# 0.08907f
C198 a_4383_2153# a_4215_2153# 0
C199 VDPWR a_16275_5839# 0
C200 VDPWR a_8700_2159# 0.02101f
C201 a_5269_1787# VDPWR 1.41387f
C202 a_16297_2159# a_16660_2159# 0.00847f
C203 a_18846_5265# a_17425_5473# 0
C204 a_5942_1761# a_2187_1765# 0.001f
C205 a_14281_5833# a_14152_5441# 0.00792f
C206 VDPWR a_12655_4553# 0
C207 VDPWR a_10289_4963# 0
C208 a_13186_4553# a_13709_4553# 0
C209 VDPWR ui_in[0] 0.81315f
C210 VDPWR a_15522_4547# 0
C211 a_10289_4963# a_10108_4597# 0
C212 VDPWR a_5890_1787# 0.13948f
C213 VDPWR a_9453_13111# 0.0252f
C214 a_4505_13107# a_4847_14525# 0
C215 a_16033_2159# a_16297_2159# 0
C216 a_15852_1793# VDPWR 0.14229f
C217 a_12194_5433# a_12533_5715# 0.04737f
C218 VDPWR ua[6] 0.00159f
C219 a_17210_4529# a_17733_4529# 0
C220 a_16454_4503# a_15711_4547# 0.11874f
C221 a_9317_5049# a_14491_5723# 0
C222 a_12587_5825# sky130_fd_sc_hd__mux4_1_0.A3 0.00113f
C223 uio_out[3] uio_out[2] 0.03102f
C224 ui_in[2] ui_in[3] 0.03102f
C225 a_2049_2157# a_2187_1765# 0
C226 a_10888_5837# a_10525_5837# 0.00847f
C227 VDPWR a_14561_4547# 0.00121f
C228 a_15242_5833# sky130_fd_sc_hd__mux4_1_0.A3 0
C229 a_14771_4803# VDPWR 0.48481f
C230 VDPWR a_11671_15239# 0.00149f
C231 a_10525_5471# a_10471_5727# 0.00386f
C232 a_6389_13769# a_6862_13645# 0.24537f
C233 a_16146_5447# a_16371_5839# 0.00559f
C234 sky130_fd_sc_hd__mux4_1_0.A2 a_12227_2049# 0.00304f
C235 a_6129_12927# a_4905_12113# 0
C236 a_6036_5017# sky130_fd_sc_hd__mux4_1_0.A3 0
C237 a_9579_12145# a_9771_12117# 0
C238 VDPWR a_12559_4553# 0.00128f
C239 a_6862_13645# a_4837_16089# 0
C240 a_2079_5417# a_1950_5025# 0.00792f
C241 a_12769_4809# a_15188_4547# 0
C242 a_4637_10577# a_4515_11543# 0.00144f
C243 a_8263_5415# a_8038_5023# 0.00559f
C244 VDPWR a_10471_5727# 0.46251f
C245 a_11255_13773# a_9769_15349# 0
C246 VDPWR a_4746_2153# 0.02101f
C247 a_4513_14775# a_4595_14775# 0.00641f
C248 a_4215_1787# a_4329_2043# 0
C249 VDPWR a_4839_12857# 1.15655f
C250 a_8794_5049# sky130_fd_sc_hd__mux4_1_0.A3 0
C251 a_12615_14007# a_9705_12861# 0
C252 a_12950_5459# a_12587_5459# 0.00985f
C253 a_9461_14779# VDPWR 0.02519f
C254 VDPWR a_12655_4919# 0
C255 sky130_fd_sc_hd__mux4_1_0.A2 a_13788_1793# 0.00121f
C256 a_16146_5447# a_14491_5723# 0.00354f
C257 a_16402_4529# a_15431_5467# 0
C258 a_10953_14739# a_11195_12931# 0
C259 VDPWR a_14908_5467# 0.21934f
C260 sky130_fd_sc_hd__mux4_1_0.A2 a_13186_4553# 0
C261 VDPWR a_9631_11297# 0.00377f
C262 a_3040_5051# a_2289_5307# 0.00682f
C263 a_2343_5417# a_2217_5025# 0.0517f
C264 uo_out[5] uo_out[4] 0.03102f
C265 a_10986_2159# a_11175_1793# 0
C266 VDPWR a_5174_5409# 0
C267 a_6089_11935# a_6281_11907# 0
C268 a_17236_5473# a_16485_5729# 0.00682f
C269 a_6629_15387# VDPWR 1.62533f
C270 a_24234_14385# a_23731_14309# 0.12294f
C271 a_24234_14385# a_24318_14385# 0.0296f
C272 sky130_fd_sc_hd__mux4_1_0.A2 a_10025_2159# 0
C273 a_10888_5471# sky130_fd_sc_hd__mux4_1_0.A3 0
C274 a_6375_5299# a_7986_5049# 0
C275 a_6281_11907# a_4915_10549# 0.43338f
C276 a_9619_16093# a_9369_16343# 0.00723f
C277 VDPWR a_14657_4547# 0
C278 a_4763_14775# a_4635_13809# 0
C279 a_11255_13773# a_12039_15239# 0.00147f
C280 a_10160_4571# sky130_fd_sc_hd__mux4_1_0.A3 0
C281 a_6389_13769# a_7749_14003# 0.00184f
C282 a_10953_14739# a_9779_13785# 0
C283 VDPWR a_9713_14529# 0.52688f
C284 clk ena 0.03102f
C285 a_13840_1767# a_13167_1793# 0.11878f
C286 a_9769_15349# a_10761_14767# 0
C287 VDPWR a_4329_2043# 0.45129f
C288 a_4721_13809# a_4913_13781# 0.00222f
C289 a_12950_5459# sky130_fd_sc_hd__mux4_1_0.A3 0
C290 a_15188_4547# a_13709_4553# 0.08907f
C291 a_10160_4571# a_10499_4853# 0.04737f
C292 a_12823_4919# a_13186_4919# 0.00847f
C293 a_9501_13813# a_4915_10549# 0.00129f
C294 a_4625_15373# a_4847_14525# 0.00215f
C295 VDPWR a_14179_2049# 0.45022f
C296 VDPWR a_10080_5471# 0.14372f
C297 a_6698_1787# a_7221_1787# 0
C298 VDPWR a_8167_5049# 0.00117f
C299 a_9779_13785# a_9703_16093# 0.01745f
C300 sky130_fd_sc_hd__mux4_1_0.A2 a_7032_2153# 0
C301 a_8377_5305# sky130_fd_sc_hd__mux4_1_0.A3 0.00302f
C302 a_4627_12141# a_4765_11543# 0
C303 a_18553_4938# VDPWR 0
C304 a_14908_5467# a_14545_5467# 0.00985f
C305 a_24234_14385# VDPWR 0.28851f
C306 ui_in[0] a_23677_14701# 0.02095f
C307 a_8337_1793# a_8283_2049# 0.00386f
C308 a_15431_5467# a_13709_4553# 0
C309 a_7113_13395# a_6635_15235# 0
C310 a_12430_4527# a_10916_4963# 0
C311 a_24241_14651# ui_in[0] 0.06316f
C312 a_13709_4553# a_14545_5833# 0
C313 VDPWR a_1898_5051# 0.14607f
C314 a_12039_15239# a_10761_14767# 0
C315 VDPWR a_10986_2159# 0
C316 a_2289_5307# a_3229_5051# 0.13963f
C317 sky130_fd_sc_hd__mux4_1_0.A2 a_8283_2049# 0.00304f
C318 a_6281_2043# a_6698_2153# 0.06611f
C319 sky130_fd_sc_hd__mux4_1_0.A2 a_17733_4529# 0
C320 a_10289_4963# a_10553_4963# 0
C321 a_5363_5043# a_5984_5043# 0.05218f
C322 a_4423_5299# a_4840_5409# 0.06611f
C323 a_4847_14525# a_5809_14763# 0.00178f
C324 a_6429_5409# a_6792_5409# 0.00847f
C325 VDPWR a_17210_4529# 0.21928f
C326 a_15242_5467# a_14491_5723# 0.00682f
C327 a_4383_1787# a_3199_1791# 0.08312f
C328 VDPWR a_16402_4529# 0.1525f
C329 a_9705_12861# a_10995_12931# 0.00312f
C330 a_10869_11939# a_9705_12861# 0
C331 a_5851_13769# a_4915_10549# 0.00192f
C332 a_11255_13773# a_10953_14739# 0
C333 a_15431_5467# a_16094_5473# 0.05191f
C334 VDPWR a_2676_1791# 0.22056f
C335 sky130_fd_sc_hd__mux4_1_0.A2 a_15188_4547# 0
C336 a_6911_15235# a_6087_14735# 0.00651f
C337 a_12769_4809# VDPWR 0.46013f
C338 a_7113_13395# a_7173_15235# 0.40674f
C339 a_9779_13785# a_4915_10549# 0.00435f
C340 VDPWR a_4477_5409# 0.0096f
C341 a_11979_13399# a_12697_14007# 0.00223f
C342 VDPWR a_12823_4553# 0.1883f
C343 a_6375_5299# sky130_fd_sc_hd__mux4_1_0.A3 0.00299f
C344 a_10841_12931# a_9705_12861# 0.29952f
C345 a_4746_1787# VDPWR 0.21796f
C346 VDPWR a_3040_5417# 0
C347 VDPWR a_6261_5043# 0
C348 a_11222_5471# sky130_fd_sc_hd__mux4_1_0.A3 0
C349 a_4119_1787# a_2187_1765# 0
C350 a_9705_12861# a_9371_13111# 0.16952f
C351 a_9896_1767# a_10025_1793# 0.00758f
C352 VDPWR a_3010_1791# 0
C353 sky130_fd_sc_hd__mux4_1_0.A3 a_10132_5445# 0.00451f
C354 sky130_fd_sc_hd__mux4_1_0.A2 a_16994_1793# 0
C355 a_9491_15377# a_9713_14529# 0.00215f
C356 a_11255_13773# a_9703_16093# 0.00515f
C357 VDPWR a_11728_13649# 0.16044f
C358 VDPWR a_16129_1793# 0
C359 a_11255_13773# a_9781_10553# 0.00248f
C360 a_4847_14525# a_4503_16339# 0
C361 a_12978_2159# a_12227_2049# 0.00696f
C362 a_3010_2157# a_3199_1791# 0
C363 a_12194_5433# a_12323_5825# 0.00792f
C364 VDPWR a_7315_5043# 1.41429f
C365 a_14771_4803# a_9317_5049# 0
C366 a_9577_15377# a_9713_14529# 0
C367 ui_in[1] a_24774_14701# 0.63058f
C368 a_6281_11907# a_6862_13645# 0.00254f
C369 a_10235_2049# a_10986_2159# 0.00696f
C370 a_4913_13781# a_5975_12927# 0.08477f
C371 a_6389_13769# a_6127_13769# 0
C372 a_16146_5447# a_16275_5839# 0.00792f
C373 a_10953_14739# a_10761_14767# 0
C374 VDPWR a_10675_14767# 0.21214f
C375 a_8337_1793# a_7944_1767# 0.02283f
C376 a_6335_2153# sky130_fd_sc_hd__mux4_1_0.A2 0
C377 sky130_fd_sc_hd__mux4_1_0.A2 a_11175_1793# 0.00285f
C378 a_9705_12861# a_9381_11547# 0
C379 a_6127_13769# a_4837_16089# 0.00702f
C380 a_9317_5049# a_10471_5727# 0
C381 ui_in[0] a_23511_14701# 0.00322f
C382 a_4839_12857# a_6129_12927# 0.00312f
C383 a_9631_11547# a_9503_10581# 0
C384 uio_in[4] uio_in[3] 0.03102f
C385 sky130_fd_sc_hd__mux4_1_0.A2 a_7944_1767# 0.00211f
C386 sky130_fd_sc_hd__mux4_1_0.A2 a_23731_14309# 0
C387 a_10261_5471# sky130_fd_sc_hd__mux4_1_0.A3 0
C388 VDPWR a_13709_4553# 1.42843f
C389 a_5269_1787# a_5080_2153# 0
C390 a_16583_4895# sky130_fd_sc_hd__mux4_1_0.A3 0
C391 a_9379_14779# a_9369_16343# 0.00102f
C392 sky130_fd_sc_hd__mux4_1_0.A2 a_24318_14385# 0.05111f
C393 VDPWR a_11147_11911# 0.30098f
C394 a_10761_14767# a_9703_16093# 0
C395 a_16902_5473# a_16539_5473# 0.00985f
C396 VDPWR a_11250_4963# 0
C397 a_9621_12861# a_4915_10549# 0
C398 VDPWR a_12194_5433# 0.35585f
C399 a_8794_5049# a_10160_4571# 0
C400 a_4765_11293# a_4515_11543# 0.00723f
C401 a_14179_2049# a_14065_1793# 0
C402 a_23511_14335# a_23677_14335# 0.00648f
C403 a_9705_12861# a_9453_13111# 0
C404 a_6165_5043# a_6036_5017# 0.00758f
C405 a_24234_14385# a_24241_14651# 0.13413f
C406 a_16902_5473# a_15711_4547# 0
C407 sky130_fd_sc_hd__mux4_1_0.A2 a_6335_1787# 0
C408 uio_in[0] ui_in[7] 0.03102f
C409 a_10841_12931# a_10923_12931# 0.00517f
C410 a_14908_5833# a_14491_5723# 0.06611f
C411 a_4763_14775# a_4847_14525# 0.07979f
C412 VDPWR a_14432_4521# 0.35559f
C413 sky130_fd_sc_hd__mux4_1_0.A2 a_12113_1793# 0
C414 a_4839_12857# a_6087_14735# 0.02474f
C415 a_6335_1787# a_6071_1787# 0
C416 a_16033_1793# VDPWR 0.00118f
C417 a_6281_11907# a_7749_14003# 0.19234f
C418 a_4585_16339# a_4837_16089# 0
C419 a_12281_2159# a_12227_2049# 0.03622f
C420 a_4637_10577# a_4915_10549# 0.1296f
C421 VDPWR a_16094_5473# 0.14176f
C422 a_10385_4597# a_10499_4853# 0
C423 a_4913_13781# a_4905_12113# 0.00627f
C424 a_2289_5307# a_2217_5025# 0.25757f
C425 a_13520_4919# sky130_fd_sc_hd__mux4_1_0.A3 0
C426 a_7999_14003# a_6281_11907# 0
C427 a_14561_4913# sky130_fd_sc_hd__mux4_1_0.A3 0
C428 a_2145_2157# a_1920_1765# 0.00559f
C429 a_14596_1793# a_14179_2049# 0.03016f
C430 a_12823_4919# a_12655_4919# 0
C431 a_9629_14779# a_9769_15349# 0.00327f
C432 VDPWR a_4753_16089# 0.00472f
C433 a_16679_4895# sky130_fd_sc_hd__mux4_1_0.A3 0
C434 a_16371_5473# sky130_fd_sc_hd__mux4_1_0.A3 0
C435 a_8337_1793# VDPWR 0.18611f
C436 a_7892_1793# a_7221_1787# 0.05168f
C437 a_8794_5049# a_8377_5305# 0.03016f
C438 a_6629_15387# a_6087_14735# 0.09734f
C439 a_16146_5447# a_14908_5467# 0
C440 a_15852_1793# a_15904_1767# 0.1439f
C441 a_15711_4547# a_15522_4913# 0
C442 a_5942_1761# a_6071_2153# 0.00792f
C443 a_8431_5415# a_8038_5023# 0.02301f
C444 a_14065_2159# a_14179_2049# 0
C445 a_5851_13769# a_6862_13645# 0
C446 sky130_fd_sc_hd__mux4_1_0.A2 VDPWR 0.50362f
C447 a_6089_11935# a_6003_11935# 0.00658f
C448 a_9501_13813# a_7749_14003# 0
C449 sky130_fd_sc_hd__mux4_1_0.A2 a_10108_4597# 0
C450 VDPWR a_6389_13769# 0.47275f
C451 a_9461_14779# a_9705_12861# 0
C452 a_16793_4785# a_17733_4529# 0.14301f
C453 a_14545_5467# a_13709_4553# 0
C454 a_14825_4913# sky130_fd_sc_hd__mux4_1_0.A3 0
C455 VDPWR a_6071_1787# 0.00122f
C456 a_18839_4938# a_18625_4938# 0.00557f
C457 a_18553_4938# a_9317_5049# 0.00526f
C458 VDPWR a_4837_16089# 1.41996f
C459 a_24774_14701# ua[0] 0.00399f
C460 a_6003_11935# a_4915_10549# 0
C461 a_10888_5471# a_8377_5305# 0
C462 a_10887_13773# a_10717_13773# 0.00167f
C463 a_10525_5837# sky130_fd_sc_hd__mux4_1_0.A3 0.0014f
C464 a_4505_13107# a_4765_11543# 0
C465 VDPWR a_7126_5409# 0
C466 a_20384_16179# a_19510_16177# 0.10112f
C467 a_6911_15235# a_6635_15235# 0.00119f
C468 a_10160_4571# a_8377_5305# 0
C469 a_8263_5415# a_8431_5415# 0
C470 uio_oe[4] uio_oe[5] 0.03102f
C471 a_6375_5299# a_6036_5017# 0.04737f
C472 a_20384_16179# VDPWR 0.47674f
C473 a_12419_5459# a_12533_5715# 0
C474 a_4903_15345# a_4513_14775# 0.00566f
C475 a_9705_12861# a_9713_14529# 0.18435f
C476 a_6329_12927# a_6862_13645# 0.10646f
C477 a_10499_4853# a_10525_5837# 0
C478 a_2289_5307# a_2175_5051# 0
C479 a_5080_2153# a_4329_2043# 0.00696f
C480 a_15431_5467# a_16485_5729# 0.21187f
C481 a_15119_1793# a_16297_1793# 0.08312f
C482 a_5851_13769# a_7749_14003# 0
C483 sky130_fd_sc_hd__mux4_1_0.A1 sky130_fd_sc_hd__mux4_1_0.A3 0.00503f
C484 a_8038_5023# a_8263_5049# 0.00487f
C485 a_14377_5467# a_14491_5723# 0
C486 a_12769_4809# a_9317_5049# 0
C487 a_16793_4785# a_15431_5467# 0
C488 a_6911_15235# a_7173_15235# 0
C489 a_5363_5043# VDPWR 1.41627f
C490 a_6429_5409# a_6165_5409# 0
C491 a_13709_4553# a_14152_5441# 0
C492 a_16539_5839# sky130_fd_sc_hd__mux4_1_0.A3 0.00117f
C493 a_4505_13107# a_4627_12141# 0.00144f
C494 a_10235_2049# sky130_fd_sc_hd__mux4_1_0.A2 0.00304f
C495 a_3938_1787# a_2187_1765# 0.00121f
C496 a_14771_4803# a_15711_4547# 0.13762f
C497 a_11411_5471# a_11222_5837# 0
C498 a_2343_5417# a_4084_5017# 0
C499 ui_in[1] sky130_fd_sc_hd__mux4_1_0.A3 0.07335f
C500 a_14930_1793# a_14179_2049# 0.00682f
C501 a_7113_13395# a_5975_12927# 0
C502 uo_out[6] uo_out[5] 0.03102f
C503 a_15188_4913# sky130_fd_sc_hd__mux4_1_0.A3 0
C504 ui_in[0] a_24407_14651# 0.00109f
C505 a_11979_13399# a_10717_13773# 0
C506 a_2217_5025# sky130_fd_sc_hd__mux4_1_0.A3 0.11807f
C507 a_9493_12145# a_9579_12145# 0.00658f
C508 a_18839_4938# sky130_fd_sc_hd__mux4_1_0.A3 0.0023f
C509 a_14432_4521# a_14152_5441# 0
C510 a_12865_14007# a_11979_13399# 0.00205f
C511 a_12769_4809# a_12823_4919# 0.03622f
C512 a_3990_1761# a_4329_2043# 0.04737f
C513 a_4627_12141# a_4713_12141# 0.00658f
C514 a_7315_5043# a_9317_5049# 0
C515 a_4755_12857# a_4505_13107# 0.00723f
C516 a_15904_1767# a_14179_2049# 0.00358f
C517 a_3938_1787# a_4119_2153# 0
C518 a_10160_4571# a_10132_5445# 0
C519 a_4839_12857# a_4755_13107# 0.08134f
C520 a_4215_1787# a_2187_1765# 0
C521 VDPWR a_11583_15239# 0
C522 a_9317_5049# a_13709_4553# 0.0303f
C523 a_12793_14007# a_12615_14007# 0.00412f
C524 a_16902_5839# sky130_fd_sc_hd__mux4_1_0.A3 0.00192f
C525 a_2175_5417# a_2343_5417# 0
C526 a_1898_5051# a_2079_5417# 0
C527 sky130_fd_sc_hd__mux4_1_0.A2 a_24241_14651# 0.03575f
C528 VDPWR a_16486_16197# 0.49757f
C529 a_9379_14779# a_9371_13111# 0
C530 a_14657_4913# sky130_fd_sc_hd__mux4_1_0.A3 0
C531 ui_in[0] a_24962_14701# 0.02482f
C532 a_8377_5305# a_10132_5445# 0
C533 a_21506_16181# sky130_fd_sc_hd__mux4_1_0.A1 0
C534 a_12194_5433# a_9317_5049# 0
C535 sky130_fd_sc_hd__mux4_1_0.A2 a_14065_1793# 0
C536 a_24152_14385# a_24774_14701# 0
C537 a_8431_5415# a_8794_5415# 0.00847f
C538 a_6792_5043# VDPWR 0.21801f
C539 a_6629_15387# a_6635_15235# 0.16833f
C540 a_16847_4895# sky130_fd_sc_hd__mux4_1_0.A3 0
C541 a_9223_1793# a_10289_1793# 0.08312f
C542 a_14432_4521# a_9317_5049# 0
C543 VDPWR a_16485_5729# 0.43938f
C544 a_9705_12861# a_11728_13649# 0.00327f
C545 sky130_fd_sc_hd__mux4_1_0.A2 a_12017_1793# 0
C546 VDPWR a_2187_1765# 1.68953f
C547 ui_in[4] ui_in[3] 0.03102f
C548 a_10385_4597# a_10160_4571# 0.00487f
C549 a_12430_4527# a_12533_5715# 0
C550 a_4839_12857# a_7173_15235# 0.00685f
C551 VDPWR a_16660_2159# 0.0192f
C552 VDPWR a_16793_4785# 0.46738f
C553 a_2259_2047# a_2145_2157# 0
C554 a_1950_5025# a_2079_5051# 0.00758f
C555 a_12281_2159# a_11175_1793# 0.04534f
C556 sky130_fd_sc_hd__mux4_1_0.A2 a_14596_1793# 0
C557 a_5975_12927# a_4905_12113# 0
C558 a_5895_14763# a_4903_15345# 0
C559 a_16485_5729# a_17425_5473# 0.13858f
C560 VDPWR a_12978_2159# 0
C561 a_9705_12861# a_10675_14767# 0.21957f
C562 sky130_fd_sc_hd__mux4_1_0.A3 a_10916_4963# 0
C563 a_9631_11547# a_9371_13111# 0
C564 sky130_fd_sc_hd__mux4_1_0.A2 a_10652_1793# 0
C565 a_16793_4785# a_17425_5473# 0
C566 a_16033_2159# VDPWR 0
C567 a_5942_1761# a_6167_2153# 0.00559f
C568 a_4839_12857# a_4913_13781# 0.44871f
C569 a_6629_15387# a_7173_15235# 0.002f
C570 sky130_fd_sc_hd__mux4_1_0.A2 a_14065_2159# 0
C571 VDPWR a_6281_11907# 0.30528f
C572 VDPWR a_4119_2153# 0
C573 a_5851_13769# a_6127_13769# 0.00119f
C574 a_2049_2157# a_1920_1765# 0.00792f
C575 sky130_fd_sc_hd__mux4_1_0.A2 a_17544_4529# 0
C576 a_6281_2043# a_7221_1787# 0.13739f
C577 a_15904_1767# a_16129_1793# 0.00487f
C578 a_14432_4521# a_12823_4919# 0
C579 a_8337_2159# a_6281_2043# 0
C580 sky130_fd_sc_hd__mux4_1_0.A2 a_9034_2159# 0
C581 a_2259_2047# a_3199_1791# 0.13962f
C582 a_10499_4853# a_10916_4963# 0.06611f
C583 VDPWR a_4753_16339# 0.33641f
C584 sky130_fd_sc_hd__mux4_1_0.A2 a_10916_4597# 0
C585 a_11147_11911# a_9705_12861# 0.02321f
C586 a_8431_5049# sky130_fd_sc_hd__mux4_1_0.A3 0
C587 sky130_fd_sc_hd__mux4_1_0.A2 a_10553_4597# 0
C588 a_4625_15373# a_4903_15345# 0.12165f
C589 a_4765_11543# a_4515_11543# 0.02504f
C590 a_9631_11547# a_9381_11547# 0.02504f
C591 a_16146_5447# a_16094_5473# 0.1439f
C592 a_23511_14335# a_23731_14309# 0.0457f
C593 a_16583_4529# VDPWR 0.00132f
C594 sky130_fd_sc_hd__mux4_1_0.A2 a_7032_1787# 0
C595 a_4119_1787# a_4383_1787# 0
C596 a_24234_14385# a_24407_14651# 0.00222f
C597 a_17210_4529# a_15711_4547# 0.08907f
C598 sky130_fd_sc_hd__mux4_1_0.A2 a_9896_1767# 0.00211f
C599 a_16402_4529# a_15711_4547# 0.05149f
C600 VDPWR a_9501_13813# 0.43873f
C601 a_16454_4503# a_14771_4803# 0.00271f
C602 a_9503_10581# a_9381_11547# 0.00144f
C603 a_4505_13107# a_4513_14775# 0
C604 a_6087_14735# a_6389_13769# 0
C605 a_11810_13649# a_11728_13649# 0.00477f
C606 a_6087_14735# a_4837_16089# 0.29394f
C607 a_11222_5837# sky130_fd_sc_hd__mux4_1_0.A3 0
C608 a_10993_13773# a_10717_13773# 0.00119f
C609 a_6036_5017# a_2217_5025# 0
C610 a_12281_2159# VDPWR 0.0097f
C611 a_4903_15345# a_5809_14763# 0.00346f
C612 a_7944_1767# a_8073_2159# 0.00792f
C613 a_8038_5023# a_8167_5049# 0.00758f
C614 VDPWR a_11195_12931# 0.31314f
C615 a_14233_1793# a_13969_1793# 0
C616 a_9461_14779# a_9379_14779# 0.00641f
C617 a_4627_12141# a_4515_11543# 0
C618 a_14419_5441# a_12533_5715# 0
C619 a_7831_14003# a_4915_10549# 0
C620 a_10261_5471# a_10132_5445# 0.00758f
C621 a_16033_1793# a_15904_1767# 0.00758f
C622 a_4839_12857# a_4721_13809# 0
C623 a_2289_5307# a_2343_5051# 0.00386f
C624 a_18371_4938# a_17733_4529# 0.15188f
C625 a_24234_14385# a_24962_14701# 0.1456f
C626 a_14930_1793# sky130_fd_sc_hd__mux4_1_0.A2 0
C627 VDPWR a_5851_13769# 0.44589f
C628 VDPWR a_23511_14335# 0.05794f
C629 a_13840_1767# a_14179_2049# 0.04737f
C630 a_17236_5839# a_17425_5473# 0
C631 a_14100_5467# a_12533_5715# 0
C632 a_11810_13649# a_11147_11911# 0
C633 VDPWR a_9779_13785# 0.76122f
C634 a_13284_5459# a_12533_5715# 0.00682f
C635 a_17254_16187# a_16486_16197# 0.1036f
C636 a_9713_14529# a_9379_14779# 0.1679f
C637 VDPWR a_12419_5459# 0
C638 sky130_fd_sc_hd__mux4_1_0.A2 a_11888_1767# 0.00211f
C639 sky130_fd_sc_hd__mux4_1_0.A2 a_15904_1767# 0.00324f
C640 a_12281_1793# a_12227_2049# 0.00386f
C641 a_4903_15345# a_4503_16339# 0
C642 a_2289_5307# a_4084_5017# 0.00286f
C643 a_5984_5043# a_6165_5409# 0
C644 sky130_fd_sc_hd__mux4_1_0.A1 a_11979_13399# 0.03491f
C645 a_15711_4547# a_13709_4553# 0
C646 a_6429_5409# sky130_fd_sc_hd__mux4_1_0.A3 0
C647 VDPWR a_6792_5409# 0.02103f
C648 a_9493_12145# a_9771_12117# 0.12057f
C649 a_13167_1793# a_14179_2049# 0.21187f
C650 a_8700_1793# a_7221_1787# 0.08907f
C651 VDPWR a_14380_4547# 0.141f
C652 VDPWR a_8073_2159# 0
C653 VDPWR a_14233_2159# 0.00967f
C654 a_24152_14385# sky130_fd_sc_hd__mux4_1_0.A3 0.01336f
C655 a_18742_16187# sky130_fd_sc_hd__mux4_1_0.A1 0
C656 a_9579_12145# a_4915_10549# 0
C657 a_11439_4597# a_12533_5715# 0
C658 a_10887_13773# a_9769_15349# 0.00818f
C659 uio_oe[3] uio_oe[2] 0.03102f
C660 sky130_fd_sc_hd__mux4_1_0.A2 a_11250_4597# 0
C661 a_13186_4553# a_11439_4597# 0.08907f
C662 VDPWR a_6329_12927# 0.31314f
C663 a_16847_4529# VDPWR 0.18788f
C664 VDPWR a_4840_5409# 0.02103f
C665 a_16243_2049# a_16129_1793# 0
C666 a_14281_5467# a_14419_5441# 0
C667 uio_in[1] uio_in[0] 0.03102f
C668 a_12865_14007# sky130_fd_sc_hd__mux4_1_0.A1 0
C669 a_9491_15377# a_9501_13813# 0
C670 VDPWR a_6021_13769# 0
C671 VDPWR a_10289_4597# 0.00151f
C672 a_10525_5837# a_10132_5445# 0.02301f
C673 a_4625_15373# a_4513_14775# 0
C674 a_7315_5043# a_8038_5023# 0.11881f
C675 a_10471_5727# a_10357_5837# 0
C676 uio_oe[5] uio_oe[6] 0.03102f
C677 a_11411_5471# a_12533_5715# 0.21188f
C678 VDPWR a_4635_13809# 0.43865f
C679 a_12769_4809# a_13520_4553# 0.00682f
C680 a_19510_16177# a_18128_16189# 0
C681 a_9317_5049# a_16485_5729# 0
C682 a_2175_5417# a_2289_5307# 0
C683 a_17544_4529# a_16793_4785# 0.00682f
C684 a_7113_13395# a_4839_12857# 0.00446f
C685 clk rst_n 0.03102f
C686 a_16793_4785# a_9317_5049# 0
C687 a_4763_14775# a_4903_15345# 0.00327f
C688 a_9781_10553# a_12697_14007# 0
C689 VDPWR a_18128_16189# 0.3744f
C690 a_5942_1761# a_6281_2043# 0.04737f
C691 a_11255_13773# VDPWR 0.47275f
C692 a_9621_12861# VDPWR 0.00415f
C693 a_8283_2049# a_9034_1793# 0.00682f
C694 sky130_fd_sc_hd__mux4_1_0.A2 a_15711_4547# 0.00101f
C695 a_6717_15235# VDPWR 0
C696 a_17236_5473# sky130_fd_sc_hd__mux4_1_0.A3 0
C697 a_16454_4503# a_16402_4529# 0.1439f
C698 sky130_fd_sc_hd__mux4_1_0.A2 a_16129_2159# 0
C699 VDPWR a_22274_16171# 0.57061f
C700 VDPWR a_8167_5415# 0
C701 a_17544_4895# a_17733_4529# 0
C702 a_8794_5049# a_8431_5049# 0.00985f
C703 a_3040_5051# a_2217_5025# 0
C704 a_4513_14775# a_5809_14763# 0
C705 a_4839_12857# a_5975_12927# 0.29952f
C706 a_10289_2159# a_10121_2159# 0
C707 a_2313_1791# a_2145_1791# 0
C708 VDPWR a_4637_10577# 0.43168f
C709 a_11979_13399# a_9769_15349# 0
C710 a_6335_2153# a_6071_2153# 0
C711 a_14908_5833# a_13709_4553# 0
C712 a_6698_1787# a_7944_1767# 0
C713 a_14419_5441# a_14545_5833# 0.04534f
C714 a_16146_5447# a_16485_5729# 0.04737f
C715 a_10869_11939# a_10841_12931# 0
C716 a_10841_12931# a_10995_12931# 0.00401f
C717 a_14419_5441# a_15431_5467# 0
C718 a_6635_15235# a_4837_16089# 0.23067f
C719 a_9713_14529# a_9369_16343# 0
C720 a_14771_4803# a_14491_5723# 0
C721 a_4597_11543# a_4515_11543# 0.00641f
C722 a_10717_13773# a_9769_15349# 0.16757f
C723 VDPWR a_5933_13769# 0
C724 VDPWR a_10761_14767# 0
C725 sky130_fd_sc_hd__mux4_1_0.A3 a_16275_5473# 0
C726 a_12430_4527# VDPWR 0.36801f
C727 a_14825_4913# a_14561_4913# 0
C728 a_10160_4571# a_8431_5049# 0
C729 a_10955_11939# a_10869_11939# 0.00658f
C730 a_6698_1787# a_6335_1787# 0.00985f
C731 a_5080_2153# a_2187_1765# 0
C732 a_10675_14767# a_9379_14779# 0
C733 VDPWR a_6003_11935# 0.22336f
C734 VDPWR a_18371_4938# 0.15241f
C735 sky130_fd_sc_hd__mux4_1_0.A2 a_16243_2049# 0.15654f
C736 a_10841_12931# a_9371_13111# 0
C737 sky130_fd_sc_hd__mux4_1_0.A1 a_8193_13753# 0.14763f
C738 a_6389_13769# a_7173_15235# 0.00147f
C739 a_18625_5265# sky130_fd_sc_hd__mux4_1_0.A3 0
C740 a_2313_2157# a_2187_1765# 0.05199f
C741 VDPWR a_16660_1793# 0.21452f
C742 a_12039_15239# a_11979_13399# 0.40674f
C743 a_12644_1793# a_12227_2049# 0.03016f
C744 a_7173_15235# a_4837_16089# 0.04818f
C745 VDPWR a_2343_5417# 0.00939f
C746 a_4513_14775# a_4503_16339# 0.00102f
C747 a_1898_5051# a_1950_5025# 0.1439f
C748 a_4215_1787# a_4383_1787# 0
C749 a_4423_5299# a_6036_5017# 0.00419f
C750 a_23677_14335# sky130_fd_sc_hd__mux4_1_0.A3 0
C751 a_14908_5467# a_14491_5723# 0.03016f
C752 a_4477_5043# a_2289_5307# 0
C753 a_18371_4938# a_17425_5473# 0.08028f
C754 sky130_fd_sc_hd__mux4_1_0.A2 a_24962_14701# 0.00234f
C755 a_4839_12857# a_4905_12113# 0.04364f
C756 a_4913_13781# a_6389_13769# 0
C757 a_12039_15239# a_10717_13773# 0
C758 a_4383_2153# a_3199_1791# 0.04534f
C759 VDPWR a_10888_5837# 0.02103f
C760 a_8431_5049# a_8377_5305# 0.00386f
C761 a_7831_14003# a_7749_14003# 0.00695f
C762 a_12865_14007# a_12039_15239# 0
C763 a_12323_5459# a_12194_5433# 0.00758f
C764 a_4913_13781# a_4837_16089# 0.01745f
C765 a_6698_1787# VDPWR 0.21798f
C766 a_12587_5459# a_12533_5715# 0.00386f
C767 a_9128_5049# sky130_fd_sc_hd__mux4_1_0.A3 0
C768 a_6429_5409# a_6036_5017# 0.02301f
C769 a_4505_13107# a_4515_11543# 0.00102f
C770 a_3229_5051# a_2217_5025# 0.00478f
C771 sky130_fd_sc_hd__mux4_1_0.A2 a_13840_1767# 0.00211f
C772 a_3990_1761# a_2187_1765# 0.00211f
C773 a_8700_1793# a_9223_1793# 0
C774 a_9371_13111# a_9381_11547# 0.00102f
C775 VDPWR a_6071_2153# 0
C776 uio_oe[1] uio_oe[2] 0.03102f
C777 sky130_fd_sc_hd__mux4_1_0.A2 a_13520_4553# 0
C778 a_10887_13773# a_9703_16093# 0.00246f
C779 a_16033_2159# a_15904_1767# 0.00792f
C780 a_7927_14003# a_4915_10549# 0
C781 a_9705_12861# a_9501_13813# 0.00246f
C782 a_9771_12117# a_9703_16093# 0
C783 VDPWR a_4383_1787# 0.18611f
C784 a_2313_1791# VDPWR 0.18286f
C785 a_7315_5043# a_8794_5415# 0.03325f
C786 a_12281_1793# a_11175_1793# 0.08312f
C787 VDPWR a_6805_15235# 0.00149f
C788 a_9781_10553# a_9771_12117# 0.0298f
C789 a_4763_14775# a_4513_14775# 0.02504f
C790 a_10121_1793# a_9223_1793# 0
C791 sky130_fd_sc_hd__mux4_1_0.A2 a_13167_1793# 0.00282f
C792 a_2343_5417# a_2706_5417# 0.00847f
C793 a_9453_13111# a_9371_13111# 0.00641f
C794 a_6281_2043# a_6167_1787# 0
C795 a_4119_2153# a_3990_1761# 0.00792f
C796 a_12644_2159# a_12227_2049# 0.06611f
C797 VDPWR a_14419_5441# 1.26078f
C798 a_14065_2159# a_14233_2159# 0
C799 a_5851_13769# a_6087_14735# 0
C800 a_16485_5729# a_16539_5473# 0.00386f
C801 a_11195_12931# a_9705_12861# 0.08252f
C802 a_17254_16187# a_18128_16189# 0.10464f
C803 a_9769_15349# a_8193_13753# 0.00127f
C804 sky130_fd_sc_hd__mux4_1_0.A2 a_16454_4503# 0
C805 a_12533_5715# sky130_fd_sc_hd__mux4_1_0.A3 0.00752f
C806 a_11501_15239# a_11979_13399# 0
C807 a_5895_14763# a_5809_14763# 0.00658f
C808 a_4847_14525# a_4711_15373# 0
C809 VDPWR a_2676_2157# 0.02202f
C810 a_23511_14335# a_23511_14701# 0.00987f
C811 a_14825_4913# a_15188_4913# 0.00847f
C812 a_15711_4547# a_16485_5729# 0
C813 VDPWR a_6165_5409# 0
C814 a_14771_4803# a_15522_4913# 0.00696f
C815 a_18625_4938# a_17733_4529# 0.19558f
C816 VDPWR a_9034_1793# 0
C817 a_24774_14701# a_23731_14309# 0.00253f
C818 a_10357_5471# sky130_fd_sc_hd__mux4_1_0.A3 0
C819 a_13969_2159# a_13788_1793# 0
C820 a_16847_4895# a_16583_4895# 0
C821 a_16793_4785# a_15711_4547# 0.21188f
C822 VDPWR a_17544_4895# 0
C823 VDPWR a_4847_14525# 0.52692f
C824 a_24318_14385# a_24774_14701# 0.01242f
C825 a_10953_14739# a_10717_13773# 0
C826 VDPWR a_13284_5459# 0
C827 a_3010_2157# VDPWR 0
C828 a_10471_5727# a_12142_5459# 0
C829 a_9771_12117# a_4915_10549# 0.00452f
C830 a_12281_2159# a_11888_1767# 0.02301f
C831 VDPWR a_14100_5467# 0.13366f
C832 a_12281_1793# a_12113_1793# 0
C833 VDPWR a_4763_14525# 0.00474f
C834 sky130_fd_sc_hd__mux4_1_0.A2 a_8169_2159# 0
C835 a_10993_13773# a_9769_15349# 0
C836 a_2145_1791# a_1920_1765# 0.00487f
C837 a_9779_13785# a_9705_12861# 0.44871f
C838 a_10553_4597# a_10289_4597# 0
C839 sky130_fd_sc_hd__mux4_1_0.A2 a_11836_1793# 0.00121f
C840 VDPWR a_6429_5043# 0.18614f
C841 a_11979_13399# a_9703_16093# 0
C842 a_2217_5025# a_4309_5409# 0
C843 VDPWR a_4215_2153# 0
C844 a_5269_1787# a_5890_1787# 0.05218f
C845 a_9781_10553# a_11979_13399# 0.20109f
C846 a_6329_12927# a_6087_14735# 0
C847 a_12039_15239# a_8193_13753# 0.002f
C848 VDPWR a_12559_4919# 0
C849 ui_in[1] sky130_fd_sc_hd__mux4_1_0.A1 0.00113f
C850 a_10717_13773# a_9703_16093# 0.08387f
C851 a_7892_1793# a_7944_1767# 0.1439f
C852 VDPWR a_11439_4597# 1.63906f
C853 VDPWR a_12281_1793# 0.18611f
C854 a_16679_4895# a_16847_4895# 0
C855 a_14419_5441# a_14545_5467# 0.08312f
C856 a_9781_10553# a_10717_13773# 0.00192f
C857 a_6944_13645# a_6862_13645# 0.00477f
C858 a_14657_4913# a_14825_4913# 0
C859 sky130_fd_sc_hd__mux4_1_0.A2 a_10652_2159# 0
C860 a_16583_4529# a_15711_4547# 0
C861 uio_in[2] uio_in[3] 0.03102f
C862 a_12194_5433# a_12419_5825# 0.00559f
C863 a_6335_2153# a_6167_2153# 0
C864 a_12865_14007# a_9781_10553# 0
C865 a_6792_5043# a_8038_5023# 0
C866 a_14281_5467# sky130_fd_sc_hd__mux4_1_0.A3 0
C867 a_14771_4803# a_15522_4547# 0.00682f
C868 a_11147_11911# a_12793_14007# 0.00264f
C869 VDPWR a_24774_14701# 0.226f
C870 a_16243_2049# a_16660_2159# 0.06611f
C871 a_9713_14529# a_9371_13111# 0
C872 a_9631_11297# a_9381_11547# 0.00723f
C873 VDPWR a_11411_5471# 1.44192f
C874 a_6717_15235# a_6087_14735# 0.00232f
C875 a_4625_15373# a_4503_16339# 0.00144f
C876 a_17733_4529# sky130_fd_sc_hd__mux4_1_0.A3 0.01989f
C877 a_12430_4527# a_9317_5049# 0
C878 a_11147_11911# a_12615_14007# 0.19234f
C879 VDPWR a_4765_11293# 0.00377f
C880 VDPWR a_9629_14779# 0.33336f
C881 VDPWR a_12017_2159# 0
C882 a_6281_11907# a_7173_15235# 0.09952f
C883 a_10080_5471# a_10261_5837# 0
C884 a_4840_5043# a_3229_5051# 0.08907f
C885 a_6429_5409# a_6375_5299# 0.03622f
C886 a_12769_4809# a_13186_4919# 0.06611f
C887 a_7113_13395# a_6389_13769# 0.0615f
C888 a_9317_5049# a_18371_4938# 0.24923f
C889 a_9779_13785# a_10799_13773# 0
C890 VDPWR a_13969_1793# 0.00118f
C891 a_15188_4547# a_14825_4547# 0.00985f
C892 a_11255_13773# a_9705_12861# 0.04676f
C893 a_9621_12861# a_9705_12861# 0.00208f
C894 VDPWR a_4595_14775# 0.02519f
C895 a_7113_13395# a_4837_16089# 0
C896 a_16485_5729# a_17210_4895# 0
C897 a_14491_5723# a_13709_4553# 0.00129f
C898 VDPWR a_7892_1793# 0.13939f
C899 a_12644_1793# a_11175_1793# 0.08907f
C900 a_2289_5307# a_4032_5043# 0
C901 a_16243_2049# a_16994_2159# 0.00696f
C902 a_16902_5839# a_16539_5839# 0.00847f
C903 a_14419_5441# a_14152_5441# 0.11855f
C904 a_14419_5441# a_13473_5459# 0.00633f
C905 a_10953_14739# a_8193_13753# 0.09734f
C906 a_16793_4785# a_17210_4895# 0.06611f
C907 a_11501_15239# a_8193_13753# 0.16833f
C908 a_7315_5043# a_8431_5415# 0.04534f
C909 VDPWR a_10289_1793# 0.18613f
C910 a_12587_5825# a_12533_5715# 0.03622f
C911 a_5269_1787# a_4329_2043# 0.13739f
C912 a_12430_4527# a_12823_4919# 0.02301f
C913 a_14377_5833# sky130_fd_sc_hd__mux4_1_0.A3 0
C914 VDPWR a_1920_1765# 0.36069f
C915 a_4903_15345# a_6862_13645# 0
C916 a_9501_13813# a_7173_15235# 0
C917 VDPWR a_2289_5307# 0.4493f
C918 a_5975_12927# a_4837_16089# 0
C919 sky130_fd_sc_hd__mux4_1_0.A3 a_14545_5833# 0.00115f
C920 a_15431_5467# sky130_fd_sc_hd__mux4_1_0.A3 0.00685f
C921 a_7032_2153# a_6281_2043# 0.00696f
C922 VDPWR a_7986_5049# 0.13941f
C923 uo_out[7] uio_out[0] 0.03102f
C924 a_14432_4521# a_14491_5723# 0
C925 a_5890_1787# a_4329_2043# 0
C926 VDPWR a_6167_2153# 0
C927 a_16094_5473# a_14491_5723# 0
C928 a_4763_14775# a_4625_15373# 0
C929 a_14100_5467# a_14152_5441# 0.1439f
C930 a_14100_5467# a_13473_5459# 0.00621f
C931 a_4423_5299# a_3229_5051# 0.21187f
C932 a_12039_15239# sky130_fd_sc_hd__mux4_1_0.A1 0.04277f
C933 a_8337_2159# a_7221_1787# 0.04534f
C934 a_8193_13753# a_9703_16093# 0.35109f
C935 a_16454_4503# a_16485_5729# 0
C936 a_14771_4803# a_14657_4547# 0
C937 a_9705_12861# a_10761_14767# 0
C938 VDPWR a_7831_14003# 0
C939 a_11671_15239# a_9713_14529# 0.00624f
C940 a_7927_14003# a_7749_14003# 0.00412f
C941 a_16454_4503# a_16793_4785# 0.04737f
C942 VDPWR a_18625_4938# 0.11951f
C943 a_12978_2159# a_13167_1793# 0
C944 a_10289_2159# a_9223_1793# 0.04534f
C945 a_2049_1791# VDPWR 0.00125f
C946 a_15852_1793# a_14179_2049# 0
C947 a_12978_1793# a_12227_2049# 0.00682f
C948 a_16847_4529# a_15711_4547# 0.08312f
C949 a_24234_14385# ui_in[0] 0.28585f
C950 ui_in[1] ua[0] 0.48995f
C951 a_18625_4938# a_17425_5473# 0.06919f
C952 a_14419_5441# a_9317_5049# 0.00543f
C953 a_10841_12931# a_11728_13649# 0
C954 sky130_fd_sc_hd__mux4_1_0.A3 a_23731_14309# 0.1036f
C955 a_5984_5043# a_6036_5017# 0.1439f
C956 a_10993_13773# a_9703_16093# 0.00702f
C957 a_7315_5043# a_8263_5049# 0
C958 a_11255_13773# a_10799_13773# 0
C959 a_5851_13769# a_7173_15235# 0
C960 a_11255_13773# a_11810_13649# 0.00183f
C961 a_4505_13107# a_4587_13107# 0.00641f
C962 a_12644_2159# a_11175_1793# 0.03325f
C963 a_24318_14385# sky130_fd_sc_hd__mux4_1_0.A3 0.04268f
C964 a_4746_2153# a_4329_2043# 0.06611f
C965 a_9128_5049# a_8377_5305# 0.00682f
C966 a_9461_14779# a_9713_14529# 0
C967 VDPWR a_12644_1793# 0.21796f
C968 VDPWR a_12587_5459# 0.18755f
C969 a_12323_5825# sky130_fd_sc_hd__mux4_1_0.A3 0
C970 a_10385_4963# sky130_fd_sc_hd__mux4_1_0.A3 0
C971 a_16297_2159# a_15119_1793# 0.04534f
C972 a_4635_13809# a_4755_13107# 0
C973 a_9621_13111# a_9493_12145# 0
C974 a_9491_15377# a_9629_14779# 0
C975 a_10235_2049# a_10289_1793# 0.00386f
C976 a_10841_12931# a_10675_14767# 0
C977 a_6087_14735# a_6805_15235# 0.00366f
C978 a_2289_5307# a_2706_5417# 0.06611f
C979 a_4837_16089# a_4905_12113# 0
C980 a_14432_4521# a_13186_4919# 0
C981 a_11147_11911# a_10869_11939# 0.11706f
C982 a_4915_10549# a_8193_13753# 0.14293f
C983 a_5851_13769# a_4913_13781# 0.00386f
C984 a_9501_13813# a_9379_14779# 0.00144f
C985 a_11411_5471# a_13473_5459# 0
C986 a_24241_14651# a_24774_14701# 0.0098f
C987 a_2259_2047# a_2145_1791# 0
C988 a_16583_4529# a_16454_4503# 0.00758f
C989 VDPWR a_9579_12145# 0.00297f
C990 a_12281_1793# a_12017_1793# 0
C991 a_6261_5409# sky130_fd_sc_hd__mux4_1_0.A3 0
C992 a_12950_5459# a_12533_5715# 0.03016f
C993 a_10385_4963# a_10499_4853# 0
C994 a_12769_4809# a_12655_4553# 0
C995 a_2343_5417# a_2079_5417# 0
C996 a_4213_5409# a_2217_5025# 0
C997 a_11147_11911# a_10841_12931# 0
C998 a_12655_4553# a_12823_4553# 0
C999 a_14771_4803# a_17210_4529# 0
C1000 a_4423_5299# a_4309_5409# 0
C1001 a_5269_1787# a_4746_1787# 0
C1002 a_10525_5471# sky130_fd_sc_hd__mux4_1_0.A3 0
C1003 a_12039_15239# a_9769_15349# 0
C1004 a_3938_1787# a_2259_2047# 0
C1005 a_14771_4803# a_16402_4529# 0
C1006 a_12113_2159# a_12227_2049# 0
C1007 a_12194_5433# a_12142_5459# 0.1439f
C1008 a_4763_14775# a_4503_16339# 0
C1009 a_9317_5049# a_11439_4597# 0.04098f
C1010 a_6335_2153# a_6281_2043# 0.03622f
C1011 a_9501_13813# a_9587_13813# 0.00658f
C1012 a_4840_5043# a_2217_5025# 0
C1013 VDPWR a_14825_4547# 0.18753f
C1014 a_6717_15235# a_6635_15235# 0.00578f
C1015 a_10955_11939# a_11147_11911# 0
C1016 VDPWR sky130_fd_sc_hd__mux4_1_0.A3 0.64914f
C1017 a_4847_14525# a_6087_14735# 0.31937f
C1018 a_10916_4597# a_11439_4597# 0
C1019 a_6329_12927# a_4913_13781# 0.02039f
C1020 a_10108_4597# sky130_fd_sc_hd__mux4_1_0.A3 0
C1021 a_10499_4853# a_10525_5471# 0
C1022 a_6281_2043# a_7944_1767# 0.0035f
C1023 a_12559_4553# a_12823_4553# 0
C1024 a_13969_2159# VDPWR 0
C1025 a_6021_13769# a_4913_13781# 0.00104f
C1026 VDPWR a_12644_2159# 0.02101f
C1027 sky130_fd_sc_hd__mux4_1_0.A1 a_9703_16093# 0
C1028 a_17425_5473# sky130_fd_sc_hd__mux4_1_0.A3 0.00921f
C1029 a_13840_1767# a_14233_2159# 0.02301f
C1030 a_9779_13785# a_9379_14779# 0
C1031 a_4084_5017# a_3229_5051# 0.11874f
C1032 VDPWR a_10499_4853# 0.71231f
C1033 a_2313_2157# a_2676_2157# 0.00847f
C1034 a_11411_5471# a_9317_5049# 0.05343f
C1035 a_9781_10553# sky130_fd_sc_hd__mux4_1_0.A1 0.15936f
C1036 a_4635_13809# a_4913_13781# 0.12049f
C1037 a_6717_15235# a_7173_15235# 0
C1038 a_12559_4919# a_12823_4919# 0
C1039 a_8700_1793# a_8283_2049# 0.03016f
C1040 a_12769_4809# a_12655_4919# 0
C1041 a_3990_1761# a_4383_1787# 0.02283f
C1042 a_8337_1793# a_8169_1793# 0
C1043 a_12823_4919# a_11439_4597# 0.04534f
C1044 a_4723_10577# a_4915_10549# 0
C1045 VDPWR a_12378_4553# 0.15193f
C1046 a_15431_5467# a_15242_5833# 0
C1047 a_6335_1787# a_6281_2043# 0.00386f
C1048 a_4423_5299# a_2217_5025# 0.00303f
C1049 a_5174_5043# a_2217_5025# 0
C1050 a_7113_13395# a_6281_11907# 0.19568f
C1051 VDPWR a_16297_1793# 0.18609f
C1052 sky130_fd_sc_hd__mux4_1_0.A2 a_8169_1793# 0
C1053 a_8167_5415# a_8038_5023# 0.00792f
C1054 a_9779_13785# a_9587_13813# 0.00222f
C1055 uio_oe[7] uio_oe[6] 0.03102f
C1056 a_13167_1793# a_14233_2159# 0.04534f
C1057 a_16485_5729# a_16371_5839# 0
C1058 VDPWR a_12697_14007# 0
C1059 a_10289_1793# a_10652_1793# 0.00985f
C1060 a_24152_14385# ui_in[1] 0.02237f
C1061 a_9223_1793# a_7221_1787# 0
C1062 a_14561_4547# a_13709_4553# 0
C1063 a_6911_15235# a_4837_16089# 0.00241f
C1064 a_14771_4803# a_13709_4553# 0.21188f
C1065 a_10953_14739# a_9769_15349# 0
C1066 a_14545_5467# sky130_fd_sc_hd__mux4_1_0.A3 0
C1067 a_16094_5473# a_16275_5839# 0
C1068 a_2259_2047# VDPWR 0.44967f
C1069 a_6281_11907# a_5975_12927# 0
C1070 a_15119_1793# a_14930_2159# 0
C1071 VDPWR a_16679_4529# 0.00101f
C1072 a_16847_4529# a_16454_4503# 0.02283f
C1073 a_12587_5459# a_14152_5441# 0
C1074 a_21506_16181# a_19510_16177# 0
C1075 VDPWR a_6281_2043# 0.45202f
C1076 a_4903_15345# a_6127_13769# 0
C1077 a_7113_13395# a_9501_13813# 0
C1078 a_12587_5825# a_12323_5825# 0
C1079 a_10357_5471# a_10132_5445# 0.00487f
C1080 sky130_fd_sc_hd__mux4_1_0.A2 a_10025_1793# 0
C1081 a_21506_16181# VDPWR 0.4426f
C1082 a_4746_1787# a_4329_2043# 0.03016f
C1083 sky130_fd_sc_hd__mux4_1_0.A2 a_8700_2159# 0
C1084 a_16243_2049# a_16660_1793# 0.03016f
C1085 a_14432_4521# a_14561_4547# 0.00758f
C1086 a_14771_4803# a_14432_4521# 0.04737f
C1087 a_4913_13781# a_5933_13769# 0
C1088 a_5269_1787# sky130_fd_sc_hd__mux4_1_0.A2 0.00234f
C1089 a_1868_1791# a_2187_1765# 0.0073f
C1090 VDPWR a_6944_13645# 0.0014f
C1091 VDPWR a_4765_11543# 0.33144f
C1092 a_3990_1761# a_4215_2153# 0.00559f
C1093 a_12281_1793# a_11888_1767# 0.02283f
C1094 a_12194_5433# a_10471_5727# 0.00291f
C1095 a_9769_15349# a_9703_16093# 0.50558f
C1096 a_4084_5017# a_4309_5409# 0.00559f
C1097 a_9619_16343# a_8193_13753# 0
C1098 a_9896_1767# a_10289_1793# 0.02283f
C1099 uio_out[6] uio_out[5] 0.03102f
C1100 a_5269_1787# a_6071_1787# 0
C1101 a_9705_12861# a_9629_14779# 0.00187f
C1102 sky130_fd_sc_hd__mux4_1_0.A2 a_12655_4553# 0
C1103 sky130_fd_sc_hd__mux4_1_0.A2 a_15522_4547# 0
C1104 a_14908_5467# a_13709_4553# 0
C1105 a_9317_5049# a_18625_4938# 0.31816f
C1106 sky130_fd_sc_hd__mux4_1_0.A2 ui_in[0] 0.0357f
C1107 a_4913_13781# a_6003_11935# 0
C1108 a_6335_2153# a_6698_2153# 0.00847f
C1109 a_10953_14739# a_12039_15239# 0.00407f
C1110 sky130_fd_sc_hd__mux4_1_0.A2 a_15852_1793# 0.00174f
C1111 a_4635_13809# a_4721_13809# 0.00658f
C1112 a_11501_15239# a_12039_15239# 0.08446f
C1113 a_8073_1793# a_7221_1787# 0
C1114 a_10675_14767# a_9713_14529# 0.00178f
C1115 a_6635_15235# a_6805_15235# 0.00167f
C1116 a_12039_15239# a_11777_15239# 0
C1117 a_6261_5409# a_6036_5017# 0.00559f
C1118 a_4515_11543# a_4915_10549# 0
C1119 sky130_fd_sc_hd__mux4_1_0.A2 a_14561_4547# 0
C1120 a_13473_5459# sky130_fd_sc_hd__mux4_1_0.A3 0.00209f
C1121 sky130_fd_sc_hd__mux4_1_0.A2 a_14771_4803# 0
C1122 sky130_fd_sc_hd__mux4_1_0.A3 a_14152_5441# 0.0052f
C1123 a_14657_4547# a_13709_4553# 0
C1124 a_9493_12145# a_4915_10549# 0.00128f
C1125 sky130_fd_sc_hd__mux4_1_0.A3 a_23677_14701# 0
C1126 a_2343_5051# a_2217_5025# 0.0842f
C1127 a_7113_13395# a_5851_13769# 0
C1128 VDPWR a_12587_5825# 0.01034f
C1129 a_7315_5043# a_8167_5049# 0
C1130 VDPWR a_7927_14003# 0
C1131 a_12017_2159# a_11888_1767# 0.00792f
C1132 a_6281_11907# a_4905_12113# 0.03573f
C1133 a_24241_14651# sky130_fd_sc_hd__mux4_1_0.A3 0.03341f
C1134 sky130_fd_sc_hd__mux4_1_0.A2 a_12559_4553# 0
C1135 a_12039_15239# a_9703_16093# 0.04818f
C1136 VDPWR a_15242_5833# 0
C1137 VDPWR a_4627_12141# 0.44464f
C1138 a_10553_4963# sky130_fd_sc_hd__mux4_1_0.A3 0
C1139 a_9781_10553# a_12039_15239# 0.09278f
C1140 a_7749_14003# a_8193_13753# 0.10797f
C1141 a_4903_15345# a_4711_15373# 0.00101f
C1142 VDPWR a_6036_5017# 0.35183f
C1143 a_2313_2157# a_1920_1765# 0.02301f
C1144 a_5851_13769# a_5975_12927# 0
C1145 a_4839_12857# a_6389_13769# 0.04676f
C1146 a_12769_4809# a_12823_4553# 0.00386f
C1147 a_7173_15235# a_6805_15235# 0
C1148 a_4847_14525# a_6635_15235# 0.17821f
C1149 a_14432_4521# a_14657_4547# 0.00487f
C1150 a_4084_5017# a_2217_5025# 0.0021f
C1151 a_9629_14529# a_9769_15349# 0
C1152 a_10385_4963# a_10160_4571# 0.00559f
C1153 a_4839_12857# a_4837_16089# 0.4639f
C1154 VDPWR a_4903_15345# 0.40883f
C1155 a_7999_14003# a_8193_13753# 0
C1156 a_10289_2159# a_10025_2159# 0
C1157 VDPWR a_8794_5049# 0.21794f
C1158 a_4477_5043# a_3229_5051# 0.08312f
C1159 a_16902_5473# a_16485_5729# 0.03016f
C1160 a_10499_4853# a_10553_4963# 0.03622f
C1161 a_4755_12857# VDPWR 0.00415f
C1162 a_7113_13395# a_6329_12927# 0
C1163 a_6629_15387# a_6389_13769# 0
C1164 VDPWR a_14596_2159# 0.02101f
C1165 VDPWR a_10887_13773# 0
C1166 a_10888_5471# a_10525_5471# 0.00985f
C1167 a_9844_1793# a_9223_1793# 0.05218f
C1168 a_9621_13111# a_4915_10549# 0
C1169 a_6629_15387# a_4837_16089# 0.26097f
C1170 ui_in[1] a_23677_14335# 0
C1171 VDPWR a_9771_12117# 0.45645f
C1172 a_9317_5049# sky130_fd_sc_hd__mux4_1_0.A3 0.02471f
C1173 sky130_fd_sc_hd__mux4_1_0.A2 a_14657_4547# 0
C1174 a_4423_5299# a_4840_5043# 0.03016f
C1175 a_8700_1793# VDPWR 0.21796f
C1176 VDPWR a_6698_2153# 0.02101f
C1177 a_4847_14525# a_7173_15235# 0
C1178 a_14908_5833# a_14419_5441# 0.03325f
C1179 a_10953_14739# a_11501_15239# 0.08698f
C1180 a_2175_5051# a_2343_5051# 0
C1181 a_10888_5471# VDPWR 0.21774f
C1182 a_10953_14739# a_11777_15239# 0.00651f
C1183 a_12978_1793# VDPWR 0
C1184 a_6329_12927# a_5975_12927# 0.09582f
C1185 a_9463_11547# a_4915_10549# 0
C1186 a_11501_15239# a_11777_15239# 0.00119f
C1187 VDPWR a_10160_4571# 0.4471f
C1188 sky130_fd_sc_hd__mux4_1_0.A1 a_9619_16343# 0
C1189 a_10499_4853# a_9317_5049# 0
C1190 a_4847_14525# a_4913_13781# 0.0012f
C1191 a_6429_5043# a_8038_5023# 0
C1192 a_10160_4571# a_10108_4597# 0.1439f
C1193 a_2175_5417# a_2217_5025# 0
C1194 VDPWR a_10121_1793# 0
C1195 a_12769_4809# a_13709_4553# 0.13741f
C1196 VDPWR a_12950_5459# 0.21529f
C1197 a_24407_14651# a_24774_14701# 0
C1198 sky130_fd_sc_hd__mux4_1_0.A2 a_14179_2049# 0.00304f
C1199 a_10953_14739# a_9703_16093# 0.29394f
C1200 a_10499_4853# a_10916_4597# 0.03016f
C1201 a_12823_4919# sky130_fd_sc_hd__mux4_1_0.A3 0
C1202 a_10553_4597# a_10499_4853# 0.00386f
C1203 a_11501_15239# a_9703_16093# 0.23067f
C1204 VDPWR a_6165_5043# 0.00122f
C1205 a_6281_11907# a_9371_13111# 0
C1206 a_10525_5471# a_8377_5305# 0
C1207 uio_out[4] uio_out[5] 0.03102f
C1208 a_11777_15239# a_9703_16093# 0.00241f
C1209 a_24234_14385# sky130_fd_sc_hd__mux4_1_0.A2 0.04346f
C1210 a_23511_14701# sky130_fd_sc_hd__mux4_1_0.A3 0.00138f
C1211 a_16146_5447# sky130_fd_sc_hd__mux4_1_0.A3 0.00525f
C1212 a_5363_5043# a_5174_5409# 0
C1213 a_5174_5043# a_4423_5299# 0.00682f
C1214 a_12769_4809# a_14432_4521# 0.00352f
C1215 VDPWR a_11979_13399# 0.501f
C1216 VDPWR a_8377_5305# 0.45194f
C1217 a_18742_16187# a_19510_16177# 0.1036f
C1218 sky130_fd_sc_hd__mux4_1_0.A2 a_10986_2159# 0
C1219 a_10108_4597# a_8377_5305# 0
C1220 a_2289_5307# a_2706_5051# 0.03016f
C1221 a_5269_1787# a_2187_1765# 0.00133f
C1222 a_16679_4895# a_17733_4529# 0
C1223 a_18742_16187# VDPWR 0.4418f
C1224 a_11147_11911# a_11728_13649# 0.00254f
C1225 a_11255_13773# a_12615_14007# 0.00184f
C1226 uio_oe[4] uio_oe[3] 0.03102f
C1227 VDPWR a_12113_2159# 0
C1228 a_9781_10553# a_9703_16093# 0.01618f
C1229 a_9501_13813# a_9371_13111# 0.00115f
C1230 sky130_fd_sc_hd__mux4_1_0.A2 a_17210_4529# 0
C1231 VDPWR a_10717_13773# 0.4459f
C1232 a_2187_1765# a_5890_1787# 0.00121f
C1233 sky130_fd_sc_hd__mux4_1_0.A2 a_16402_4529# 0
C1234 VDPWR a_12865_14007# 0
C1235 a_24774_14701# a_24962_14701# 0.10432f
C1236 a_2343_5417# a_1950_5025# 0.02301f
C1237 a_6261_5409# a_6375_5299# 0
C1238 a_12769_4809# sky130_fd_sc_hd__mux4_1_0.A2 0
C1239 a_11195_12931# a_10841_12931# 0.09582f
C1240 sky130_fd_sc_hd__mux4_1_0.A2 a_12823_4553# 0
C1241 a_14419_5441# a_14377_5467# 0
C1242 a_4119_1787# a_3199_1791# 0
C1243 VDPWR a_3040_5051# 0
C1244 a_7032_1787# a_6281_2043# 0.00682f
C1245 a_11195_12931# a_9371_13111# 0
C1246 a_10235_2049# a_10121_1793# 0
C1247 a_5984_5043# a_2217_5025# 0.00121f
C1248 a_9779_13785# a_10995_12931# 0
C1249 a_4084_5017# a_4213_5409# 0.00792f
C1250 a_9779_13785# a_10869_11939# 0
C1251 a_16033_2159# a_15852_1793# 0
C1252 VDPWR a_4597_11543# 0.02518f
C1253 a_5080_1787# VDPWR 0
C1254 VDPWR a_4513_14775# 0.51083f
C1255 a_6003_11935# a_5975_12927# 0
C1256 a_16371_5473# a_15431_5467# 0
C1257 VDPWR a_6375_5299# 0.4517f
C1258 a_4477_5043# a_2217_5025# 0
C1259 a_10525_5471# a_10132_5445# 0.02283f
C1260 a_9779_13785# a_10841_12931# 0.08477f
C1261 a_9713_14529# a_11583_15239# 0.00159f
C1262 a_4746_2153# a_2187_1765# 0
C1263 VDPWR a_4383_2153# 0.0097f
C1264 sky130_fd_sc_hd__mux4_1_0.A2 a_16129_1793# 0
C1265 a_4213_5043# a_3229_5051# 0
C1266 a_9781_10553# a_4915_10549# 0.00418f
C1267 a_14432_4521# a_13709_4553# 0.11874f
C1268 VDPWR a_11222_5471# 0
C1269 VDPWR a_10132_5445# 0.35088f
C1270 a_9779_13785# a_9371_13111# 0
C1271 a_13840_1767# a_13969_1793# 0.00758f
C1272 a_10108_4597# a_10132_5445# 0
C1273 a_7986_5049# a_8038_5023# 0.1439f
C1274 a_15904_1767# a_16297_1793# 0.02283f
C1275 a_12323_5459# a_11411_5471# 0
C1276 a_2259_2047# a_2313_2157# 0.03622f
C1277 a_10499_4853# a_11250_4597# 0.00682f
C1278 a_15242_5467# sky130_fd_sc_hd__mux4_1_0.A3 0
C1279 a_4839_12857# a_6281_11907# 0.02321f
C1280 a_7315_5043# a_7126_5409# 0
C1281 a_8167_5415# a_8431_5415# 0
C1282 a_9379_14779# a_9629_14779# 0.02504f
C1283 a_16539_5473# sky130_fd_sc_hd__mux4_1_0.A3 0
C1284 a_10525_5471# a_10261_5471# 0
C1285 a_6089_11935# a_4915_10549# 0
C1286 a_12950_5459# a_14152_5441# 0
C1287 sky130_fd_sc_hd__mux4_1_0.A2 a_13709_4553# 0
C1288 a_13473_5459# a_12950_5459# 0
C1289 a_4505_13107# VDPWR 0.51474f
C1290 VDPWR a_10986_1793# 0
C1291 a_4032_5043# a_3229_5051# 0.05073f
C1292 a_4423_5299# a_4084_5017# 0.04737f
C1293 a_18839_4938# a_17733_4529# 0
C1294 a_13167_1793# a_13969_1793# 0
C1295 a_8794_5049# a_9317_5049# 0
C1296 a_7032_2153# a_7221_1787# 0
C1297 a_15711_4547# sky130_fd_sc_hd__mux4_1_0.A3 0
C1298 a_10160_4571# a_10553_4963# 0.02301f
C1299 a_2187_1765# a_4329_2043# 0.00305f
C1300 VDPWR a_10261_5471# 0.00116f
C1301 VDPWR a_16583_4895# 0
C1302 a_5363_5043# a_6261_5043# 0
C1303 a_6003_11935# a_4905_12113# 0.18489f
C1304 VDPWR a_8193_13753# 2.59438f
C1305 a_9629_14529# a_4915_10549# 0
C1306 VDPWR a_3229_5051# 1.42184f
C1307 a_6629_15387# a_4753_16339# 0
C1308 a_5942_1761# a_6167_1787# 0.00487f
C1309 a_10385_4597# VDPWR 0.00132f
C1310 sky130_fd_sc_hd__mux4_1_0.A2 a_14432_4521# 0
C1311 a_7221_1787# a_8283_2049# 0.21187f
C1312 a_2259_2047# a_3990_1761# 0.00332f
C1313 VDPWR a_4713_12141# 0.00297f
C1314 sky130_fd_sc_hd__mux4_1_0.A2 a_16033_1793# 0
C1315 uio_out[1] uio_out[0] 0.03102f
C1316 a_23511_14335# ui_in[0] 0.01792f
C1317 a_5363_5043# a_7315_5043# 0
C1318 a_11836_1793# a_12017_2159# 0
C1319 sky130_fd_sc_hd__mux4_1_0.A3 a_9128_5415# 0
C1320 a_8337_2159# a_8283_2049# 0.03622f
C1321 a_24407_14651# sky130_fd_sc_hd__mux4_1_0.A3 0
C1322 a_15431_5467# a_16539_5839# 0.04534f
C1323 a_4903_15345# a_6087_14735# 0
C1324 sky130_fd_sc_hd__mux4_1_0.A2 a_8337_1793# 0
C1325 a_8377_5305# a_10553_4963# 0
C1326 a_10121_2159# VDPWR 0
C1327 VDPWR a_10993_13773# 0.0014f
C1328 a_10160_4571# a_9317_5049# 0
C1329 VDPWR ua[4] 0.00173f
C1330 a_10289_2159# VDPWR 0.00967f
C1331 a_4753_16089# a_4837_16089# 0.00234f
C1332 VDPWR a_13520_4919# 0
C1333 VDPWR a_14561_4913# 0
C1334 a_9621_12861# a_9371_13111# 0.00723f
C1335 a_16679_4895# VDPWR 0
C1336 a_18742_16187# a_17254_16187# 0
C1337 uo_out[6] uo_out[7] 0.03102f
C1338 a_10553_4597# a_10160_4571# 0.02283f
C1339 VDPWR a_16371_5473# 0
C1340 a_9713_14529# a_9501_13813# 0
C1341 a_16847_4895# a_17733_4529# 0
C1342 a_6389_13769# a_4837_16089# 0.00515f
C1343 a_17210_4529# a_16485_5729# 0
C1344 a_9844_1793# a_10025_2159# 0
C1345 a_14419_5441# a_14491_5723# 0.21187f
C1346 a_4839_12857# a_5851_13769# 0.13054f
C1347 a_10235_2049# a_10986_1793# 0.00682f
C1348 a_16793_4785# a_17210_4529# 0.03016f
C1349 uio_in[5] uio_in[6] 0.03102f
C1350 VDPWR a_14825_4913# 0.01165f
C1351 a_9317_5049# a_8377_5305# 0.13758f
C1352 a_8038_5023# sky130_fd_sc_hd__mux4_1_0.A3 0.00209f
C1353 VDPWR a_15119_1793# 1.40147f
C1354 a_10887_13773# a_9705_12861# 0
C1355 a_10121_1793# a_9896_1767# 0.00487f
C1356 a_5895_14763# VDPWR 0
C1357 a_15711_4547# a_16679_4529# 0
C1358 a_2676_1791# a_2187_1765# 0.08982f
C1359 ui_in[1] a_23731_14309# 0.35239f
C1360 a_4723_10577# VDPWR 0.00176f
C1361 a_12644_1793# a_13167_1793# 0
C1362 a_9705_12861# a_9771_12117# 0.04364f
C1363 ui_in[1] a_24318_14385# 0.04767f
C1364 VDPWR a_10525_5837# 0.00694f
C1365 a_9619_16343# a_9703_16093# 0.07445f
C1366 a_14908_5833# sky130_fd_sc_hd__mux4_1_0.A3 0.0019f
C1367 a_4625_15373# a_4711_15373# 0.00658f
C1368 a_16902_5839# a_15431_5467# 0.03325f
C1369 a_16847_4529# a_14771_4803# 0
C1370 a_12323_5459# a_12587_5459# 0
C1371 a_4213_5043# a_2217_5025# 0
C1372 a_9629_14779# a_9369_16343# 0
C1373 VDPWR a_4309_5409# 0
C1374 a_4746_1787# a_2187_1765# 0
C1375 a_4477_5043# a_4840_5043# 0.00985f
C1376 a_2187_1765# a_3010_1791# 0
C1377 a_6792_5043# a_7315_5043# 0
C1378 VDPWR a_4625_15373# 0.45068f
C1379 a_16243_2049# a_16297_1793# 0.00386f
C1380 a_8263_5415# sky130_fd_sc_hd__mux4_1_0.A3 0
C1381 a_17210_4895# sky130_fd_sc_hd__mux4_1_0.A3 0
C1382 a_3938_1787# a_3199_1791# 0.05108f
C1383 ui_in[4] ui_in[5] 0.03102f
C1384 a_19510_16177# sky130_fd_sc_hd__mux4_1_0.A1 0
C1385 a_4839_12857# a_6329_12927# 0.08252f
C1386 a_10235_2049# a_10121_2159# 0
C1387 a_7221_1787# a_7944_1767# 0.11881f
C1388 a_9779_13785# a_9713_14529# 0.0012f
C1389 uio_in[7] uo_out[0] 0.03102f
C1390 a_13969_2159# a_13840_1767# 0.00792f
C1391 a_9491_15377# a_8193_13753# 0
C1392 a_10289_2159# a_10235_2049# 0.03622f
C1393 a_4839_12857# a_6021_13769# 0
C1394 VDPWR sky130_fd_sc_hd__mux4_1_0.A1 1.6285f
C1395 a_8337_2159# a_7944_1767# 0.02301f
C1396 a_2289_5307# a_1950_5025# 0.04737f
C1397 a_4032_5043# a_2217_5025# 0.00121f
C1398 a_6862_13645# a_4915_10549# 0
C1399 a_4423_5299# a_5984_5043# 0
C1400 a_4839_12857# a_4635_13809# 0.00246f
C1401 VDPWR a_16539_5839# 0.01025f
C1402 a_12323_5459# sky130_fd_sc_hd__mux4_1_0.A3 0
C1403 VDPWR a_5809_14763# 0.21213f
C1404 VDPWR ui_in[1] 0.45013f
C1405 a_9705_12861# a_11979_13399# 0.00446f
C1406 a_9844_1793# a_8283_2049# 0
C1407 a_14281_5833# a_14100_5467# 0
C1408 a_4215_1787# a_3199_1791# 0
C1409 a_4477_5043# a_4423_5299# 0.00386f
C1410 VDPWR a_15188_4913# 0.02568f
C1411 a_4627_12141# a_4755_13107# 0
C1412 a_9317_5049# a_10132_5445# 0
C1413 a_16454_4503# sky130_fd_sc_hd__mux4_1_0.A3 0
C1414 VDPWR a_2217_5025# 1.58075f
C1415 a_12430_4527# a_12655_4553# 0.00487f
C1416 a_4585_16339# a_4503_16339# 0.00641f
C1417 VDPWR a_18839_4938# 0.00182f
C1418 sky130_fd_sc_hd__mux4_1_0.A3 a_13284_5825# 0
C1419 ui_in[0] rst_n 0.03102f
C1420 VDPWR a_2145_2157# 0
C1421 a_9705_12861# a_10717_13773# 0.13054f
C1422 a_7113_13395# a_7831_14003# 0.00223f
C1423 a_4513_14775# a_6087_14735# 0
C1424 a_4309_5043# a_3229_5051# 0
C1425 VDPWR a_4515_11543# 0.50586f
C1426 a_14179_2049# a_14233_2159# 0.03622f
C1427 VDPWR a_7221_1787# 1.41106f
C1428 a_9223_1793# a_8283_2049# 0.13739f
C1429 a_14377_5467# sky130_fd_sc_hd__mux4_1_0.A3 0
C1430 VDPWR a_9493_12145# 0.44464f
C1431 ua[0] a_23731_14309# 0
C1432 a_12430_4527# a_12559_4553# 0.00758f
C1433 VDPWR a_8337_2159# 0.0097f
C1434 a_11411_5471# a_12950_5825# 0.03325f
C1435 a_7749_14003# a_4915_10549# 0.07615f
C1436 a_12113_2159# a_11888_1767# 0.00559f
C1437 a_5269_1787# a_6698_1787# 0.08907f
C1438 a_13186_4919# a_11439_4597# 0.03325f
C1439 VDPWR a_4503_16339# 0.5096f
C1440 VDPWR a_3199_1791# 1.41762f
C1441 VDPWR a_16902_5839# 0.01944f
C1442 a_9451_16343# a_9703_16093# 0
C1443 a_11255_13773# a_9713_14529# 0
C1444 a_11195_12931# a_11728_13649# 0.10646f
C1445 a_4839_12857# a_5933_13769# 0
C1446 VDPWR a_9769_15349# 0.40883f
C1447 VDPWR a_14657_4913# 0
C1448 a_7999_14003# a_4915_10549# 0
C1449 sky130_fd_sc_hd__mux4_1_0.A2 a_2187_1765# 0.11803f
C1450 a_6071_2153# a_5890_1787# 0
C1451 a_12430_4527# a_12655_4919# 0.00559f
C1452 a_6071_1787# a_2187_1765# 0
C1453 uo_out[3] uo_out[4] 0.03102f
C1454 sky130_fd_sc_hd__mux4_1_0.A2 a_16660_2159# 0.00205f
C1455 a_1868_1791# a_1920_1765# 0.1439f
C1456 a_4839_12857# a_6003_11935# 0
C1457 sky130_fd_sc_hd__mux4_1_0.A2 a_16793_4785# 0
C1458 a_8794_5415# sky130_fd_sc_hd__mux4_1_0.A3 0
C1459 VDPWR a_16847_4895# 0.01197f
C1460 a_2706_5417# a_2217_5025# 0.0357f
C1461 VDPWR a_2175_5051# 0.00105f
C1462 a_11411_5471# a_13186_4919# 0
C1463 a_11810_13649# a_11979_13399# 0
C1464 a_10553_4597# a_10385_4597# 0
C1465 a_12769_4809# a_14380_4547# 0
C1466 a_16454_4503# a_16679_4529# 0.00487f
C1467 sky130_fd_sc_hd__mux4_1_0.A2 a_12978_2159# 0
C1468 a_4903_15345# a_7173_15235# 0
C1469 a_9779_13785# a_11728_13649# 0
C1470 a_16847_4529# a_17210_4529# 0.00985f
C1471 VDPWR a_9621_13111# 0.33272f
C1472 sky130_fd_sc_hd__mux4_1_0.A2 a_16033_2159# 0
C1473 uio_out[2] uio_out[1] 0.03102f
C1474 a_10888_5837# a_10471_5727# 0.06611f
C1475 a_6281_11907# a_6389_13769# 0.00254f
C1476 a_15119_1793# a_14596_1793# 0
C1477 a_4477_5409# a_4840_5409# 0.00847f
C1478 VDPWR a_10916_4963# 0.05811f
C1479 VDPWR a_12039_15239# 0.7104f
C1480 a_11195_12931# a_11147_11911# 0.00298f
C1481 sky130_fd_sc_hd__mux4_1_0.A3 a_10357_5837# 0
C1482 a_10717_13773# a_10799_13773# 0.00578f
C1483 a_4903_15345# a_4913_13781# 0.11595f
C1484 a_9589_10581# a_9781_10553# 0
C1485 VDPWR ua[0] 0.20284f
C1486 sky130_fd_sc_hd__mux4_1_0.A1 a_23677_14701# 0
C1487 a_9779_13785# a_10675_14767# 0
C1488 sky130_fd_sc_hd__mux4_1_0.A2 a_16994_2159# 0
C1489 a_4763_14775# VDPWR 0.33336f
C1490 a_9463_11547# VDPWR 0.02518f
C1491 a_10121_2159# a_9896_1767# 0.00559f
C1492 a_5363_5043# a_6792_5043# 0.08907f
C1493 a_10289_2159# a_9896_1767# 0.02301f
C1494 a_12419_5825# sky130_fd_sc_hd__mux4_1_0.A3 0
C1495 a_4753_16339# a_4837_16089# 0.07445f
C1496 a_9223_1793# a_11175_1793# 0
C1497 a_3990_1761# a_4383_2153# 0.02301f
C1498 a_4477_5043# a_4084_5017# 0.02283f
C1499 sky130_fd_sc_hd__mux4_1_0.A2 a_16583_4529# 0
C1500 a_6335_2153# a_5942_1761# 0.02301f
C1501 a_4032_5043# a_4213_5409# 0
C1502 a_9705_12861# a_8193_13753# 0.00341f
C1503 a_14771_4803# a_14419_5441# 0
C1504 a_17254_16187# sky130_fd_sc_hd__mux4_1_0.A1 0
C1505 VDPWR a_8431_5049# 0.18611f
C1506 a_11411_5471# a_12142_5459# 0.05122f
C1507 a_8377_5305# a_9128_5415# 0.00696f
C1508 ui_in[1] a_23677_14701# 0.0594f
C1509 a_24241_14651# ui_in[1] 0.00168f
C1510 VDPWR a_4213_5409# 0
C1511 a_16146_5447# a_16371_5473# 0.00487f
C1512 a_12194_5433# a_12419_5459# 0.00487f
C1513 sky130_fd_sc_hd__mux4_1_0.A3 a_16371_5839# 0
C1514 sky130_fd_sc_hd__mux4_1_0.A2 a_12281_2159# 0
C1515 a_14380_4547# a_13709_4553# 0.05169f
C1516 a_9705_12861# a_10993_13773# 0.00253f
C1517 a_5895_14763# a_6087_14735# 0
C1518 a_13788_1793# a_12227_2049# 0
C1519 a_12655_4553# a_11439_4597# 0
C1520 a_9844_1793# VDPWR 0.13948f
C1521 VDPWR a_4840_5043# 0.21798f
C1522 a_14419_5441# a_14908_5467# 0.08907f
C1523 VDPWR a_11222_5837# 0
C1524 a_4513_14775# a_4755_13107# 0
C1525 a_5942_1761# a_6335_1787# 0.02283f
C1526 a_4309_5043# a_2217_5025# 0
C1527 a_9491_15377# a_9769_15349# 0.12165f
C1528 a_11255_13773# a_11728_13649# 0.24537f
C1529 a_14930_1793# ua[4] 0
C1530 a_14596_2159# a_13167_1793# 0.03325f
C1531 a_24152_14385# a_23731_14309# 0.01881f
C1532 a_24152_14385# a_24318_14385# 0.05583f
C1533 a_8377_5305# a_8038_5023# 0.04737f
C1534 a_4383_1787# a_4329_2043# 0.00386f
C1535 a_14491_5723# sky130_fd_sc_hd__mux4_1_0.A3 0.00768f
C1536 a_4839_12857# a_4847_14525# 0.18435f
C1537 a_14432_4521# a_14380_4547# 0.1439f
C1538 VDPWR a_10953_14739# 0.4457f
C1539 a_4839_12857# a_4763_14525# 0
C1540 a_9577_15377# a_9769_15349# 0.00101f
C1541 a_12769_4809# a_12430_4527# 0.04737f
C1542 a_5851_13769# a_6389_13769# 0.07901f
C1543 a_8073_1793# a_7944_1767# 0.00758f
C1544 VDPWR a_11501_15239# 0.4212f
C1545 ui_in[0] a_24774_14701# 0.02515f
C1546 a_18625_5265# a_17733_4529# 0.00499f
C1547 a_12430_4527# a_12823_4553# 0.02283f
C1548 a_5851_13769# a_4837_16089# 0.08387f
C1549 VDPWR a_11777_15239# 0
C1550 VDPWR a_16297_2159# 0.00966f
C1551 a_6261_5409# a_6429_5409# 0
C1552 a_12559_4553# a_11439_4597# 0
C1553 VDPWR a_9223_1793# 1.41077f
C1554 a_18839_4938# a_9317_5049# 0.00688f
C1555 a_6629_15387# a_4847_14525# 0.29211f
C1556 a_6944_13645# a_7113_13395# 0
C1557 a_4423_5299# VDPWR 0.45138f
C1558 a_5942_1761# VDPWR 0.35292f
C1559 a_8263_5415# a_8377_5305# 0
C1560 a_5174_5043# VDPWR 0
C1561 a_12615_14007# a_12697_14007# 0.00695f
C1562 a_12950_5825# sky130_fd_sc_hd__mux4_1_0.A3 0.00186f
C1563 sky130_fd_sc_hd__mux4_1_0.A2 a_14380_4547# 0
C1564 a_4505_13107# a_4755_13107# 0.02504f
C1565 a_11255_13773# a_11147_11911# 0.00254f
C1566 VDPWR a_9703_16093# 1.40253f
C1567 a_23511_14701# sky130_fd_sc_hd__mux4_1_0.A1 0.04613f
C1568 a_10289_1793# a_10025_1793# 0
C1569 sky130_fd_sc_hd__mux4_1_0.A2 a_8073_2159# 0
C1570 sky130_fd_sc_hd__mux4_1_0.A2 a_14233_2159# 0
C1571 a_15904_1767# a_15119_1793# 0.11873f
C1572 VDPWR ua[7] 0
C1573 VDPWR a_9781_10553# 0.69476f
C1574 a_14281_5833# sky130_fd_sc_hd__mux4_1_0.A3 0
C1575 a_15431_5467# a_16275_5473# 0
C1576 a_6087_14735# a_5809_14763# 0.1109f
C1577 a_16793_4785# a_16485_5729# 0
C1578 VDPWR a_6429_5409# 0.00968f
C1579 a_8431_5415# sky130_fd_sc_hd__mux4_1_0.A3 0
C1580 a_2049_2157# VDPWR 0
C1581 sky130_fd_sc_hd__mux4_1_0.A2 a_16847_4529# 0
C1582 a_16146_5447# a_16539_5839# 0.02301f
C1583 a_6329_12927# a_6389_13769# 0.20048f
C1584 a_3229_5051# a_2706_5051# 0
C1585 a_6375_5299# a_8038_5023# 0.0035f
C1586 VDPWR a_24152_14385# 0.00498f
C1587 a_11411_5471# a_10471_5727# 0.13964f
C1588 a_4513_14775# a_4913_13781# 0
C1589 ui_in[1] a_23511_14701# 0.05408f
C1590 a_6021_13769# a_6389_13769# 0
C1591 a_10675_14767# a_10761_14767# 0.00658f
C1592 a_7113_13395# a_7927_14003# 0.00121f
C1593 sky130_fd_sc_hd__mux4_1_0.A2 a_10289_4597# 0
C1594 a_13186_4919# sky130_fd_sc_hd__mux4_1_0.A3 0
C1595 a_4329_2043# a_4215_2153# 0
C1596 ua[5] a_10986_1793# 0
C1597 a_12587_5825# a_12419_5825# 0
C1598 a_6021_13769# a_4837_16089# 0.00246f
C1599 a_10553_4963# a_10916_4963# 0.00847f
C1600 a_18846_5265# a_18625_4938# 0.00783f
C1601 a_8073_1793# VDPWR 0.00117f
C1602 a_7999_14003# a_7749_14003# 0.00876f
C1603 a_16371_5473# a_16539_5473# 0
C1604 VDPWR a_6089_11935# 0
C1605 a_4119_2153# a_2187_1765# 0
C1606 a_2313_1791# a_2676_1791# 0.00985f
C1607 VDPWR a_4587_13107# 0.0252f
C1608 a_16847_4895# a_9317_5049# 0
C1609 a_16902_5473# sky130_fd_sc_hd__mux4_1_0.A3 0
C1610 VDPWR a_4915_10549# 0.86941f
C1611 a_4084_5017# a_4213_5043# 0.00758f
C1612 a_12430_4527# a_12194_5433# 0
C1613 a_10235_2049# a_9223_1793# 0.21187f
C1614 a_4839_12857# a_4595_14775# 0
C1615 a_4746_1787# a_4383_1787# 0.00985f
C1616 VDPWR a_9629_14529# 0.00474f
C1617 a_7113_13395# a_4903_15345# 0
C1618 a_5363_5043# a_6792_5409# 0.03325f
C1619 a_6717_15235# a_4837_16089# 0
C1620 sky130_fd_sc_hd__mux4_1_0.A3 a_8263_5049# 0
C1621 a_2145_2157# a_2313_2157# 0
C1622 a_7173_15235# a_8193_13753# 0.04124f
C1623 VDPWR a_17236_5473# 0
C1624 a_10261_5837# sky130_fd_sc_hd__mux4_1_0.A3 0
C1625 a_4505_13107# a_4913_13781# 0
C1626 a_12142_5459# sky130_fd_sc_hd__mux4_1_0.A3 0.003f
C1627 a_9705_12861# a_9493_12145# 0
C1628 a_9713_14529# a_9629_14779# 0.07979f
C1629 VDPWR a_2343_5051# 0.18537f
C1630 a_15522_4913# sky130_fd_sc_hd__mux4_1_0.A3 0
C1631 a_4903_15345# a_5975_12927# 0
C1632 a_17236_5473# a_17425_5473# 0
C1633 VDPWR a_14233_1793# 0.18613f
C1634 a_6335_1787# a_6167_1787# 0
C1635 a_12194_5433# a_10888_5837# 0
C1636 a_4084_5017# a_4032_5043# 0.1439f
C1637 a_2079_5417# a_2217_5025# 0
C1638 a_20384_16179# a_22274_16171# 0
C1639 VDPWR a_14930_2159# 0
C1640 a_17236_5839# a_16485_5729# 0.00696f
C1641 a_5933_13769# a_6389_13769# 0
C1642 a_9705_12861# a_9769_15349# 0.1369f
C1643 sky130_fd_sc_hd__mux4_1_0.A2 a_12430_4527# 0
C1644 a_15242_5833# a_14491_5723# 0.00696f
C1645 a_24234_14385# a_24774_14701# 0.17579f
C1646 a_8377_5305# a_8794_5415# 0.06611f
C1647 a_12533_5715# a_14545_5833# 0
C1648 a_5933_13769# a_4837_16089# 0
C1649 VDPWR a_4084_5017# 0.35048f
C1650 a_9491_15377# a_9703_16093# 0
C1651 a_11175_1793# a_12227_2049# 0.21187f
C1652 VDPWR a_6057_12927# 0
C1653 VDPWR a_16275_5473# 0.00119f
C1654 sky130_fd_sc_hd__mux4_1_0.A2 a_16660_1793# 0.00236f
C1655 a_7126_5043# sky130_fd_sc_hd__mux4_1_0.A3 0
C1656 a_18846_5265# sky130_fd_sc_hd__mux4_1_0.A3 0.00101f
C1657 a_12769_4809# a_11439_4597# 0.21189f
C1658 a_6261_5043# a_6429_5043# 0
C1659 a_6003_11935# a_4837_16089# 0
C1660 a_12823_4553# a_11439_4597# 0.08312f
C1661 a_12587_5825# a_12950_5825# 0.00847f
C1662 a_16275_5839# sky130_fd_sc_hd__mux4_1_0.A3 0
C1663 VDPWR a_6167_1787# 0
C1664 a_4627_12141# a_4905_12113# 0.12057f
C1665 a_10471_5727# a_12587_5459# 0
C1666 a_9621_13111# a_9705_12861# 0.08134f
C1667 a_14419_5441# a_13709_4553# 0.00111f
C1668 VDPWR a_18625_5265# 0
C1669 a_15711_4547# a_16539_5839# 0
C1670 a_16243_2049# a_15119_1793# 0.21187f
C1671 a_5895_14763# a_7173_15235# 0
C1672 a_9705_12861# a_12039_15239# 0.00685f
C1673 a_10289_4963# sky130_fd_sc_hd__mux4_1_0.A3 0
C1674 ui_in[0] sky130_fd_sc_hd__mux4_1_0.A3 0.08699f
C1675 a_3990_1761# a_3199_1791# 0.11873f
C1676 VDPWR a_23677_14335# 0
C1677 a_4423_5299# a_4309_5043# 0
C1678 sky130_fd_sc_hd__mux4_1_0.A2 a_6698_1787# 0
C1679 a_18625_5265# a_17425_5473# 0.0056f
C1680 a_12769_4809# a_11411_5471# 0
C1681 a_9379_14779# a_8193_13753# 0.00206f
C1682 a_14561_4547# a_14825_4547# 0
C1683 a_5851_13769# a_6281_11907# 0
C1684 a_2217_5025# a_2706_5051# 0.08994f
C1685 a_12227_2049# a_12113_1793# 0
C1686 a_16454_4503# a_16583_4895# 0.00792f
C1687 a_14771_4803# a_14825_4547# 0.00386f
C1688 a_9223_1793# a_10652_1793# 0.08907f
C1689 a_14419_5441# a_14432_4521# 0.00135f
C1690 a_12793_14007# a_11979_13399# 0.00121f
C1691 VDPWR a_9128_5049# 0
C1692 a_9844_1793# a_9896_1767# 0.1439f
C1693 a_14771_4803# sky130_fd_sc_hd__mux4_1_0.A3 0
C1694 a_2175_5417# VDPWR 0
C1695 a_6375_5299# a_8794_5415# 0
C1696 a_9223_1793# a_9034_2159# 0
C1697 a_2706_5417# a_4084_5017# 0
C1698 a_16847_4529# a_16793_4785# 0.00386f
C1699 a_9769_15349# a_10799_13773# 0.0035f
C1700 a_8794_5415# a_10132_5445# 0
C1701 a_12615_14007# a_11979_13399# 0.27996f
C1702 a_18553_4938# a_18625_4938# 0
C1703 a_10471_5727# sky130_fd_sc_hd__mux4_1_0.A3 0.00739f
C1704 VDPWR a_6862_13645# 0.16049f
C1705 a_16486_16197# a_18128_16189# 0
C1706 a_6805_15235# a_4837_16089# 0
C1707 VDPWR a_12227_2049# 0.45076f
C1708 a_11439_4597# a_13709_4553# 0
C1709 a_9779_13785# a_9501_13813# 0.12049f
C1710 VDPWR a_9619_16343# 0.33721f
C1711 VDPWR a_4119_1787# 0.00118f
C1712 a_6329_12927# a_6281_11907# 0.00298f
C1713 a_16679_4895# a_16454_4503# 0.00559f
C1714 a_4477_5043# a_4213_5043# 0
C1715 a_12655_4919# sky130_fd_sc_hd__mux4_1_0.A3 0
C1716 a_16902_5839# a_15711_4547# 0
C1717 a_9896_1767# a_9223_1793# 0.11878f
C1718 a_14908_5467# sky130_fd_sc_hd__mux4_1_0.A3 0
C1719 a_8700_2159# a_6281_2043# 0
C1720 a_11250_4963# a_11439_4597# 0
C1721 a_7173_15235# a_5809_14763# 0
C1722 a_5269_1787# a_6281_2043# 0.21187f
C1723 a_10499_4853# a_10471_5727# 0.00177f
C1724 a_10357_5837# a_10132_5445# 0.00559f
C1725 a_12615_14007# a_10717_13773# 0
C1726 a_15119_1793# a_13167_1793# 0
C1727 a_12615_14007# a_12865_14007# 0.00876f
C1728 VDPWR a_12533_5715# 0.44177f
C1729 a_13788_1793# VDPWR 0.13948f
C1730 a_10357_5471# a_10525_5471# 0
C1731 sky130_fd_sc_hd__mux4_1_0.A2 a_9034_1793# 0
C1732 VDPWR a_13186_4553# 0.21831f
C1733 a_11195_12931# a_9779_13785# 0.02039f
C1734 a_15711_4547# a_16847_4895# 0.04534f
C1735 a_16454_4503# a_14825_4913# 0
C1736 a_14657_4547# a_14825_4547# 0
C1737 a_10953_14739# a_9705_12861# 0.02474f
C1738 ua[6] a_6281_2043# 0
C1739 a_4847_14525# a_6389_13769# 0
C1740 a_4913_13781# a_5809_14763# 0
C1741 a_4847_14525# a_4837_16089# 0.46419f
C1742 VDPWR a_10357_5471# 0
C1743 VDPWR a_10025_2159# 0
C1744 a_2289_5307# a_3040_5417# 0.00696f
C1745 a_16847_4529# a_16583_4529# 0
C1746 ui_in[1] a_24962_14701# 0.12838f
C1747 a_14233_1793# a_14065_1793# 0
C1748 a_12194_5433# a_11411_5471# 0.11876f
C1749 a_8283_2049# a_7944_1767# 0.04737f
C1750 a_10995_12931# a_9771_12117# 0
C1751 a_10869_11939# a_9771_12117# 0.18489f
C1752 a_14377_5833# a_14545_5833# 0
C1753 VDPWR a_7749_14003# 0.13676f
C1754 VDPWR a_5984_5043# 0.13952f
C1755 a_7315_5043# a_7986_5049# 0.05168f
C1756 sky130_fd_sc_hd__mux4_1_0.A2 a_11439_4597# 0.00102f
C1757 a_10289_2159# a_10652_2159# 0.00847f
C1758 a_8377_5305# a_8431_5415# 0.03622f
C1759 a_9705_12861# a_9703_16093# 0.4639f
C1760 a_4477_5043# VDPWR 0.18615f
C1761 a_10841_12931# a_9771_12117# 0
C1762 a_7999_14003# VDPWR 0
C1763 sky130_fd_sc_hd__mux4_1_0.A2 a_12281_1793# 0
C1764 a_14233_1793# a_14596_1793# 0.00985f
C1765 a_8167_5049# sky130_fd_sc_hd__mux4_1_0.A3 0
C1766 a_10080_5471# sky130_fd_sc_hd__mux4_1_0.A3 0.00331f
C1767 a_7113_13395# a_8193_13753# 0.03479f
C1768 a_8193_13753# a_9369_16343# 0.00257f
C1769 a_9705_12861# a_9781_10553# 0.00242f
C1770 a_4309_5043# a_4084_5017# 0.00487f
C1771 a_12769_4809# a_12587_5459# 0
C1772 a_4505_13107# a_5975_12927# 0
C1773 a_18553_4938# sky130_fd_sc_hd__mux4_1_0.A3 0
C1774 ui_in[2] ui_in[1] 0.03102f
C1775 a_9371_13111# a_9771_12117# 0
C1776 a_15904_1767# a_16297_2159# 0.02301f
C1777 a_24234_14385# sky130_fd_sc_hd__mux4_1_0.A3 0.07599f
C1778 a_16793_4785# a_18371_4938# 0
C1779 a_10955_11939# a_9771_12117# 0
C1780 a_2049_2157# a_2313_2157# 0
C1781 sky130_fd_sc_hd__mux4_1_0.A2 a_24774_14701# 0.00262f
C1782 a_7032_2153# VDPWR 0
C1783 uio_oe[0] uio_out[7] 0.03102f
C1784 a_6944_13645# a_4839_12857# 0
C1785 a_5851_13769# a_6329_12927# 0
C1786 a_14281_5467# VDPWR 0.00106f
C1787 sky130_fd_sc_hd__mux4_1_0.A2 a_12017_2159# 0
C1788 uo_out[1] uo_out[2] 0.03102f
C1789 a_11255_13773# a_11195_12931# 0.20048f
C1790 a_5851_13769# a_6021_13769# 0.00167f
C1791 a_5363_5043# a_6429_5043# 0.08312f
C1792 a_16454_4503# a_15188_4913# 0
C1793 VDPWR a_9451_16343# 0.02516f
C1794 a_6281_11907# a_6003_11935# 0.11706f
C1795 VDPWR a_8283_2049# 0.45076f
C1796 a_9381_11547# a_9771_12117# 0
C1797 a_9491_15377# a_9619_16343# 0
C1798 a_16402_4529# sky130_fd_sc_hd__mux4_1_0.A3 0
C1799 VDPWR a_17733_4529# 0.41856f
C1800 a_12769_4809# a_14825_4547# 0
C1801 a_9705_12861# a_4915_10549# 0
C1802 sky130_fd_sc_hd__mux4_1_0.A2 a_13969_1793# 0
C1803 a_4635_13809# a_5851_13769# 0
C1804 a_8377_5305# a_8263_5049# 0
C1805 a_12769_4809# sky130_fd_sc_hd__mux4_1_0.A3 0
C1806 a_6375_5299# a_8431_5415# 0
C1807 a_9629_14529# a_9705_12861# 0
C1808 a_10841_12931# a_11979_13399# 0
C1809 a_6071_2153# a_2187_1765# 0
C1810 sky130_fd_sc_hd__mux4_1_0.A2 a_7892_1793# 0.00121f
C1811 a_5269_1787# a_6698_2153# 0.03325f
C1812 a_17733_4529# a_17425_5473# 0.39935f
C1813 a_16847_4895# a_17210_4895# 0.00847f
C1814 a_10525_5837# a_10357_5837# 0
C1815 a_8431_5415# a_10132_5445# 0
C1816 a_11255_13773# a_9779_13785# 0
C1817 sky130_fd_sc_hd__mux4_1_0.A2 a_10289_1793# 0
C1818 VDPWR a_15188_4547# 0.22144f
C1819 ua[0] a_24962_14701# 0.13396f
C1820 uo_out[2] uo_out[3] 0.03102f
C1821 a_4505_13107# a_4905_12113# 0
C1822 a_4383_1787# a_2187_1765# 0
C1823 a_10841_12931# a_10717_13773# 0
C1824 a_6261_5043# sky130_fd_sc_hd__mux4_1_0.A3 0
C1825 a_4839_12857# a_4627_12141# 0
C1826 a_9619_16093# a_9703_16093# 0.00234f
C1827 a_2313_1791# a_2187_1765# 0.08436f
C1828 a_10799_13773# a_9703_16093# 0
C1829 a_24318_14385# a_23731_14309# 0.02707f
C1830 a_12533_5715# a_14152_5441# 0.00359f
C1831 a_13473_5459# a_12533_5715# 0.13739f
C1832 a_9379_14779# a_9769_15349# 0.00566f
C1833 VDPWR a_9589_10581# 0.00176f
C1834 a_10499_4853# a_12823_4553# 0
C1835 a_8431_5049# a_8038_5023# 0.02283f
C1836 VDPWR a_14377_5833# 0
C1837 a_12194_5433# a_12587_5459# 0.02283f
C1838 a_16297_2159# a_16129_2159# 0
C1839 a_10160_4571# a_10289_4963# 0.00792f
C1840 VDPWR a_15431_5467# 1.4342f
C1841 a_14281_5467# a_14545_5467# 0
C1842 a_4839_12857# a_4903_15345# 0.1369f
C1843 a_11175_1793# a_12113_1793# 0
C1844 VDPWR a_14545_5833# 0.00865f
C1845 a_7315_5043# sky130_fd_sc_hd__mux4_1_0.A3 0.00284f
C1846 a_16146_5447# a_16275_5473# 0.00758f
C1847 a_6335_1787# a_7944_1767# 0
C1848 VDPWR a_16994_1793# 0
C1849 VDPWR a_2145_1791# 0.00107f
C1850 a_4713_12141# a_4905_12113# 0
C1851 a_7831_14003# a_6389_13769# 0
C1852 a_8337_2159# a_8169_2159# 0
C1853 a_4755_12857# a_4839_12857# 0.00208f
C1854 a_2676_2157# a_2187_1765# 0.03547f
C1855 a_9631_11547# a_9493_12145# 0
C1856 a_16454_4503# a_16847_4895# 0.02301f
C1857 a_15431_5467# a_17425_5473# 0
C1858 sky130_fd_sc_hd__mux4_1_0.A1 a_9369_16343# 0
C1859 uio_out[3] uio_out[4] 0.03102f
C1860 a_6792_5043# a_6429_5043# 0.00985f
C1861 a_5851_13769# a_5933_13769# 0.00578f
C1862 VDPWR a_6127_13769# 0.0014f
C1863 a_9621_13111# a_9379_14779# 0
C1864 a_3938_1787# VDPWR 0.1394f
C1865 a_6629_15387# a_4903_15345# 0
C1866 a_14825_4547# a_13709_4553# 0.08312f
C1867 a_3010_2157# a_2187_1765# 0
C1868 a_6335_2153# VDPWR 0.00967f
C1869 a_10888_5471# a_10471_5727# 0.03016f
C1870 a_9493_12145# a_9503_10581# 0
C1871 a_2259_2047# a_2676_1791# 0.03016f
C1872 VDPWR a_11175_1793# 1.4104f
C1873 a_17544_4895# a_16793_4785# 0.00696f
C1874 a_13709_4553# sky130_fd_sc_hd__mux4_1_0.A3 0
C1875 a_2217_5025# a_1950_5025# 0.08244f
C1876 a_10160_4571# a_10471_5727# 0
C1877 sky130_fd_sc_hd__mux4_1_0.A2 a_12644_1793# 0
C1878 VDPWR a_7944_1767# 0.35009f
C1879 a_10261_5837# a_10132_5445# 0.00792f
C1880 a_2187_1765# a_4215_2153# 0
C1881 a_16297_1793# a_16129_1793# 0
C1882 VDPWR a_23731_14309# 0.46521f
C1883 a_12194_5433# sky130_fd_sc_hd__mux4_1_0.A3 0.0051f
C1884 a_9317_5049# a_12533_5715# 0
C1885 VDPWR a_4213_5043# 0.00118f
C1886 a_16243_2049# a_16297_2159# 0.03622f
C1887 VDPWR a_24318_14385# 0.00521f
C1888 a_10471_5727# a_12950_5459# 0
C1889 a_14432_4521# a_14825_4547# 0.02283f
C1890 a_6087_14735# a_6862_13645# 0
C1891 a_2259_2047# a_3010_1791# 0.00682f
C1892 VDPWR a_10385_4963# 0
C1893 a_4477_5043# a_4309_5043# 0
C1894 a_14281_5467# a_14152_5441# 0.00758f
C1895 VDPWR a_12323_5825# 0
C1896 a_14281_5467# a_13473_5459# 0
C1897 a_14432_4521# sky130_fd_sc_hd__mux4_1_0.A3 0
C1898 a_4215_1787# VDPWR 0
C1899 a_12615_14007# sky130_fd_sc_hd__mux4_1_0.A1 0.10822f
C1900 a_11250_4963# a_10499_4853# 0.00696f
C1901 a_16094_5473# sky130_fd_sc_hd__mux4_1_0.A3 0.0031f
C1902 a_4585_16339# VDPWR 0.02516f
C1903 VDPWR a_6335_1787# 0.18613f
C1904 a_5975_12927# a_5809_14763# 0
C1905 a_7126_5043# a_6375_5299# 0.00682f
C1906 VDPWR a_12113_1793# 0
C1907 a_16539_5839# a_16371_5839# 0
C1908 a_6261_5409# VDPWR 0
C1909 a_14596_2159# a_14179_2049# 0.06611f
C1910 sky130_fd_sc_hd__mux4_1_0.A2 a_14825_4547# 0
C1911 a_2343_5051# a_2706_5051# 0.00985f
C1912 a_12769_4809# a_12587_5825# 0
C1913 VDPWR a_4032_5043# 0.13943f
C1914 a_11147_11911# a_12697_14007# 0.00377f
C1915 VDPWR a_10525_5471# 0.18051f
C1916 a_10025_2159# a_9896_1767# 0.00792f
C1917 VDPWR a_4711_15373# 0.00333f
C1918 sky130_fd_sc_hd__mux4_1_0.A2 sky130_fd_sc_hd__mux4_1_0.A3 0.91673f
C1919 uio_oe[0] uio_oe[1] 0.03102f
C1920 a_9769_15349# a_9369_16343# 0
C1921 VDPWR a_19510_16177# 0.46458f
C1922 a_2175_5051# a_1950_5025# 0.00487f
C1923 a_16539_5839# a_14491_5723# 0
C1924 a_16033_1793# a_16297_1793# 0
C1925 a_10235_2049# a_11175_1793# 0.13739f
C1926 a_16539_5473# a_16275_5473# 0
C1927 a_13969_2159# sky130_fd_sc_hd__mux4_1_0.A2 0
C1928 VDPWR a_10108_4597# 0.12354f
C1929 sky130_fd_sc_hd__mux4_1_0.A2 a_12644_2159# 0
C1930 a_10953_14739# a_9379_14779# 0
C1931 sky130_fd_sc_hd__mux4_1_0.A2 a_10499_4853# 0
C1932 a_7126_5409# sky130_fd_sc_hd__mux4_1_0.A3 0
C1933 a_14377_5833# a_14152_5441# 0.00559f
C1934 a_7173_15235# a_4915_10549# 0.09278f
C1935 a_15188_4913# a_14491_5723# 0
C1936 VDPWR a_17425_5473# 0.2756f
C1937 a_12227_2049# a_11888_1767# 0.04737f
C1938 a_14545_5833# a_14152_5441# 0.02301f
C1939 sky130_fd_sc_hd__mux4_1_0.A2 a_12378_4553# 0
C1940 sky130_fd_sc_hd__mux4_1_0.A2 a_16297_1793# 0
C1941 a_6261_5043# a_6036_5017# 0.00487f
C1942 a_2187_1765# a_1920_1765# 0.08244f
C1943 a_4839_12857# a_4513_14775# 0.00442f
C1944 a_4847_14525# a_5851_13769# 0
C1945 a_9034_2159# a_8283_2049# 0.00696f
C1946 a_9317_5049# a_17733_4529# 0.37402f
C1947 a_14419_5441# a_14380_4547# 0
C1948 a_9713_14529# a_10717_13773# 0
C1949 a_9379_14779# a_9703_16093# 0
C1950 uio_in[1] uio_in[2] 0.03102f
C1951 a_11222_5471# a_10471_5727# 0.00682f
C1952 a_4119_1787# a_3990_1761# 0.00758f
C1953 a_8377_5305# a_10080_5471# 0
C1954 a_4746_2153# a_4383_2153# 0.00847f
C1955 a_10471_5727# a_10132_5445# 0.04737f
C1956 a_5363_5043# sky130_fd_sc_hd__mux4_1_0.A3 0.00183f
C1957 a_4515_11543# a_4905_12113# 0
C1958 a_9501_13813# a_9629_14779# 0
C1959 a_9896_1767# a_8283_2049# 0.00419f
C1960 a_10525_5837# a_10261_5837# 0
C1961 a_16902_5839# a_14491_5723# 0
C1962 sky130_fd_sc_hd__mux4_1_0.A2 a_6281_2043# 0.00307f
C1963 a_8794_5049# a_7315_5043# 0.08907f
C1964 sky130_fd_sc_hd__mux4_1_0.A2 a_16679_4529# 0
C1965 VDPWR a_14545_5467# 0.18449f
C1966 a_12194_5433# a_12587_5825# 0.02301f
C1967 VDPWR a_2706_5417# 0.021f
C1968 a_16793_4785# a_18625_4938# 0
C1969 a_23677_14701# a_23731_14309# 0.09132f
C1970 a_10235_2049# VDPWR 0.45058f
C1971 a_24241_14651# a_23731_14309# 0.02645f
C1972 a_12281_2159# a_12017_2159# 0
C1973 a_4505_13107# a_4839_12857# 0.16952f
C1974 a_12615_14007# a_12039_15239# 0.16707f
C1975 a_24241_14651# a_24318_14385# 0.01352f
C1976 a_5080_1787# a_4329_2043# 0.00682f
C1977 a_11175_1793# a_12017_1793# 0
C1978 a_15431_5467# a_9317_5049# 0.0454f
C1979 a_6944_13645# a_6389_13769# 0.00183f
C1980 a_7831_14003# a_6281_11907# 0.00377f
C1981 a_9223_1793# a_10652_2159# 0.03325f
C1982 a_9379_14779# a_4915_10549# 0
C1983 a_13840_1767# a_14233_1793# 0.02283f
C1984 a_4383_2153# a_4329_2043# 0.03622f
C1985 a_9629_14529# a_9379_14779# 0.00723f
C1986 a_10652_1793# a_11175_1793# 0
C1987 a_10385_4963# a_10553_4963# 0
C1988 a_21506_16181# a_20384_16179# 0.10183f
C1989 a_4635_13809# a_4847_14525# 0
C1990 a_6635_15235# a_6862_13645# 0
C1991 a_9503_10581# a_9781_10553# 0.1296f
C1992 a_11411_5471# a_12419_5459# 0
C1993 VDPWR a_9491_15377# 0.45072f
C1994 a_11147_11911# a_9771_12117# 0.03573f
C1995 a_6629_15387# a_8193_13753# 0.05689f
C1996 a_10080_5471# a_10132_5445# 0.1439f
C1997 a_9587_13813# a_4915_10549# 0
C1998 a_15852_1793# a_15119_1793# 0.05087f
C1999 VDPWR a_9577_15377# 0.00333f
C2000 a_6717_15235# a_4847_14525# 0.00159f
C2001 a_14233_1793# a_13167_1793# 0.08312f
C2002 VDPWR a_23677_14701# 0.21646f
C2003 VDPWR a_14152_5441# 0.34016f
C2004 VDPWR a_13473_5459# 0.12977f
C2005 a_6792_5043# sky130_fd_sc_hd__mux4_1_0.A3 0
C2006 a_16146_5447# a_15431_5467# 0.11891f
C2007 a_10869_11939# a_9493_12145# 0
C2008 a_9631_11547# a_4915_10549# 0
C2009 a_14771_4803# a_14825_4913# 0.03622f
C2010 a_11979_13399# a_11728_13649# 0.10945f
C2011 a_24241_14651# VDPWR 0.27727f
C2012 a_7315_5043# a_8377_5305# 0.21187f
C2013 a_17254_16187# a_19510_16177# 0
C2014 a_16485_5729# sky130_fd_sc_hd__mux4_1_0.A3 0.00779f
C2015 VDPWR a_14065_1793# 0
C2016 a_9713_14529# a_8193_13753# 0.29837f
C2017 a_16793_4785# sky130_fd_sc_hd__mux4_1_0.A3 0
C2018 VDPWR a_17254_16187# 0.4937f
C2019 a_9703_16093# a_9369_16343# 0.16891f
C2020 VDPWR a_10553_4963# 0.05574f
C2021 a_9503_10581# a_4915_10549# 0.001f
C2022 a_10717_13773# a_11728_13649# 0
C2023 a_4903_15345# a_6389_13769# 0
C2024 VDPWR a_12017_1793# 0.00118f
C2025 VDPWR a_4309_5043# 0
C2026 a_8169_1793# a_7221_1787# 0
C2027 ui_in[0] sky130_fd_sc_hd__mux4_1_0.A1 0.00242f
C2028 a_8700_1793# a_8337_1793# 0.00985f
C2029 a_16539_5839# a_16275_5839# 0
C2030 a_5895_14763# a_4839_12857# 0
C2031 a_9493_12145# a_9371_13111# 0.00144f
C2032 a_4903_15345# a_4837_16089# 0.50558f
C2033 sky130_fd_sc_hd__mux4_1_0.A2 a_14596_2159# 0
C2034 a_4913_13781# a_6862_13645# 0
C2035 a_10525_5837# a_10471_5727# 0.03622f
C2036 a_7892_1793# a_8073_2159# 0
C2037 VDPWR a_14596_1793# 0.21795f
C2038 a_10675_14767# a_10717_13773# 0
C2039 a_10841_12931# a_9769_15349# 0
C2040 a_23511_14701# a_23731_14309# 0.00549f
C2041 sky130_fd_sc_hd__mux4_1_0.A2 a_6698_2153# 0
C2042 a_11147_11911# a_11979_13399# 0.19568f
C2043 VDPWR a_10652_1793# 0.21796f
C2044 sky130_fd_sc_hd__mux4_1_0.A2 a_8700_1793# 0
C2045 a_12793_14007# a_9781_10553# 0
C2046 a_6261_5043# a_6375_5299# 0
C2047 a_12978_1793# sky130_fd_sc_hd__mux4_1_0.A2 0
C2048 VDPWR a_14065_2159# 0
C2049 ui_in[1] ui_in[0] 5.58248f
C2050 VDPWR a_9317_5049# 2.60485f
C2051 a_17544_4529# VDPWR 0
C2052 VDPWR a_6129_12927# 0
C2053 a_13840_1767# a_12227_2049# 0.00419f
C2054 a_9493_12145# a_9381_11547# 0
C2055 VDPWR a_9034_2159# 0
C2056 a_12430_4527# a_12559_4919# 0.00792f
C2057 a_14545_5467# a_14152_5441# 0.02283f
C2058 a_14545_5467# a_13473_5459# 0
C2059 sky130_fd_sc_hd__mux4_1_0.A2 a_10160_4571# 0
C2060 a_11147_11911# a_10717_13773# 0
C2061 VDPWR a_10916_4597# 0.31242f
C2062 a_7315_5043# a_6375_5299# 0.13739f
C2063 a_12430_4527# a_11439_4597# 0.1189f
C2064 a_14908_5833# a_12533_5715# 0
C2065 ua[4] a_14179_2049# 0
C2066 a_7113_13395# a_4915_10549# 0.20109f
C2067 a_11147_11911# a_12865_14007# 0
C2068 a_15711_4547# a_17733_4529# 0.00125f
C2069 a_5363_5043# a_6036_5017# 0.11878f
C2070 sky130_fd_sc_hd__mux4_1_0.A2 a_10121_1793# 0
C2071 a_12615_14007# a_9781_10553# 0.07615f
C2072 a_7173_15235# a_7749_14003# 0.16707f
C2073 a_10553_4597# VDPWR 0.27571f
C2074 a_9317_5049# a_17425_5473# 0.24941f
C2075 a_8700_2159# a_7221_1787# 0.03325f
C2076 a_5269_1787# a_7221_1787# 0
C2077 a_11175_1793# a_11888_1767# 0.11874f
C2078 a_6629_15387# a_4625_15373# 0
C2079 a_16402_4529# a_16583_4895# 0
C2080 a_14771_4803# a_15188_4913# 0.06611f
C2081 a_8337_2159# a_8700_2159# 0.00847f
C2082 a_9621_13111# a_9371_13111# 0.02504f
C2083 a_7999_14003# a_7173_15235# 0
C2084 a_2343_5051# a_1950_5025# 0.02283f
C2085 a_2259_2047# a_2187_1765# 0.25757f
C2086 VDPWR a_7032_1787# 0
C2087 a_13788_1793# a_13840_1767# 0.1439f
C2088 VDPWR a_9896_1767# 0.35015f
C2089 a_13167_1793# a_12227_2049# 0.13739f
C2090 a_3938_1787# a_3990_1761# 0.1439f
C2091 a_12419_5459# a_12587_5459# 0
C2092 a_5269_1787# a_3199_1791# 0
C2093 VDPWR a_6087_14735# 0.4457f
C2094 VDPWR a_12823_4919# 0.01321f
C2095 a_15119_1793# a_14179_2049# 0.13739f
C2096 a_15188_4547# a_15711_4547# 0
C2097 ua[6] a_7221_1787# 0
C2098 a_4477_5409# a_3229_5051# 0.04534f
C2099 a_16793_4785# a_16679_4529# 0
C2100 a_4839_12857# a_5809_14763# 0.21957f
C2101 a_6629_15387# sky130_fd_sc_hd__mux4_1_0.A1 0.10747f
C2102 a_12430_4527# a_11411_5471# 0
C2103 a_9491_15377# a_9577_15377# 0.00658f
C2104 a_16146_5447# VDPWR 0.35424f
C2105 a_15431_5467# a_16539_5473# 0.08313f
C2106 a_8431_5049# a_8263_5049# 0
C2107 VDPWR a_23511_14701# 0.19914f
C2108 a_17236_5839# sky130_fd_sc_hd__mux4_1_0.A3 0
C2109 a_1868_1791# a_2049_2157# 0
C2110 a_4847_14525# a_6805_15235# 0.00624f
C2111 sky130_fd_sc_hd__mux4_1_0.A2 a_12113_2159# 0
C2112 a_13788_1793# a_13167_1793# 0.05218f
C2113 a_3040_5417# a_3229_5051# 0
C2114 a_12281_2159# a_12644_2159# 0.00847f
C2115 a_8167_5415# a_7986_5049# 0
C2116 a_6629_15387# a_5809_14763# 0
C2117 a_15711_4547# a_15431_5467# 0
C2118 a_10235_2049# a_10652_1793# 0.03016f
C2119 VDPWR a_5080_2153# 0
C2120 a_13473_5459# a_14152_5441# 0
C2121 a_11888_1767# a_12113_1793# 0.00487f
C2122 VDPWR a_9705_12861# 1.15673f
C2123 a_4839_12857# a_4515_11543# 0
C2124 a_5174_5409# a_2217_5025# 0
C2125 a_23511_14335# sky130_fd_sc_hd__mux4_1_0.A3 0.00544f
C2126 a_4215_1787# a_3990_1761# 0.00487f
C2127 a_12769_4809# a_13520_4919# 0.00696f
C2128 a_14419_5441# a_14100_5467# 0.0459f
C2129 a_14771_4803# a_14657_4913# 0
C2130 a_6944_13645# a_6281_11907# 0
C2131 VDPWR a_2313_2157# 0.00827f
C2132 a_9463_11547# a_9381_11547# 0.00641f
C2133 a_14930_1793# VDPWR 0
C2134 a_12533_5715# a_13284_5825# 0.00696f
C2135 a_12419_5459# sky130_fd_sc_hd__mux4_1_0.A3 0
C2136 a_10675_14767# a_8193_13753# 0
C2137 a_18742_16187# a_20384_16179# 0
C2138 a_5363_5043# a_6165_5043# 0
C2139 a_6089_11935# a_4905_12113# 0
C2140 a_4746_2153# a_3199_1791# 0.03325f
C2141 a_6057_12927# a_5975_12927# 0.00517f
C2142 a_15904_1767# VDPWR 0.34973f
C2143 ui_in[0] ua[0] 0.38436f
C2144 a_6792_5409# sky130_fd_sc_hd__mux4_1_0.A3 0
C2145 VDPWR a_11888_1767# 0.35008f
C2146 a_4915_10549# a_4905_12113# 0.0298f
C2147 a_14380_4547# sky130_fd_sc_hd__mux4_1_0.A3 0
C2148 a_4847_14525# a_4763_14525# 0.00206f
C2149 a_10235_2049# a_9896_1767# 0.04737f
C2150 a_4513_14775# a_4837_16089# 0
C2151 a_9461_14779# a_9769_15349# 0
C2152 a_16146_5447# a_14545_5467# 0
C2153 VDPWR a_2079_5417# 0
C2154 a_2175_5417# a_1950_5025# 0.00559f
C2155 a_6281_11907# a_7927_14003# 0.00264f
C2156 a_6629_15387# a_4503_16339# 0
C2157 a_2289_5307# a_2343_5417# 0.03622f
C2158 VDPWR a_3990_1761# 0.35029f
C2159 a_11671_15239# a_12039_15239# 0
C2160 a_10869_11939# a_9703_16093# 0
C2161 a_4477_5409# a_4309_5409# 0
C2162 a_17210_4895# a_17733_4529# 0
C2163 a_13969_2159# a_14233_2159# 0
C2164 a_10869_11939# a_9781_10553# 0
C2165 VDPWR a_11250_4597# 0
C2166 a_9317_5049# a_14152_5441# 0
C2167 a_24234_14385# ui_in[1] 0.34724f
C2168 a_13473_5459# a_9317_5049# 0.00435f
C2169 a_7126_5409# a_6375_5299# 0.00696f
C2170 ua[5] a_11175_1793# 0
C2171 a_4627_12141# a_6281_11907# 0
C2172 a_15119_1793# a_16129_1793# 0
C2173 a_16243_2049# a_16994_1793# 0.00682f
C2174 a_14419_5441# a_11411_5471# 0
C2175 a_10841_12931# a_9703_16093# 0
C2176 a_13520_4919# a_13709_4553# 0
C2177 a_3199_1791# a_4329_2043# 0.21188f
C2178 a_1898_5051# a_2217_5025# 0.0073f
C2179 a_7113_13395# a_6862_13645# 0.10945f
C2180 a_9713_14529# a_9769_15349# 0.15227f
C2181 VDPWR a_9619_16093# 0.00495f
C2182 VDPWR a_11810_13649# 0.0014f
C2183 a_24318_14385# a_24407_14651# 0
C2184 VDPWR a_10799_13773# 0
C2185 a_14908_5833# a_14545_5833# 0.00847f
C2186 sky130_fd_sc_hd__mux4_1_0.A2 a_10986_1793# 0
C2187 a_9619_16343# a_9369_16343# 0.02504f
C2188 VDPWR a_15242_5467# 0
C2189 a_4763_14775# a_4839_12857# 0.00187f
C2190 VDPWR a_10923_12931# 0
C2191 VDPWR a_16539_5473# 0.18678f
C2192 a_16454_4503# a_17733_4529# 0
C2193 a_2313_1791# a_1920_1765# 0.02283f
C2194 a_8167_5415# sky130_fd_sc_hd__mux4_1_0.A3 0
C2195 a_4913_13781# a_6127_13769# 0
C2196 a_10955_11939# a_9781_10553# 0
C2197 a_2343_5051# a_2079_5051# 0
C2198 a_5363_5043# a_6375_5299# 0.21187f
C2199 a_14432_4521# a_14561_4913# 0.00792f
C2200 a_9223_1793# a_10025_1793# 0
C2201 a_14825_4913# a_13709_4553# 0.04534f
C2202 VDPWR a_2706_5051# 0.21783f
C2203 VDPWR a_15711_4547# 1.4869f
C2204 a_5975_12927# a_6862_13645# 0
C2205 a_10235_2049# a_11888_1767# 0.00395f
C2206 sky130_fd_sc_hd__mux4_1_0.A2 a_10385_4597# 0
C2207 VDPWR a_4755_13107# 0.33272f
C2208 a_4477_5409# a_2217_5025# 0
C2209 a_23511_14701# a_23677_14701# 0.05551f
C2210 VDPWR a_16129_2159# 0
C2211 a_12419_5825# a_12533_5715# 0
C2212 a_9713_14529# a_12039_15239# 0
C2213 a_15711_4547# a_17425_5473# 0
C2214 a_8169_2159# a_8283_2049# 0
C2215 a_5269_1787# a_5942_1761# 0.11878f
C2216 a_4847_14525# a_4595_14775# 0
C2217 a_9781_10553# a_9381_11547# 0
C2218 a_24962_14701# a_23731_14309# 0
C2219 a_11411_5471# a_11439_4597# 0
C2220 a_12194_5433# a_10525_5837# 0
C2221 a_14432_4521# a_14825_4913# 0.02301f
C2222 a_16033_1793# a_15119_1793# 0
C2223 a_16847_4529# a_16679_4529# 0
C2224 sky130_fd_sc_hd__mux4_1_0.A2 a_10121_2159# 0
C2225 VDPWR a_6635_15235# 0.42119f
C2226 a_10471_5727# a_11222_5837# 0.00696f
C2227 a_10953_14739# a_11671_15239# 0.00366f
C2228 a_9371_13111# a_4915_10549# 0.00232f
C2229 uio_in[5] uio_in[4] 0.03102f
C2230 VDPWR a_9128_5415# 0
C2231 a_3040_5417# a_2217_5025# 0
C2232 a_10289_2159# sky130_fd_sc_hd__mux4_1_0.A2 0
C2233 a_11501_15239# a_11671_15239# 0.00167f
C2234 a_5942_1761# a_5890_1787# 0.1439f
C2235 a_7113_13395# a_7749_14003# 0.27996f
C2236 VDPWR a_24407_14651# 0.00293f
C2237 a_12430_4527# sky130_fd_sc_hd__mux4_1_0.A3 0
C2238 a_2049_1791# a_2313_1791# 0
C2239 a_11255_13773# a_12697_14007# 0
C2240 ua[5] VDPWR 0.00172f
C2241 a_16454_4503# a_15431_5467# 0
C2242 a_10553_4597# a_10916_4597# 0.00985f
C2243 a_2676_1791# a_3199_1791# 0
C2244 a_7999_14003# a_7113_13395# 0.00205f
C2245 a_18371_4938# sky130_fd_sc_hd__mux4_1_0.A3 0.00367f
C2246 a_11147_11911# sky130_fd_sc_hd__mux4_1_0.A1 0.00289f
C2247 a_24152_14385# ui_in[0] 0.03464f
C2248 a_12430_4527# a_10499_4853# 0.00138f
C2249 a_24234_14385# ua[0] 0
C2250 a_13167_1793# a_11175_1793# 0
C2251 sky130_fd_sc_hd__mux4_1_0.A2 a_15119_1793# 0.00765f
C2252 a_9381_11547# a_4915_10549# 0.00227f
C2253 a_11671_15239# a_9703_16093# 0
C2254 VDPWR a_7173_15235# 0.7127f
C2255 a_16243_2049# VDPWR 0.43625f
C2256 a_4903_15345# a_5851_13769# 0.16757f
C2257 a_5363_5043# a_3229_5051# 0
C2258 a_16146_5447# a_9317_5049# 0
C2259 a_4746_1787# a_3199_1791# 0.08907f
C2260 uo_out[1] uo_out[0] 0.03102f
C2261 a_8431_5049# a_8167_5049# 0
C2262 a_10888_5837# sky130_fd_sc_hd__mux4_1_0.A3 0.00192f
C2263 a_5895_14763# a_4837_16089# 0
C2264 a_12430_4527# a_12378_4553# 0.1439f
C2265 a_15188_4913# a_13709_4553# 0.03325f
C2266 VDPWR a_8038_5023# 0.35038f
C2267 a_6792_5043# a_6375_5299# 0.03016f
C2268 a_21506_16181# a_22274_16171# 0.1036f
C2269 VDPWR a_4913_13781# 0.76099f
C2270 VDPWR a_24962_14701# 0.29288f
C2271 a_9589_10581# a_9503_10581# 0.00658f
C2272 a_9779_13785# a_10887_13773# 0.00104f
C2273 a_9451_16343# a_9369_16343# 0.00641f
C2274 a_12017_1793# a_11888_1767# 0.00758f
C2275 VDPWR a_14908_5833# 0.02196f
C2276 a_9769_15349# a_11728_13649# 0
C2277 a_5080_1787# a_2187_1765# 0
C2278 a_9453_13111# a_4915_10549# 0
C2279 a_9779_13785# a_9771_12117# 0.00627f
C2280 a_16297_1793# a_16660_1793# 0.00985f
C2281 a_10953_14739# a_9713_14529# 0.31937f
C2282 a_4625_15373# a_4837_16089# 0
C2283 a_4423_5299# a_5174_5409# 0.00696f
C2284 a_4383_2153# a_2187_1765# 0
C2285 VDPWR a_17210_4895# 0.02205f
C2286 a_11836_1793# a_11175_1793# 0.05174f
C2287 a_12950_5825# a_12533_5715# 0.06611f
C2288 a_13840_1767# VDPWR 0.35015f
C2289 a_4637_10577# a_4765_11543# 0
C2290 a_11501_15239# a_9713_14529# 0.17821f
C2291 VDPWR a_8263_5415# 0
C2292 a_10675_14767# a_9769_15349# 0.00346f
C2293 a_10235_2049# ua[5] 0
C2294 a_11147_11911# a_9493_12145# 0
C2295 a_8169_2159# a_7944_1767# 0.00559f
C2296 a_9501_13813# a_10717_13773# 0
C2297 VDPWR a_13520_4553# 0
C2298 a_11195_12931# a_11979_13399# 0
C2299 a_4635_13809# a_4627_12141# 0
C2300 a_14596_2159# a_14233_2159# 0.00847f
C2301 a_4903_15345# a_6021_13769# 0.00818f
C2302 a_14419_5441# sky130_fd_sc_hd__mux4_1_0.A3 0.00398f
C2303 a_5942_1761# a_4329_2043# 0.00419f
C2304 sky130_fd_sc_hd__mux4_1_0.A2 ui_in[1] 0.24408f
C2305 a_4119_2153# a_4383_2153# 0
C2306 a_9713_14529# a_9703_16093# 0.46419f
C2307 a_12281_2159# a_12113_2159# 0
C2308 a_12587_5459# a_11439_4597# 0
C2309 a_4903_15345# a_4635_13809# 0.00159f
C2310 a_4839_12857# a_4587_13107# 0
C2311 VDPWR a_13167_1793# 1.41083f
C2312 a_11195_12931# a_10717_13773# 0
C2313 VDPWR a_9379_14779# 0.51116f
C2314 a_4839_12857# a_4915_10549# 0.00242f
C2315 a_12281_1793# a_12644_1793# 0.00985f
C2316 a_12323_5459# VDPWR 0.0012f
C2317 a_20384_16179# sky130_fd_sc_hd__mux4_1_0.A1 0
C2318 a_4477_5409# a_4213_5409# 0
C2319 a_5809_14763# a_4837_16089# 0.03093f
C2320 a_16454_4503# VDPWR 0.37148f
C2321 a_10675_14767# a_12039_15239# 0
C2322 a_8337_1793# a_7221_1787# 0.08313f
C2323 a_9631_11297# a_4915_10549# 0
C2324 a_4627_12141# a_4637_10577# 0
C2325 a_17544_4895# sky130_fd_sc_hd__mux4_1_0.A3 0
C2326 a_6698_1787# a_6281_2043# 0.03016f
C2327 a_14432_4521# a_14657_4913# 0.00559f
C2328 a_14100_5467# sky130_fd_sc_hd__mux4_1_0.A3 0.00306f
C2329 a_5269_1787# a_6167_1787# 0
C2330 a_13284_5459# sky130_fd_sc_hd__mux4_1_0.A3 0
C2331 a_11255_13773# a_10887_13773# 0
C2332 VDPWR a_4721_13809# 0.003f
C2333 sky130_fd_sc_hd__mux4_1_0.A2 a_7221_1787# 0.00286f
C2334 a_24241_14651# a_24407_14651# 0.00988f
C2335 a_6429_5043# sky130_fd_sc_hd__mux4_1_0.A3 0
C2336 a_11411_5471# a_12587_5459# 0.08312f
C2337 a_7315_5043# a_8431_5049# 0.08313f
C2338 a_4503_16339# a_4753_16089# 0.00723f
C2339 VDPWR a_9587_13813# 0.003f
C2340 a_9779_13785# a_10717_13773# 0.00386f
C2341 sky130_fd_sc_hd__mux4_1_0.A2 a_8337_2159# 0
C2342 a_10160_4571# a_10289_4597# 0.00758f
C2343 a_11147_11911# a_12039_15239# 0.09952f
C2344 a_2259_2047# a_2313_1791# 0.00386f
C2345 a_12559_4919# sky130_fd_sc_hd__mux4_1_0.A3 0
C2346 VDPWR a_14377_5467# 0
C2347 VDPWR a_11836_1793# 0.13944f
C2348 VDPWR a_8169_2159# 0
C2349 a_9713_14529# a_4915_10549# 0
C2350 a_6281_11907# a_8193_13753# 0.00288f
C2351 VDPWR a_9631_11547# 0.33144f
C2352 a_11439_4597# sky130_fd_sc_hd__mux4_1_0.A3 0
C2353 a_15188_4547# a_14491_5723# 0
C2354 a_2049_1791# a_1920_1765# 0.00758f
C2355 a_24234_14385# a_24152_14385# 0.04662f
C2356 a_15711_4547# a_9317_5049# 0.03084f
C2357 a_4627_12141# a_6003_11935# 0
C2358 a_4503_16339# a_4837_16089# 0.16891f
C2359 a_16371_5473# a_16485_5729# 0
C2360 a_9629_14529# a_9713_14529# 0.00206f
C2361 ui_in[6] ui_in[7] 0.03102f
C2362 a_4903_15345# a_5933_13769# 0.0035f
C2363 VDPWR a_9503_10581# 0.43168f
C2364 a_4839_12857# a_6057_12927# 0.00148f
C2365 a_5363_5043# a_2217_5025# 0.0013f
C2366 a_16679_4895# a_16793_4785# 0
C2367 a_10499_4853# a_12559_4919# 0
C2368 a_4423_5299# a_4477_5409# 0.03622f
C2369 ua[1] VGND 0.14696f
C2370 ua[2] VGND 0.14696f
C2371 ua[3] VGND 0.14696f
C2372 ua[4] VGND 0.14481f
C2373 ua[5] VGND 0.14481f
C2374 ua[6] VGND 0.1449f
C2375 ua[7] VGND 0.14552f
C2376 ena VGND 0.07038f
C2377 clk VGND 0.04288f
C2378 rst_n VGND 0.04288f
C2379 ui_in[2] VGND 0.04288f
C2380 ui_in[3] VGND 0.04288f
C2381 ui_in[4] VGND 0.04288f
C2382 ui_in[5] VGND 0.04288f
C2383 ui_in[6] VGND 0.04288f
C2384 ui_in[7] VGND 0.04288f
C2385 uio_in[0] VGND 0.04288f
C2386 uio_in[1] VGND 0.04288f
C2387 uio_in[2] VGND 0.04288f
C2388 uio_in[3] VGND 0.04288f
C2389 uio_in[4] VGND 0.04288f
C2390 uio_in[5] VGND 0.04288f
C2391 uio_in[6] VGND 0.04288f
C2392 uio_in[7] VGND 0.04288f
C2393 uo_out[0] VGND 0.04288f
C2394 uo_out[1] VGND 0.04288f
C2395 uo_out[2] VGND 0.04288f
C2396 uo_out[3] VGND 0.04288f
C2397 uo_out[4] VGND 0.04288f
C2398 uo_out[5] VGND 0.04288f
C2399 uo_out[6] VGND 0.04288f
C2400 uo_out[7] VGND 0.04288f
C2401 uio_out[0] VGND 0.04288f
C2402 uio_out[1] VGND 0.04288f
C2403 uio_out[2] VGND 0.04288f
C2404 uio_out[3] VGND 0.04288f
C2405 uio_out[4] VGND 0.04288f
C2406 uio_out[5] VGND 0.04288f
C2407 uio_out[6] VGND 0.04288f
C2408 uio_out[7] VGND 0.04288f
C2409 uio_oe[0] VGND 0.04288f
C2410 uio_oe[1] VGND 0.04288f
C2411 uio_oe[2] VGND 0.04288f
C2412 uio_oe[3] VGND 0.04288f
C2413 uio_oe[4] VGND 0.04288f
C2414 uio_oe[5] VGND 0.04288f
C2415 uio_oe[6] VGND 0.04288f
C2416 uio_oe[7] VGND 0.07038f
C2417 ua[0] VGND 9.56443f
C2418 ui_in[1] VGND 9.1369f
C2419 ui_in[0] VGND 9.30843f
C2420 VDPWR VGND 0.22134p
C2421 a_16994_1793# VGND 0
C2422 a_16660_1793# VGND 0.01465f
C2423 a_16297_1793# VGND 0.02017f
C2424 a_16129_1793# VGND 0
C2425 a_16033_1793# VGND 0
C2426 a_14930_1793# VGND 0
C2427 a_14596_1793# VGND 0.01679f
C2428 a_14233_1793# VGND 0.02017f
C2429 a_14065_1793# VGND 0
C2430 a_13969_1793# VGND 0
C2431 a_16994_2159# VGND 0.00217f
C2432 a_16660_2159# VGND 0.1985f
C2433 a_16297_2159# VGND 0.21682f
C2434 a_16129_2159# VGND 0.00234f
C2435 a_16033_2159# VGND 0.00307f
C2436 a_15852_1793# VGND 0.15057f
C2437 a_12978_1793# VGND 0
C2438 a_12644_1793# VGND 0.01679f
C2439 a_12281_1793# VGND 0.02014f
C2440 a_12113_1793# VGND 0
C2441 a_12017_1793# VGND 0
C2442 a_14930_2159# VGND 0.00244f
C2443 a_14596_2159# VGND 0.20226f
C2444 a_14233_2159# VGND 0.21682f
C2445 a_14065_2159# VGND 0.00233f
C2446 a_13969_2159# VGND 0.00307f
C2447 a_13788_1793# VGND 0.14753f
C2448 a_10986_1793# VGND 0
C2449 a_10652_1793# VGND 0.01679f
C2450 a_10289_1793# VGND 0.02017f
C2451 a_10121_1793# VGND 0
C2452 a_10025_1793# VGND 0
C2453 a_12978_2159# VGND 0.00242f
C2454 a_12644_2159# VGND 0.20221f
C2455 a_12281_2159# VGND 0.21675f
C2456 a_12113_2159# VGND 0.00232f
C2457 a_12017_2159# VGND 0.00306f
C2458 a_11836_1793# VGND 0.14801f
C2459 a_9034_1793# VGND 0
C2460 a_8700_1793# VGND 0.01679f
C2461 a_8337_1793# VGND 0.02015f
C2462 a_8169_1793# VGND 0
C2463 a_8073_1793# VGND 0
C2464 a_10986_2159# VGND 0.00244f
C2465 a_10652_2159# VGND 0.20227f
C2466 a_10289_2159# VGND 0.21687f
C2467 a_10121_2159# VGND 0.00233f
C2468 a_10025_2159# VGND 0.00307f
C2469 a_9844_1793# VGND 0.14753f
C2470 a_7032_1787# VGND 0
C2471 a_6698_1787# VGND 0.01676f
C2472 a_6335_1787# VGND 0.02015f
C2473 a_6167_1787# VGND 0
C2474 a_6071_1787# VGND 0
C2475 a_9034_2159# VGND 0.00242f
C2476 a_8700_2159# VGND 0.20221f
C2477 a_8337_2159# VGND 0.21675f
C2478 a_8169_2159# VGND 0.00232f
C2479 a_8073_2159# VGND 0.00307f
C2480 a_7892_1793# VGND 0.14822f
C2481 a_5080_1787# VGND 0
C2482 a_4746_1787# VGND 0.01677f
C2483 a_4383_1787# VGND 0.02013f
C2484 a_4215_1787# VGND 0
C2485 a_4119_1787# VGND 0
C2486 a_7032_2153# VGND 0.00244f
C2487 a_6698_2153# VGND 0.20225f
C2488 a_6335_2153# VGND 0.21685f
C2489 a_6167_2153# VGND 0.00233f
C2490 a_6071_2153# VGND 0.00307f
C2491 a_5890_1787# VGND 0.14746f
C2492 a_3010_1791# VGND 0
C2493 a_2676_1791# VGND 0.01809f
C2494 a_2313_1791# VGND 0.01957f
C2495 a_2145_1791# VGND 0
C2496 a_2049_1791# VGND 0
C2497 a_5080_2153# VGND 0.00242f
C2498 a_4746_2153# VGND 0.20219f
C2499 a_4383_2153# VGND 0.21674f
C2500 a_4215_2153# VGND 0.00231f
C2501 a_4119_2153# VGND 0.00305f
C2502 a_3938_1787# VGND 0.14876f
C2503 a_16243_2049# VGND 1.4551f
C2504 a_15119_1793# VGND 1.28484f
C2505 a_15904_1767# VGND 0.53144f
C2506 a_14179_2049# VGND 1.46678f
C2507 a_13167_1793# VGND 1.23052f
C2508 a_13840_1767# VGND 0.53063f
C2509 a_12227_2049# VGND 1.46549f
C2510 a_11175_1793# VGND 1.25081f
C2511 a_11888_1767# VGND 0.53079f
C2512 a_10235_2049# VGND 1.46621f
C2513 a_9223_1793# VGND 1.23055f
C2514 a_9896_1767# VGND 0.53063f
C2515 a_8283_2049# VGND 1.46549f
C2516 a_7221_1787# VGND 1.25589f
C2517 a_7944_1767# VGND 0.53132f
C2518 a_6281_2043# VGND 1.46554f
C2519 a_5269_1787# VGND 1.22942f
C2520 a_5942_1761# VGND 0.53013f
C2521 a_4329_2043# VGND 1.46531f
C2522 a_3990_1761# VGND 0.5313f
C2523 a_3199_1791# VGND 1.29168f
C2524 a_3010_2157# VGND 0.00242f
C2525 a_2676_2157# VGND 0.20473f
C2526 a_2313_2157# VGND 0.21441f
C2527 a_2145_2157# VGND 0.0024f
C2528 a_2049_2157# VGND 0.00314f
C2529 a_1868_1791# VGND 0.1642f
C2530 a_2259_2047# VGND 1.46637f
C2531 a_1920_1765# VGND 0.54304f
C2532 a_2187_1765# VGND 3.37991f
C2533 a_17544_4529# VGND 0
C2534 a_17210_4529# VGND 0.01738f
C2535 a_16847_4529# VGND 0.01904f
C2536 a_18839_4938# VGND 0
C2537 a_18553_4938# VGND 0
C2538 a_15522_4547# VGND 0
C2539 a_15188_4547# VGND 0.01467f
C2540 a_14825_4547# VGND 0.02052f
C2541 a_14657_4547# VGND 0
C2542 a_14561_4547# VGND 0
C2543 a_17544_4895# VGND 0.00238f
C2544 a_17210_4895# VGND 0.20252f
C2545 a_16847_4895# VGND 0.21482f
C2546 a_16679_4895# VGND 0.00207f
C2547 a_16583_4895# VGND 0.0029f
C2548 a_16402_4529# VGND 0.14149f
C2549 a_16793_4785# VGND 1.46252f
C2550 a_16454_4503# VGND 0.51858f
C2551 a_15711_4547# VGND 1.21435f
C2552 a_13520_4553# VGND 0
C2553 a_13186_4553# VGND 0.01746f
C2554 a_12823_4553# VGND 0.01889f
C2555 a_15522_4913# VGND 0.00221f
C2556 a_15188_4913# VGND 0.19864f
C2557 a_14825_4913# VGND 0.21708f
C2558 a_14657_4913# VGND 0.00233f
C2559 a_14561_4913# VGND 0.00306f
C2560 a_14380_4547# VGND 0.1495f
C2561 a_14771_4803# VGND 1.45136f
C2562 a_14432_4521# VGND 0.53166f
C2563 a_13709_4553# VGND 1.22178f
C2564 a_11250_4597# VGND 0
C2565 a_10916_4597# VGND 0.01491f
C2566 a_10553_4597# VGND 0.01744f
C2567 a_10385_4597# VGND 0
C2568 a_10289_4597# VGND 0
C2569 a_13520_4919# VGND 0.00245f
C2570 a_13186_4919# VGND 0.20276f
C2571 a_12823_4919# VGND 0.21461f
C2572 a_12655_4919# VGND 0.00207f
C2573 a_12559_4919# VGND 0.0029f
C2574 a_12378_4553# VGND 0.14264f
C2575 a_12769_4809# VGND 1.46426f
C2576 a_12430_4527# VGND 0.51961f
C2577 a_11439_4597# VGND 1.26233f
C2578 a_11250_4963# VGND 0.00219f
C2579 a_10916_4963# VGND 0.19899f
C2580 a_10553_4963# VGND 0.21133f
C2581 a_10385_4963# VGND 0.00223f
C2582 a_10289_4963# VGND 0.00325f
C2583 a_10108_4597# VGND 0.18458f
C2584 a_10499_4853# VGND 1.43509f
C2585 a_10160_4571# VGND 0.54628f
C2586 a_9128_5049# VGND 0
C2587 a_8794_5049# VGND 0.01792f
C2588 a_8431_5049# VGND 0.02049f
C2589 a_8263_5049# VGND 0
C2590 a_8167_5049# VGND 0
C2591 a_18846_5265# VGND 0.00346f
C2592 a_18625_5265# VGND 0.00367f
C2593 a_18625_4938# VGND 0.30751f
C2594 a_17733_4529# VGND 0.64714f
C2595 a_18371_4938# VGND 0.36105f
C2596 a_17236_5473# VGND 0
C2597 a_16902_5473# VGND 0.02117f
C2598 a_16539_5473# VGND 0.0211f
C2599 a_16371_5473# VGND 0
C2600 a_16275_5473# VGND 0
C2601 a_17425_5473# VGND 1.04149f
C2602 a_15242_5467# VGND 0
C2603 a_14908_5467# VGND 0.01858f
C2604 a_14545_5467# VGND 0.02292f
C2605 a_14377_5467# VGND 0
C2606 a_14281_5467# VGND 0
C2607 a_17236_5839# VGND 0.00267f
C2608 a_16902_5839# VGND 0.20496f
C2609 a_16539_5839# VGND 0.21767f
C2610 a_16371_5839# VGND 0.00238f
C2611 a_16275_5839# VGND 0.0031f
C2612 a_16094_5473# VGND 0.14905f
C2613 a_13284_5459# VGND 0
C2614 a_12950_5459# VGND 0.02272f
C2615 a_12587_5459# VGND 0.02074f
C2616 a_12419_5459# VGND 0
C2617 a_12323_5459# VGND 0
C2618 a_15242_5833# VGND 0.00246f
C2619 a_14908_5833# VGND 0.20339f
C2620 a_14545_5833# VGND 0.21882f
C2621 a_14377_5833# VGND 0.00261f
C2622 a_14281_5833# VGND 0.00325f
C2623 a_14100_5467# VGND 0.1613f
C2624 a_13473_5459# VGND 0.17099f
C2625 a_11222_5471# VGND 0
C2626 a_10888_5471# VGND 0.10793f
C2627 a_10525_5471# VGND 0.10701f
C2628 a_10357_5471# VGND 0
C2629 a_10261_5471# VGND 0
C2630 a_13284_5825# VGND 0.00274f
C2631 a_12950_5825# VGND 0.20604f
C2632 a_12587_5825# VGND 0.21777f
C2633 a_12419_5825# VGND 0.00238f
C2634 a_12323_5825# VGND 0.00309f
C2635 a_12142_5459# VGND 0.14936f
C2636 a_16485_5729# VGND 1.49806f
C2637 a_15431_5467# VGND 1.21826f
C2638 a_16146_5447# VGND 0.53334f
C2639 a_14491_5723# VGND 1.47276f
C2640 a_14419_5441# VGND 0.9778f
C2641 a_14152_5441# VGND 0.55038f
C2642 a_12533_5715# VGND 1.49467f
C2643 a_12194_5433# VGND 0.53334f
C2644 a_11411_5471# VGND 1.25016f
C2645 a_9317_5049# VGND 4.06732f
C2646 a_7126_5043# VGND 0
C2647 a_6792_5043# VGND 0.01675f
C2648 a_6429_5043# VGND 0.02015f
C2649 a_6261_5043# VGND 0
C2650 a_6165_5043# VGND 0
C2651 a_9128_5415# VGND 0.00245f
C2652 a_8794_5415# VGND 0.20264f
C2653 a_8431_5415# VGND 0.21692f
C2654 a_8263_5415# VGND 0.00232f
C2655 a_8167_5415# VGND 0.00307f
C2656 a_7986_5049# VGND 0.14823f
C2657 a_5174_5043# VGND 0
C2658 a_4840_5043# VGND 0.01675f
C2659 a_4477_5043# VGND 0.02018f
C2660 a_4309_5043# VGND 0
C2661 a_4213_5043# VGND 0
C2662 a_7126_5409# VGND 0.00244f
C2663 a_6792_5409# VGND 0.20224f
C2664 a_6429_5409# VGND 0.21685f
C2665 a_6261_5409# VGND 0.00234f
C2666 a_6165_5409# VGND 0.00308f
C2667 a_5984_5043# VGND 0.14749f
C2668 a_3040_5051# VGND 0
C2669 a_2706_5051# VGND 0.01704f
C2670 a_2343_5051# VGND 0.02075f
C2671 a_2175_5051# VGND 0
C2672 a_2079_5051# VGND 0
C2673 a_5174_5409# VGND 0.00247f
C2674 a_4840_5409# VGND 0.20252f
C2675 a_4477_5409# VGND 0.21723f
C2676 a_4309_5409# VGND 0.00233f
C2677 a_4213_5409# VGND 0.00308f
C2678 a_4032_5043# VGND 0.1494f
C2679 a_8377_5305# VGND 1.47482f
C2680 a_7315_5043# VGND 1.25819f
C2681 a_8038_5023# VGND 0.53153f
C2682 a_6375_5299# VGND 1.46572f
C2683 a_5363_5043# VGND 1.23026f
C2684 a_6036_5017# VGND 0.53057f
C2685 a_4423_5299# VGND 1.46661f
C2686 a_4084_5017# VGND 0.5324f
C2687 a_3229_5051# VGND 1.32496f
C2688 a_3040_5417# VGND 0.00243f
C2689 a_2706_5417# VGND 0.20241f
C2690 a_2343_5417# VGND 0.21713f
C2691 a_2175_5417# VGND 0.0024f
C2692 a_2079_5417# VGND 0.00312f
C2693 a_1898_5051# VGND 0.16186f
C2694 a_2289_5307# VGND 1.46694f
C2695 a_1950_5025# VGND 0.54265f
C2696 a_11222_5837# VGND 0.00261f
C2697 a_10888_5837# VGND 0.23876f
C2698 a_10525_5837# VGND 0.27025f
C2699 a_10357_5837# VGND 0.00294f
C2700 a_10261_5837# VGND 0.00349f
C2701 a_10080_5471# VGND 0.19211f
C2702 a_10471_5727# VGND 1.73075f
C2703 a_10132_5445# VGND 0.65067f
C2704 a_2217_5025# VGND 3.40166f
C2705 a_9589_10581# VGND 0.00699f
C2706 a_4723_10577# VGND 0.00697f
C2707 a_9503_10581# VGND 0.41388f
C2708 a_4637_10577# VGND 0.41376f
C2709 a_9631_11297# VGND 0.0104f
C2710 a_4765_11293# VGND 0.0104f
C2711 a_9631_11547# VGND 0.11016f
C2712 a_9463_11547# VGND 0.00246f
C2713 a_4765_11543# VGND 0.11016f
C2714 a_4597_11543# VGND 0.00246f
C2715 a_9381_11547# VGND 0.67614f
C2716 a_4515_11543# VGND 0.67611f
C2717 a_10955_11939# VGND 0.00634f
C2718 a_6089_11935# VGND 0.00634f
C2719 a_9579_12145# VGND 0.00681f
C2720 a_10869_11939# VGND 0.40486f
C2721 a_9771_12117# VGND 1.21463f
C2722 a_4713_12141# VGND 0.00681f
C2723 a_6003_11935# VGND 0.40484f
C2724 a_4905_12113# VGND 1.21953f
C2725 a_9493_12145# VGND 0.40968f
C2726 a_4627_12141# VGND 0.40967f
C2727 a_10995_12931# VGND 0.00334f
C2728 a_10923_12931# VGND 0.00447f
C2729 a_9621_12861# VGND 0.00877f
C2730 a_6129_12927# VGND 0.00334f
C2731 a_6057_12927# VGND 0.00447f
C2732 a_4755_12857# VGND 0.00877f
C2733 a_9621_13111# VGND 0.02732f
C2734 a_9453_13111# VGND 0.00177f
C2735 a_9371_13111# VGND 0.50789f
C2736 a_10841_12931# VGND 0.48715f
C2737 a_4755_13107# VGND 0.02732f
C2738 a_4587_13107# VGND 0.00177f
C2739 a_4505_13107# VGND 0.50789f
C2740 a_5975_12927# VGND 0.48715f
C2741 a_11810_13649# VGND 0
C2742 a_11195_12931# VGND 0.66309f
C2743 a_11728_13649# VGND 0.2862f
C2744 a_10993_13773# VGND 0.00435f
C2745 a_10887_13773# VGND 0.0051f
C2746 a_10799_13773# VGND 0.00448f
C2747 a_9587_13813# VGND 0.00661f
C2748 a_12865_14007# VGND 0
C2749 a_12793_14007# VGND 0
C2750 a_12697_14007# VGND 0
C2751 a_11979_13399# VGND 0.68151f
C2752 a_11147_11911# VGND 1.75603f
C2753 a_9781_10553# VGND 4.42967f
C2754 a_12615_14007# VGND 0.39508f
C2755 a_11255_13773# VGND 0.58592f
C2756 a_10717_13773# VGND 0.49652f
C2757 a_9779_13785# VGND 1.449f
C2758 a_6944_13645# VGND 0
C2759 a_6329_12927# VGND 0.66309f
C2760 a_6862_13645# VGND 0.28619f
C2761 a_6127_13769# VGND 0.00435f
C2762 a_6021_13769# VGND 0.0051f
C2763 a_5933_13769# VGND 0.00448f
C2764 a_4721_13809# VGND 0.00661f
C2765 a_7999_14003# VGND 0
C2766 a_7927_14003# VGND 0
C2767 a_7831_14003# VGND 0
C2768 a_7113_13395# VGND 0.68113f
C2769 a_6281_11907# VGND 1.75628f
C2770 a_4915_10549# VGND 4.31757f
C2771 a_7749_14003# VGND 0.39537f
C2772 a_6389_13769# VGND 0.58592f
C2773 a_9501_13813# VGND 0.4112f
C2774 a_5851_13769# VGND 0.49652f
C2775 a_4913_13781# VGND 1.45376f
C2776 a_4635_13809# VGND 0.41276f
C2777 a_24318_14385# VGND 0.11977f
C2778 a_24152_14385# VGND 0.24786f
C2779 a_23677_14335# VGND 0.00194f
C2780 a_23511_14335# VGND 0.27853f
C2781 a_24962_14701# VGND 0.3508f
C2782 a_24774_14701# VGND 0.28066f
C2783 a_24234_14385# VGND 0.09472f
C2784 a_24241_14651# VGND 0.00666f
C2785 sky130_fd_sc_hd__mux4_1_0.A2 VGND 12.6154f
C2786 sky130_fd_sc_hd__mux4_1_0.A3 VGND 12.5454f
C2787 a_9629_14529# VGND 0.00834f
C2788 a_4763_14525# VGND 0.00834f
C2789 a_23731_14309# VGND 0.45844f
C2790 a_23677_14701# VGND 0.00775f
C2791 a_23511_14701# VGND 0.03067f
C2792 a_10761_14767# VGND 0.00739f
C2793 a_9629_14779# VGND 0.02799f
C2794 a_9461_14779# VGND 0.00172f
C2795 a_5895_14763# VGND 0.00739f
C2796 a_9379_14779# VGND 0.50862f
C2797 a_9705_12861# VGND 3.42826f
C2798 a_4763_14775# VGND 0.02799f
C2799 a_4595_14775# VGND 0.00172f
C2800 a_4513_14775# VGND 0.50862f
C2801 a_4839_12857# VGND 3.43216f
C2802 a_10675_14767# VGND 0.4031f
C2803 a_5809_14763# VGND 0.40306f
C2804 a_11777_15239# VGND 0.00388f
C2805 a_11671_15239# VGND 0.00341f
C2806 a_11583_15239# VGND 0.0016f
C2807 a_12039_15239# VGND 1.08912f
C2808 a_9577_15377# VGND 0.00661f
C2809 a_6911_15235# VGND 0.00388f
C2810 a_6805_15235# VGND 0.00341f
C2811 a_6717_15235# VGND 0.0016f
C2812 a_11501_15239# VGND 0.30451f
C2813 a_10953_14739# VGND 0.7804f
C2814 a_9713_14529# VGND 1.04741f
C2815 a_8193_13753# VGND 2.99982f
C2816 a_9769_15349# VGND 1.95556f
C2817 a_7173_15235# VGND 1.09008f
C2818 a_4711_15373# VGND 0.00661f
C2819 a_6635_15235# VGND 0.30451f
C2820 a_6087_14735# VGND 0.77977f
C2821 a_4847_14525# VGND 1.05454f
C2822 a_4903_15345# VGND 1.95885f
C2823 a_9491_15377# VGND 0.41115f
C2824 a_4625_15373# VGND 0.41117f
C2825 a_9619_16093# VGND 0.00773f
C2826 a_4753_16089# VGND 0.00773f
C2827 a_22274_16171# VGND 0.70974f
C2828 a_21506_16181# VGND 0.64559f
C2829 a_20384_16179# VGND 0.77824f
C2830 a_19510_16177# VGND 0.70725f
C2831 a_18742_16187# VGND 0.64249f
C2832 a_18128_16189# VGND 0.58889f
C2833 a_17254_16187# VGND 0.70665f
C2834 a_16486_16197# VGND 0.65717f
C2835 a_9703_16093# VGND 2.28703f
C2836 a_9619_16343# VGND 0.01843f
C2837 a_9451_16343# VGND 0.00117f
C2838 a_4837_16089# VGND 2.38983f
C2839 a_4753_16339# VGND 0.01843f
C2840 a_4585_16339# VGND 0.00117f
C2841 a_9369_16343# VGND 0.49623f
C2842 a_4503_16339# VGND 0.49694f
C2843 a_6629_15387# VGND 2.82353f
C2844 sky130_fd_sc_hd__mux4_1_0.A1 VGND 9.00165f
.ends

