* NGSPICE file created from tt_um_ohmy90_flat_adders.ext - technology: sky130A

.subckt tt_um_ohmy90_flat_adders clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5]
+ ua[6] ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7]
+ uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
+ uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
+ uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
+ VDPWR VGND
X0 a_4183_1787# a_4129_2043# a_3790_1761# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X1 a_15255_4841# a_14325_4589# a_15672_4585# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X2 a_24234_14385# ui_in[0] a_24152_14385# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.10855 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X3 VGND a_14888_5433# a_14836_5459# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X4 a_15113_5825# VDPWR a_15017_5825# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X5 a_13732_1769# VGND VDPWR w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X6 a_4711_15373# VGND a_4625_15373# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X7 a_11202_5441# a_10611_5471# a_11427_5467# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X8 VDPWR VGND a_2313_1791# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X9 VGND a_5636_5017# a_5584_5043# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X10 a_9865_15329# a_9587_15357# VDPWR w_9490_15543# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X11 a_1950_5025# a_2217_5025# a_2175_5051# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X12 VDPWR VDPWR a_15644_5459# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X13 a_5999_1783# a_5069_1787# VDPWR w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X14 VDPWR VDPWR a_9587_15357# w_9490_15543# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X15 a_4513_14775# VDPWR VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X16 a_6129_12927# a_4913_13781# a_6057_12927# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=1764,126
X17 VDPWR VDPWR a_6392_5043# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X18 a_11623_4959# a_11569_4849# a_11230_4567# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X19 VDPWR VDPWR a_11595_5467# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X20 sky130_fd_sc_hd__mux4_1_0.A3 a_17125_4938# VDPWR w_16764_4814# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=6334,279 d=10400,504
X21 a_13802_4955# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X22 a_7113_13395# a_6862_13645# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4010,197 d=6760,364
X23 VDPWR VGND a_15239_1765# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X24 a_3820_5021# a_3229_5051# a_4045_5413# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X25 VDPWR VGND a_4587_13107# w_4432_13071# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X26 a_13439_4955# a_12509_4593# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X27 a_15045_4951# a_14946_4905# a_14946_4905# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.07384 ps=0.80236 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X28 a_22274_16171# a_21506_16181# VDPWR w_22086_16385# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X29 a_2175_5417# VDPWR a_2079_5417# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X30 a_6089_11935# a_4849_11293# a_6003_11935# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X31 VDPWR VGND a_4597_11543# w_4442_11507# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X32 VDPWR a_9867_12097# a_10965_11919# w_10868_12105# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X33 a_14946_4905# a_14946_4905# a_15309_4951# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.07384 pd=0.80236 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X34 a_17346_5265# a_16195_4585# a_17125_4938# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
**devattr s=3990,179 d=2772,150
X35 VGND VGND a_9467_13091# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X36 a_15936_2131# VDPWR a_15185_2021# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X37 VGND VDPWR a_4213_5413# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X38 a_9671_5727# VGND a_10088_5471# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X39 a_11553_1773# a_11499_2029# a_11160_1747# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X40 a_13774_5463# VGND VDPWR w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X41 a_3949_5047# VGND VDPWR w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X42 VGND VGND a_8566_2145# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X43 a_9715_16323# VGND VDPWR w_9392_16287# sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X44 a_9725_14509# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X45 VGND a_1920_1765# a_1868_1791# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X46 VDPWR a_12075_13379# a_12881_13987# w_12566_13951# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=5930,268
X47 a_10422_5837# VDPWR a_9671_5727# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X48 VDPWR sky130_fd_sc_hd__mux4_1_0.A1 a_6629_15387# w_9392_17212# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X49 VDPWR VDPWR a_4753_16339# w_4430_16303# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X50 a_9332_5445# VGND a_9557_5837# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X51 VDPWR a_5606_1757# a_5554_1783# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X52 VDPWR a_12976_1743# a_12924_1769# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X53 a_4880_1787# VDPWR a_4129_2043# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X54 a_5945_2039# a_5069_1787# a_6362_2149# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X55 a_12509_4593# a_11569_4849# VDPWR w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X56 a_11359_4959# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X57 VGND VDPWR a_4546_2153# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X58 a_4903_15345# a_4625_15373# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X59 a_11541_5723# a_10611_5471# a_11958_5833# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X60 a_11230_4567# a_10639_4597# a_11455_4593# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X61 a_15644_5825# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X62 a_7476_1753# a_6885_1783# a_7701_2145# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X63 VDPWR VDPWR a_4763_14775# w_4440_14739# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X64 a_11291_12911# a_10937_12911# VDPWR w_10872_13125# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5689,267 d=10400,504
X65 a_8232_2145# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X66 a_7869_1779# a_7815_2035# a_7476_1753# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X67 a_5831_2149# VDPWR a_5735_2149# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X68 a_4913_13781# a_4635_13809# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X69 a_10813_13753# a_9799_16073# VDPWR w_10748_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X70 a_5735_1783# VGND VDPWR w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X71 VGND VDPWR a_9725_5837# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X72 VDPWR a_11202_5441# a_11150_5467# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X73 a_11499_2029# a_10569_1777# a_11916_2139# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X74 a_11986_4593# VGND VDPWR w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X75 VDPWR VDPWR a_9727_11527# w_9404_11491# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X76 a_9753_4597# VDPWR VDPWR w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X77 a_4723_10577# VGND a_4637_10577# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X78 VDPWR VDPWR a_11623_4593# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X79 a_4587_13107# VDPWR a_4505_13107# w_4432_13071# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X80 a_2079_5051# VGND VDPWR w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X81 VGND a_9360_4571# a_9308_4597# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X82 VDPWR VDPWR a_9599_10561# w_9502_10747# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X83 a_11331_5467# VGND VDPWR w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X84 a_4597_11543# VDPWR a_4515_11543# w_4442_11507# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X85 a_6944_13645# a_6329_12927# a_6862_13645# w_6756_13609# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X86 a_7669_14003# a_7173_15235# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X87 a_9467_13091# VDPWR VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X88 a_16195_4585# a_15255_4841# a_14946_4905# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.11427 ps=1.24175 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X89 VDPWR VGND a_11595_5467# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X90 a_4635_13809# VGND VDPWR w_4538_13995# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X91 a_2706_5417# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X92 VDPWR VGND a_2343_5051# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X93 a_15281_5459# a_14297_5463# VDPWR w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X94 VGND a_4513_14775# a_4847_14525# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X95 a_5975_5299# a_5099_5047# a_6392_5409# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X96 VGND a_4503_16339# a_4837_16089# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X97 VGND a_9475_14759# a_9809_14509# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X98 a_13315_2025# a_12439_1773# a_13732_2135# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X99 VGND VDPWR a_4576_5413# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X100 VGND VGND a_10422_5837# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X101 a_6029_5043# a_5975_5299# a_5636_5017# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X102 a_12135_15219# a_11597_15219# VDPWR w_11532_15433# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X103 a_15602_2131# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X104 VDPWR VGND a_4880_1787# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X105 VGND a_8785_5039# a_16871_4938# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=5796,222
X106 a_11385_1773# VDPWR a_11289_1773# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X107 VGND sky130_fd_sc_hd__mux4_1_0.A1 a_23511_14335# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X108 VGND VGND a_4213_5413# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X109 VDPWR VGND a_14136_4589# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X110 VGND VGND a_15978_5825# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X111 a_6805_15235# a_4847_14525# a_6717_15235# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X112 a_7899_5405# a_6915_5043# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X113 VDPWR VDPWR a_13411_5463# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X114 a_15239_2131# a_14255_1769# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X115 a_9727_11527# VGND VDPWR w_9404_11491# sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X116 a_1920_1765# a_2187_1765# a_2145_2157# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X117 a_14325_4589# a_13385_4845# VDPWR w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X118 VDPWR a_11230_4567# a_11178_4593# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X119 VGND VDPWR a_9753_4963# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X120 a_16486_16197# sky130_fd_sc_hd__mux4_1_0.A0 VDPWR w_16298_16411# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X121 a_4546_1787# VGND VDPWR w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X122 a_23677_14701# ui_in[0] ui_in[1] sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.36 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=4316,272
X123 a_4905_12113# a_4627_12141# VDPWR w_4530_12327# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X124 a_4915_10549# a_4637_10577# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X125 a_9461_5837# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X126 a_14888_5433# a_14297_5463# a_15113_5825# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X127 a_7815_2035# a_6885_1783# a_8232_1779# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X128 a_7605_2145# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X129 VDPWR a_9809_14509# a_11597_15219# w_11532_15433# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X130 a_6087_14735# a_5809_14763# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X131 VGND a_6281_11907# a_7669_14003# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2772,150 d=2268,138
X132 VGND VDPWR a_2313_2157# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X133 VGND VDPWR a_11958_5833# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X134 a_13243_5829# VDPWR a_13147_5829# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X135 a_9683_2143# a_9629_2033# a_9290_1751# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X136 VGND VGND a_9725_5837# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X137 a_15672_4585# a_14946_4905# VDPWR w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X138 a_13411_5463# a_13357_5719# a_13018_5437# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X139 VDPWR VGND a_3010_1791# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X140 a_4183_2153# a_3199_1791# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X141 a_5099_5047# a_4159_5303# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X142 a_11553_2139# a_10569_1777# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X143 VDPWR VGND a_11623_4593# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X144 a_4763_14525# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X145 a_15309_4585# a_14325_4589# VDPWR w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X146 a_24962_14701# ui_in[1] a_24234_14385# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.15102 pd=1.285 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=6041,257
X147 a_4045_5047# VDPWR a_3949_5047# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X148 a_2259_2047# a_2187_1765# a_2676_1791# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X149 VDPWR VGND a_13369_1769# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X150 a_6696_1783# VDPWR a_5945_2039# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X151 VDPWR a_9290_1751# a_9238_1777# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X152 a_1950_5025# a_2217_5025# a_2175_5417# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X153 a_12631_13987# a_9877_10533# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4368,272 d=2772,150
X154 a_9589_12125# VGND VDPWR w_9492_12311# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X155 a_11906_13629# a_11291_12911# a_11824_13629# w_11718_13593# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X156 VGND VDPWR a_6392_5409# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X157 sky130_fd_sc_hd__mux4_1_0.A2 a_15185_2021# VDPWR w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X158 a_9753_4597# a_9699_4853# a_9360_4571# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X159 VDPWR a_13018_5437# a_12966_5463# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X160 VGND VDPWR a_13732_2135# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X161 a_6915_5043# a_5975_5299# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X162 a_7635_5405# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X163 a_12292_5467# VDPWR a_11541_5723# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X164 a_14946_4905# a_14946_4905# a_16006_4951# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.07384 pd=0.80236 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X165 a_14975_2131# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X166 a_15185_2021# a_14255_1769# a_15602_1765# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X167 VDPWR VGND a_9547_16323# w_9392_16287# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X168 a_3040_5051# VDPWR a_2289_5307# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X169 a_13201_1769# VDPWR a_13105_1769# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X170 a_8755_1779# a_7815_2035# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X171 a_5895_14763# a_4849_11293# a_5809_14763# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X172 VGND VGND a_9475_14759# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X173 VGND VGND a_7899_5405# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X174 VDPWR a_3790_1761# a_3738_1787# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X175 VGND VDPWR a_4711_15373# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X176 VDPWR a_9801_12841# a_10771_14747# w_10674_14933# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X177 a_5861_5043# VDPWR a_5765_5043# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X178 a_13147_5463# VGND VDPWR w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X179 VDPWR a_9799_16073# a_11597_15219# w_11532_15433# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X180 a_14916_4559# a_14325_4589# a_15141_4951# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X181 a_5069_1787# a_4129_2043# VDPWR w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X182 a_10639_4597# a_9699_4853# VDPWR w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X183 VGND VDPWR a_2676_2157# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X184 a_13271_4955# VDPWR a_13175_4955# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X185 VGND VGND a_4513_14775# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X186 a_9671_5727# VGND a_10088_5837# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X187 VDPWR a_14916_4559# a_14864_4585# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X188 a_11051_11919# a_9811_11277# a_10965_11919# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X189 a_13774_5829# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X190 a_3790_1761# a_3199_1791# a_4015_1787# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X191 VDPWR VDPWR a_13802_4589# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X192 VDPWR VDPWR a_8232_1779# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X193 a_11351_13753# a_10813_13753# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X194 VGND VGND a_2313_2157# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X195 VDPWR a_11351_13753# a_11906_13629# w_11718_13593# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5830,267
X196 a_9515_2143# VDPWR a_9419_2143# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X197 ua[0] a_24962_14701# VDPWR sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X198 a_4755_13107# VGND VDPWR w_4432_13071# sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X199 VDPWR VGND a_6696_1783# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X200 a_5999_2149# a_5069_1787# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X201 VDPWR VDPWR a_4183_1787# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X202 a_5933_13769# a_4849_11293# a_5851_13769# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
X203 a_9673_15357# VGND a_9587_15357# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X204 a_4576_5047# VGND VDPWR w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X205 VGND VGND a_15281_5825# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X206 VGND a_11160_1747# a_11108_1773# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X207 a_11230_4567# a_10639_4597# a_11455_4959# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X208 a_11597_15219# a_8113_13753# VDPWR w_11532_15433# sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X209 a_4765_11543# VGND VDPWR w_4442_11507# sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X210 a_21506_16181# a_20384_16179# VDPWR w_21318_16395# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X211 a_6885_1783# a_5945_2039# VDPWR w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X212 a_9683_13793# VGND a_9597_13793# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X213 VDPWR VGND a_12292_5467# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X214 a_9547_16323# VDPWR a_9465_16323# w_9392_16287# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X215 a_4503_16339# VDPWR VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X216 a_5606_1757# a_5069_1787# a_5831_1783# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X217 a_11986_4959# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X218 a_9475_14759# VDPWR VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X219 a_4015_2153# VDPWR a_3919_2153# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X220 a_17339_4938# a_16167_5459# a_17125_4938# w_16764_4814# sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1932 ps=1.34 w=0.42 l=0.15
**devattr s=7728,268 d=3066,157
X221 VDPWR VGND a_3040_5051# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X222 a_11595_5833# a_11541_5723# a_11202_5441# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X223 a_6362_1783# VGND VDPWR w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X224 a_12320_4593# VDPWR a_11569_4849# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X225 VGND VDPWR a_11623_4959# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X226 VDPWR VDPWR a_9715_16323# w_9392_16287# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X227 a_10771_14747# a_9811_11277# VDPWR w_10674_14933# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X228 a_9809_14509# VDPWR a_9725_14509# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X229 a_2079_5417# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X230 a_3229_5051# a_2289_5307# VDPWR w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X231 a_9629_2033# a_8755_1779# a_10046_1777# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X232 VGND sky130_fd_sc_hd__mux4_1_0.A3 a_2217_5025# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X233 a_12481_5467# a_11541_5723# VDPWR w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X234 a_12439_1773# a_11499_2029# VDPWR w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X235 a_15309_4585# a_15255_4841# a_14916_4559# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X236 a_9585_4597# VDPWR a_9489_4597# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X237 a_11553_2139# a_11499_2029# a_11160_1747# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X238 a_11160_1747# a_10569_1777# a_11385_1773# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X239 a_14066_1769# VDPWR a_13315_2025# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X240 VGND a_7476_1753# a_7424_1779# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X241 a_2289_5307# a_2217_5025# a_2706_5051# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X242 a_15978_5459# VDPWR a_15227_5715# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X243 ui_in[1] a_23731_14309# a_23677_14335# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.09322 pd=1.07 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3409,185
X244 a_6389_13769# a_5851_13769# VDPWR w_5786_13983# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X245 a_11958_5467# VGND VDPWR w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X246 VDPWR a_4903_15345# a_5851_13769# w_5786_13983# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X247 VGND VGND a_2343_5417# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X248 VDPWR VDPWR a_15602_1765# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X249 a_7751_14003# a_4915_10549# a_7669_14003# w_7604_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2772,150
X250 VDPWR VGND a_9559_11527# w_9404_11491# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X251 a_16167_5459# a_15227_5715# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X252 VDPWR VDPWR a_2343_5051# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X253 a_9683_1777# a_8755_1779# VDPWR w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X254 a_9699_4853# VDPWR a_10116_4963# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X255 VGND VDPWR a_4723_10577# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X256 a_13369_2135# a_12439_1773# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X257 a_4625_15373# VGND VDPWR w_4528_15559# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X258 a_14136_4955# VDPWR a_13385_4845# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X259 a_19510_16177# a_18742_16187# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X260 a_11049_14719# a_10771_14747# VDPWR w_10674_14933# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X261 a_4159_5303# a_3229_5051# a_4576_5413# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X262 a_6029_5409# a_5975_5299# a_5636_5017# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X263 a_14946_4905# VDPWR a_15672_4951# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.07384 pd=0.80236 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X264 a_8596_5405# VDPWR a_7845_5295# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X265 a_5735_2149# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X266 a_24774_14701# ui_in[1] VDPWR sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X267 VDPWR a_3820_5021# a_3768_5047# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X268 a_18742_16187# a_18128_16189# VDPWR w_18554_16401# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X269 a_9865_15329# a_9587_15357# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X270 VDPWR VDPWR a_4635_13809# w_4538_13995# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X271 VGND VDPWR a_13411_5829# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X272 a_14108_5463# VDPWR a_13357_5719# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X273 a_9875_13765# a_9597_13793# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X274 a_10569_1777# a_9629_2033# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X275 VDPWR VGND a_4183_1787# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X276 a_17125_4938# a_16195_4585# a_17053_4938# w_16764_4814# sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=7728,268
X277 VDPWR VGND a_12320_4593# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X278 a_11291_12911# a_10937_12911# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=5266,228 d=6760,364
X279 VGND a_7506_5013# a_7454_5039# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X280 VDPWR sky130_fd_sc_hd__mux4_1_0.A1 a_23511_14701# sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X281 a_8113_13753# a_7669_14003# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4075,198 d=7020,368
X282 VGND a_14846_1739# a_14794_1765# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X283 a_15071_2131# VDPWR a_14975_2131# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X284 VDPWR sky130_fd_sc_hd__mux4_1_0.A2 a_2187_1765# w_6044_2758# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X285 VGND a_13046_4563# a_12994_4589# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X286 sky130_fd_sc_hd__mux4_1_0.A0 a_22274_16171# VDPWR w_22960_16387# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X287 ui_in[1] a_24774_14701# a_24962_14701# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.09322 pd=1.07 as=0.15102 ps=1.285 w=0.42 l=0.15
**devattr s=6041,257 d=4368,272
X288 a_6057_12927# a_4849_11293# a_5975_12927# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X289 a_9725_5471# VGND VDPWR w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X290 a_7869_1779# a_6885_1783# VDPWR w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X291 a_3199_1791# a_2259_2047# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X292 VDPWR VDPWR a_8262_5039# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X293 a_23677_14335# sky130_fd_sc_hd__mux4_1_0.A0 VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X294 VDPWR VGND a_14066_1769# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X295 a_13411_5829# a_13357_5719# a_13018_5437# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X296 VGND a_6389_13769# a_6862_13645# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4010,197
X297 a_9559_11527# VDPWR a_9477_11527# w_9404_11491# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X298 a_11427_5833# VDPWR a_11331_5833# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X299 a_16006_4585# VDPWR a_15255_4841# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X300 VGND VGND a_11623_4959# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X301 a_7919_14003# a_7173_15235# a_7847_14003# w_7604_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X302 a_14255_1769# a_13315_2025# VDPWR w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X303 a_11243_11891# a_10965_11919# VDPWR w_10868_12105# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X304 VDPWR VDPWR a_10046_1777# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X305 a_12976_1743# a_12439_1773# a_13201_1769# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X306 a_2313_1791# a_2187_1765# VDPWR w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X307 a_5975_12927# a_4913_13781# VDPWR w_5910_13141# sky130_fd_pr__pfet_01v8_hvt ad=0.0805 pd=0.94333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2646,147
X308 a_11385_2139# VDPWR a_11289_2139# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X309 VDPWR VDPWR a_2706_5051# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X310 a_11289_1773# VGND VDPWR w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X311 a_4213_5047# a_4159_5303# a_3820_5021# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X312 a_5636_5017# a_5099_5047# a_5861_5043# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X313 VDPWR VDPWR a_5999_1783# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X314 VDPWR VDPWR a_13369_1769# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X315 a_15141_4585# VDPWR a_15045_4585# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X316 VGND VGND a_8596_5405# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X317 a_6392_5043# VGND VDPWR w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X318 VGND a_4837_16089# a_6911_15235# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X319 VGND VGND a_15936_2131# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X320 VGND VDPWR a_10116_4963# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X321 a_13046_4563# a_12509_4593# a_13271_4955# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X322 VDPWR VGND a_11553_1773# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X323 VDPWR VGND a_14108_5463# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X324 a_4847_14525# VDPWR a_4763_14525# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X325 a_6029_5043# a_5099_5047# VDPWR w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X326 VGND VDPWR a_13439_4955# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X327 a_3040_5417# VDPWR a_2289_5307# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X328 a_7506_5013# a_6915_5043# a_7731_5405# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X329 a_8262_5405# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X330 a_10380_2143# VDPWR a_9629_2033# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X331 a_13147_5829# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X332 a_9290_1751# a_8755_1779# a_9515_2143# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X333 a_4713_12141# VGND a_4627_12141# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X334 a_5861_5409# VDPWR a_5765_5409# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X335 a_14297_5463# a_13357_5719# VDPWR w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X336 a_10983_13753# a_9865_15329# a_10895_13753# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X337 a_11089_13753# a_9799_16073# a_10983_13753# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X338 a_13018_5437# a_12481_5467# a_13243_5463# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X339 a_13369_2135# a_13315_2025# a_12976_1743# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X340 VGND VGND a_3010_2157# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X341 a_9867_12097# a_9589_12125# VDPWR w_9492_12311# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X342 a_6717_15235# a_6629_15387# a_6635_15235# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
X343 a_4837_16089# a_4503_16339# a_4753_16339# w_4430_16303# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X344 VDPWR VDPWR a_9589_12125# w_9492_12311# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X345 VDPWR VDPWR a_10088_5471# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X346 a_9877_10533# a_9599_10561# VDPWR w_9502_10747# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X347 VDPWR VGND a_7869_1779# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X348 VGND VDPWR a_9683_2143# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X349 a_2259_2047# a_2187_1765# a_2676_2157# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X350 a_4753_16089# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X351 VDPWR a_4849_11293# a_5975_12927# w_5910_13141# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0805 ps=0.94333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X352 VGND a_4839_12857# a_5895_14763# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X353 a_6696_2149# VDPWR a_5945_2039# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X354 a_15227_5715# a_14297_5463# a_15644_5825# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X355 a_10450_4597# VDPWR a_9699_4853# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X356 VDPWR a_14888_5433# a_14836_5459# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X357 a_9360_4571# VDPWR a_9585_4597# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X358 a_18128_16189# a_17254_16187# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X359 VDPWR a_5636_5017# a_5584_5043# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X360 a_7701_1779# VDPWR a_7605_1779# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X361 a_12135_15219# a_11597_15219# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X362 a_4910_5047# VDPWR a_4159_5303# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X363 a_13439_4589# a_13385_4845# a_13046_4563# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X364 a_11569_4849# a_10639_4597# a_11986_4593# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X365 VGND a_9867_12097# a_11051_11919# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X366 a_13105_1769# VGND VDPWR w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X367 VGND VDPWR a_7869_2145# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X368 a_17125_4938# a_16167_5459# a_17125_5265# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=3990,179
X369 a_15017_5459# VGND VDPWR w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X370 VGND sky130_fd_sc_hd__mux4_1_0.A1 a_6629_15387# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X371 VGND VGND a_3040_5417# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X372 VDPWR VGND a_5999_1783# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X373 a_7899_5039# a_7845_5295# a_7506_5013# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X374 a_11873_15219# a_11049_14719# a_11767_15219# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X375 VDPWR a_9801_12841# a_10813_13753# w_10748_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X376 a_5765_5043# VGND VDPWR w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X377 a_12509_4593# a_11569_4849# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X378 a_12320_4959# VDPWR a_11569_4849# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X379 VGND VGND a_10380_2143# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X380 VGND a_4505_13107# a_4839_12857# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X381 VDPWR VDPWR a_4755_13107# w_4432_13071# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X382 sky130_fd_sc_hd__mux4_1_0.A3 a_17125_4938# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4514,209 d=6760,364
X383 a_10937_12911# a_9875_13765# VDPWR w_10872_13125# sky130_fd_pr__pfet_01v8_hvt ad=0.0805 pd=0.94333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2646,147
X384 a_11595_5467# a_10611_5471# VDPWR w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X385 a_13175_4955# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X386 a_4905_12113# a_4627_12141# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X387 a_2289_5307# a_2217_5025# a_2706_5417# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X388 VDPWR VDPWR a_15281_5459# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X389 VGND VDPWR a_9673_15357# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X390 VDPWR sky130_fd_sc_hd__mux4_1_0.A3 a_24407_14651# sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.09013 ps=0.995 w=0.42 l=0.15
**devattr s=3605,199 d=2268,138
X391 VDPWR VDPWR a_4765_11543# w_4442_11507# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X392 VDPWR a_7113_13395# a_7919_14003# w_7604_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=5930,268
X393 VGND VGND a_13439_4955# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X394 VGND VDPWR a_9683_13793# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X395 a_10046_2143# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X396 VGND VGND a_4503_16339# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X397 VGND VDPWR a_2343_5417# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X398 a_9419_2143# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X399 a_12075_13379# a_11824_13629# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4010,197 d=6760,364
X400 VGND VGND a_6696_2149# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X401 sky130_fd_sc_hd__mux4_1_0.A1 a_12631_13987# VDPWR w_12566_13951# sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5930,268 d=10800,508
X402 a_12250_1773# VDPWR a_11499_2029# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X403 a_4213_5413# a_3229_5051# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X404 a_14846_1739# a_14255_1769# a_15071_2131# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X405 VDPWR VGND a_10450_4597# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X406 VDPWR VDPWR a_13774_5463# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X407 a_15239_1765# a_15185_2021# a_14846_1739# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X408 a_15281_5459# a_15227_5715# a_14888_5433# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X409 a_20384_16179# a_19510_16177# VDPWR w_20196_16393# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X410 VGND VDPWR a_7899_5405# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X411 VGND VDPWR a_15239_2131# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X412 VGND VGND a_9683_2143# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X413 a_15255_4841# a_14325_4589# a_15672_4951# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X414 a_17254_16187# a_16486_16197# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X415 a_6862_13645# a_6329_12927# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X416 VDPWR VGND a_4910_5047# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X417 VDPWR VGND a_13411_5463# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X418 a_5606_1757# a_5069_1787# a_5831_2149# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X419 a_11202_5441# a_10611_5471# a_11427_5833# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X420 a_14108_5829# VDPWR a_13357_5719# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X421 a_6362_2149# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X422 VGND a_5606_1757# a_5554_1783# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X423 a_3919_2153# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X424 a_4129_2043# a_3199_1791# a_4546_1787# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X425 a_5851_13769# a_4849_11293# VDPWR w_5786_13983# sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X426 a_4721_13809# VGND a_4635_13809# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X427 VDPWR a_9865_15329# a_10813_13753# w_10748_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X428 VDPWR a_4847_14525# a_6635_15235# w_6570_15449# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X429 VGND VDPWR a_15644_5825# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X430 a_8566_1779# VDPWR a_7815_2035# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X431 a_10116_4597# VGND VDPWR w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X432 VGND VGND a_12320_4959# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X433 VGND a_9801_12841# a_11089_13753# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X434 a_9489_4597# VGND VDPWR w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X435 VDPWR VDPWR a_4625_15373# w_4528_15559# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X436 a_12631_13987# a_12135_15219# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X437 a_9725_5837# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X438 a_11160_1747# a_10569_1777# a_11385_2139# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X439 a_13385_4845# a_12509_4593# a_13802_4589# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X440 VGND VDPWR a_11595_5833# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X441 VDPWR VDPWR a_11986_4593# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X442 a_7113_13395# a_6862_13645# VDPWR w_6756_13609# sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5830,267 d=13600,536
X443 a_11091_12911# a_9875_13765# a_11019_12911# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=1764,126
X444 a_8785_5039# a_7845_5295# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X445 a_11623_4593# a_10639_4597# VDPWR w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X446 a_7845_5295# a_6915_5043# a_8262_5039# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X447 a_14325_4589# a_13385_4845# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X448 a_9557_5471# VDPWR a_9461_5471# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X449 VDPWR VDPWR a_15309_4585# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X450 VDPWR VGND a_9753_4597# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X451 VDPWR a_8785_5039# a_17339_4938# w_16764_4814# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.07665 ps=0.785 w=0.42 l=0.15
**devattr s=3066,157 d=6334,279
X452 VGND a_11230_4567# a_11178_4593# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X453 a_7731_5039# VDPWR a_7635_5039# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X454 a_24774_14701# ui_in[1] VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X455 VDPWR VGND a_12250_1773# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X456 a_23677_14701# sky130_fd_sc_hd__mux4_1_0.A0 VDPWR sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.36 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X457 VGND VGND a_4505_13107# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X458 VGND VDPWR a_2706_5417# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X459 a_5636_5017# a_5099_5047# a_5861_5409# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X460 a_4183_2153# a_4129_2043# a_3790_1761# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X461 a_3949_5413# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X462 a_6392_5409# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X463 ua[0] a_24962_14701# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X464 a_9801_12841# a_9467_13091# a_9717_13091# w_9394_13055# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X465 a_13732_2135# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X466 a_2145_1791# VDPWR a_2049_1791# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X467 a_6726_5043# VDPWR a_5975_5299# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X468 a_15936_1765# VDPWR a_15185_2021# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X469 a_5809_14763# a_4849_11293# VDPWR w_5712_14949# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X470 a_6029_5409# a_5099_5047# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X471 VGND VGND a_14108_5829# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X472 a_11916_1773# VGND VDPWR w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X473 VGND a_9801_12841# a_11091_12911# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5266,228
X474 VDPWR VDPWR a_11553_1773# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X475 VDPWR VGND a_8566_1779# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X476 a_15113_5459# VDPWR a_15017_5459# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X477 VGND a_11243_11891# a_12631_13987# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2772,150 d=2268,138
X478 VDPWR a_4837_16089# a_6635_15235# w_6570_15449# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X479 VGND VGND a_15239_2131# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X480 a_13018_5437# a_12481_5467# a_13243_5829# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X481 a_8755_1779# a_7815_2035# VDPWR w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X482 a_9753_4963# VDPWR VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X483 VDPWR VDPWR a_4546_1787# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X484 VGND VDPWR a_10088_5837# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X485 a_7476_1753# a_6885_1783# a_7701_1779# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X486 a_13802_4589# VGND VDPWR w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X487 a_12713_13987# a_9877_10533# a_12631_13987# w_12566_13951# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2772,150
X488 a_8232_1779# VGND VDPWR w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X489 a_10611_5471# a_9671_5727# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X490 a_11331_5833# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X491 a_2313_2157# a_2187_1765# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X492 a_11767_15219# a_9809_14509# a_11679_15219# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X493 a_11824_13629# a_11291_12911# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X494 a_5099_5047# a_4159_5303# VDPWR w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X495 a_11289_2139# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X496 VGND a_9332_5445# a_9280_5471# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X497 a_3820_5021# a_3229_5051# a_4045_5047# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X498 VGND VDPWR a_5999_2149# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X499 a_22274_16171# a_21506_16181# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X500 a_10813_13753# a_9811_11277# VDPWR w_10748_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X501 a_4505_13107# VDPWR VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X502 VGND VGND a_11595_5833# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X503 a_13439_4589# a_12509_4593# VDPWR w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X504 a_15045_4585# a_14946_4905# VDPWR w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X505 a_6635_15235# a_6629_15387# VDPWR w_6570_15449# sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X506 VGND VDPWR a_4713_12141# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X507 a_15281_5825# a_14297_5463# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X508 VGND VGND a_4515_11543# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X509 a_10639_4597# a_9699_4853# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X510 VGND a_9801_12841# a_10857_14747# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X511 VDPWR a_14946_4905# a_15309_4585# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X512 a_14946_4905# a_14916_4559# a_14864_4585# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.11427 pd=1.24175 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X513 a_11049_14719# a_10771_14747# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X514 a_9597_13793# VGND VDPWR w_9500_13979# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X515 VGND VGND a_11553_2139# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X516 VDPWR VDPWR a_4213_5047# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X517 VDPWR VGND a_6726_5043# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X518 a_4880_2153# VDPWR a_4129_2043# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X519 a_11569_4849# a_10639_4597# a_11986_4959# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X520 a_9715_16073# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X521 a_2676_1791# VGND VDPWR w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X522 VDPWR a_11160_1747# a_11108_1773# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X523 a_7869_2145# a_7815_2035# a_7476_1753# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X524 a_5765_5409# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X525 VGND VGND a_14136_4955# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X526 a_4837_16089# VDPWR a_4753_16089# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X527 a_6915_5043# a_5975_5299# VDPWR w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X528 a_4913_13781# a_4635_13809# VDPWR w_4538_13995# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X529 VDPWR a_4839_12857# a_5975_12927# w_5910_13141# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0805 ps=0.94333 w=0.42 l=0.15
**devattr s=2646,147 d=5689,267
X530 a_6329_12927# a_5975_12927# VDPWR w_5910_13141# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5689,267 d=10400,504
X531 VGND a_1950_5025# a_1898_5051# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X532 a_13315_2025# a_12439_1773# a_13732_1769# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X533 VDPWR a_9811_11277# a_10937_12911# w_10872_13125# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0805 ps=0.94333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X534 VDPWR VDPWR a_11916_1773# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X535 a_11541_5723# a_10611_5471# a_11958_5467# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X536 a_15644_5459# VGND VDPWR w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X537 a_9675_12125# VGND a_9589_12125# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X538 a_15602_1765# VGND VDPWR w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X539 a_11597_15219# a_11049_14719# VDPWR w_11532_15433# sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X540 a_24234_14385# ui_in[0] a_24241_14651# sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1274 pd=1.16667 as=0.10855 ps=1.36 w=0.42 l=0.15
**devattr s=4316,272 d=2268,138
X541 VDPWR VDPWR a_9717_13091# w_9394_13055# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X542 a_6281_11907# a_6003_11935# VDPWR w_5906_12121# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X543 a_9811_11277# VDPWR a_9727_11277# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X544 VGND a_3790_1761# a_3738_1787# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X545 VDPWR a_4905_12113# a_6003_11935# w_5906_12121# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X546 a_9685_10561# VGND a_9599_10561# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X547 a_15239_1765# a_14255_1769# VDPWR w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X548 VDPWR a_7476_1753# a_7424_1779# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X549 a_4847_14525# a_4513_14775# a_4763_14775# w_4440_14739# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X550 a_5069_1787# a_4129_2043# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X551 a_15672_4951# a_14946_4905# a_14946_4905# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.07384 ps=0.80236 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X552 a_9809_14509# a_9475_14759# a_9725_14759# w_9402_14723# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X553 a_10895_13753# a_9811_11277# a_10813_13753# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
X554 a_4515_11543# VDPWR VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X555 VGND VDPWR a_13774_5829# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X556 a_10857_14747# a_9811_11277# a_10771_14747# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X557 a_7605_1779# VGND VDPWR w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X558 a_7847_14003# a_6281_11907# a_7751_14003# w_7604_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X559 a_15309_4951# a_14325_4589# a_14946_4905# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.07384 ps=0.80236 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X560 a_13357_5719# a_12481_5467# a_13774_5463# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X561 a_9683_1777# a_9629_2033# a_9290_1751# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X562 a_17125_5265# a_16871_4938# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=5796,222 d=2772,150
X563 a_24241_14651# sky130_fd_sc_hd__mux4_1_0.A2 VDPWR sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.10855 pd=1.36 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X564 a_4045_5413# VDPWR a_3949_5413# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X565 VGND VGND a_13411_5829# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X566 VGND VGND a_4880_2153# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X567 VGND a_9465_16323# a_9799_16073# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X568 VGND VGND a_5999_2149# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X569 a_4183_1787# a_3199_1791# VDPWR w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X570 VDPWR VDPWR a_4576_5047# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X571 a_6021_13769# a_4903_15345# a_5933_13769# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X572 VDPWR a_1920_1765# a_1868_1791# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X573 VGND sky130_fd_sc_hd__mux4_1_0.A3 a_24152_14385# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.10855 ps=1.36 w=0.42 l=0.15
**devattr s=4316,272 d=2268,138
X574 a_6127_13769# a_4837_16089# a_6021_13769# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X575 a_4627_12141# VGND VDPWR w_4530_12327# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X576 a_6885_1783# a_5945_2039# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X577 a_9753_4963# a_9699_4853# a_9360_4571# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X578 VDPWR VGND a_4213_5047# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X579 a_12292_5833# VDPWR a_11541_5723# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X580 a_4546_2153# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X581 VGND VDPWR a_11986_4959# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X582 a_4637_10577# VGND VDPWR w_4540_10763# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X583 VDPWR sky130_fd_sc_hd__mux4_1_0.A3 a_2217_5025# w_6074_6018# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X584 a_10569_1777# a_9629_2033# VDPWR w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X585 a_11623_4959# a_10639_4597# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X586 VDPWR VGND a_15978_5459# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X587 a_9717_13091# VGND VDPWR w_9394_13055# sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X588 a_9727_11277# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X589 a_7815_2035# a_6885_1783# a_8232_2145# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X590 a_7899_5039# a_6915_5043# VDPWR w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X591 VGND ui_in[0] a_23731_14309# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4368,272
X592 VDPWR a_14846_1739# a_14794_1765# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X593 a_6003_11935# a_4849_11293# VDPWR w_5906_12121# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X594 a_9557_5837# VDPWR a_9461_5837# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X595 VDPWR VDPWR a_6362_1783# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X596 a_12250_2139# VDPWR a_11499_2029# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X597 VDPWR VDPWR a_13732_1769# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X598 a_16486_16197# sky130_fd_sc_hd__mux4_1_0.A0 VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X599 VGND VDPWR a_4721_13809# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X600 a_9725_5471# a_9671_5727# a_9332_5445# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X601 VDPWR VDPWR a_9753_4597# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X602 a_11455_4593# VDPWR a_11359_4593# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X603 a_16167_5459# a_15227_5715# VDPWR w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X604 a_9877_10533# a_9599_10561# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X605 VGND a_11202_5441# a_11150_5467# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X606 a_14975_1765# VGND VDPWR w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X607 a_14888_5433# a_14297_5463# a_15113_5459# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X608 VGND a_12075_13379# a_12631_13987# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2268,138 d=4075,198
X609 VDPWR a_9801_12841# a_10937_12911# w_10872_13125# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0805 ps=0.94333 w=0.42 l=0.15
**devattr s=2646,147 d=5689,267
X610 VDPWR VDPWR a_11958_5467# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X611 a_2343_5051# a_2217_5025# VDPWR w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X612 VGND VGND a_13369_2135# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X613 VGND VDPWR a_13802_4955# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X614 a_7173_15235# a_6635_15235# VDPWR w_6570_15449# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X615 a_24234_14385# a_24774_14701# a_24962_14701# sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1274 pd=1.16667 as=0.09209 ps=0.99 w=0.42 l=0.15
**devattr s=3683,198 d=10752,424
X616 a_6726_5409# VDPWR a_5975_5299# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X617 VDPWR VDPWR a_6029_5043# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X618 a_2313_1791# a_2259_2047# a_1920_1765# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X619 a_12881_13987# a_12135_15219# a_12809_13987# w_12566_13951# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X620 a_4576_5413# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X621 a_4755_12857# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X622 VGND a_4515_11543# a_4849_11293# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X623 VDPWR a_7506_5013# a_7454_5039# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X624 a_9515_1777# VDPWR a_9419_1777# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X625 VGND a_12976_1743# a_12924_1769# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X626 a_13201_2135# VDPWR a_13105_2135# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X627 a_15185_2021# a_14255_1769# a_15602_2131# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X628 VGND VGND a_12292_5833# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X629 a_10088_5471# VGND VDPWR w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X630 a_4585_16339# VDPWR a_4503_16339# w_4430_16303# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X631 VGND a_9477_11527# a_9811_11277# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X632 VDPWR a_14946_4905# a_16006_4585# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X633 VDPWR a_4839_12857# a_5809_14763# w_5712_14949# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X634 a_7635_5039# VGND VDPWR w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X635 VGND VGND a_9465_16323# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X636 a_4595_14775# VDPWR a_4513_14775# w_4440_14739# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X637 VGND VGND a_12250_2139# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X638 VDPWR a_9360_4571# a_9308_4597# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X639 a_15309_4951# a_15255_4841# a_14916_4559# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X640 a_9585_4963# VDPWR a_9489_4963# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X641 VDPWR VGND a_7899_5039# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X642 a_15978_5825# VDPWR a_15227_5715# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X643 a_3790_1761# a_3199_1791# a_4015_2153# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X644 a_11958_5833# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X645 a_4015_1787# VDPWR a_3919_1787# w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X646 a_16195_4585# a_15255_4841# VDPWR w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X647 VGND VDPWR a_8232_2145# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X648 a_2049_1791# VGND VDPWR w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X649 a_2145_2157# VDPWR a_2049_2157# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X650 a_14916_4559# a_14325_4589# a_15141_4585# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X651 sky130_fd_sc_hd__mux4_1_0.A1 a_12631_13987# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4075,198 d=7020,368
X652 a_11351_13753# a_10813_13753# VDPWR w_10748_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X653 a_11916_2139# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X654 a_13271_4589# VDPWR a_13175_4589# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X655 a_6389_13769# a_5851_13769# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X656 a_4839_12857# a_4505_13107# a_4755_13107# w_4432_13071# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X657 VGND VGND a_6726_5409# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X658 VGND VDPWR a_4183_2153# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X659 VGND VDPWR a_11553_2139# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X660 a_19510_16177# a_18742_16187# VDPWR w_19322_16391# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X661 VGND a_4839_12857# a_6127_13769# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X662 VGND a_11351_13753# a_11824_13629# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4010,197
X663 a_3010_1791# VDPWR a_2259_2047# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X664 a_13369_1769# a_12439_1773# VDPWR w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X665 a_23511_14335# ui_in[0] ui_in[1] sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.09322 ps=1.07 w=0.42 l=0.15
**devattr s=3409,185 d=4368,272
X666 a_9725_14759# VGND VDPWR w_9402_14723# sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X667 a_4765_11293# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X668 VDPWR VGND a_6029_5043# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X669 a_5999_1783# a_5945_2039# a_5606_1757# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X670 VDPWR VGND a_15281_5459# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X671 a_21506_16181# a_20384_16179# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X672 VDPWR VDPWR a_9597_13793# w_9500_13979# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X673 a_4903_15345# a_4625_15373# VDPWR w_4528_15559# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X674 a_9629_2033# a_8755_1779# a_10046_2143# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X675 VGND a_9799_16073# a_11873_15219# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X676 a_9465_16323# VDPWR VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X677 a_14066_2135# VDPWR a_13315_2025# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X678 a_9799_16073# VDPWR a_9715_16073# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X679 VGND VDPWR a_8262_5405# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X680 a_11595_5467# a_11541_5723# a_11202_5441# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X681 VGND a_13018_5437# a_12966_5463# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X682 VGND VDPWR a_15602_2131# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X683 a_2343_5051# a_2289_5307# a_1950_5025# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X684 a_7669_14003# a_4915_10549# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4368,272 d=2772,150
X685 a_15071_1765# VDPWR a_14975_1765# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X686 a_9683_2143# a_8755_1779# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X687 a_16006_4951# VDPWR a_15255_4841# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X688 VDPWR a_6389_13769# a_6944_13645# w_6756_13609# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5830,267
X689 VDPWR a_8785_5039# a_16871_4938# w_16764_4814# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.1176 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2772,150
X690 a_13411_5463# a_12481_5467# VDPWR w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X691 a_13357_5719# a_12481_5467# a_13774_5829# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X692 VDPWR VGND a_9549_13091# w_9394_13055# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X693 VGND VDPWR a_9675_12125# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X694 VGND VGND a_9477_11527# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X695 a_24407_14651# a_23731_14309# a_24234_14385# sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09013 pd=0.995 as=0.1274 ps=1.16667 w=0.42 l=0.15
**devattr s=2268,138 d=3605,199
X696 VGND a_4839_12857# a_6129_12927# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5266,228
X697 a_2676_2157# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X698 a_11679_15219# a_8113_13753# a_11597_15219# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
X699 VGND VDPWR a_9685_10561# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X700 a_4213_5413# a_4159_5303# a_3820_5021# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X701 a_9699_4853# VDPWR a_10116_4597# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X702 a_15141_4951# VDPWR a_15045_4951# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X703 a_9587_15357# VGND VDPWR w_9490_15543# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X704 a_11019_12911# a_9811_11277# a_10937_12911# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=1764,126
X705 a_11243_11891# a_10965_11919# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X706 VGND VDPWR a_11916_2139# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X707 a_14136_4589# VDPWR a_13385_4845# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X708 a_4159_5303# a_3229_5051# a_4576_5047# w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X709 VDPWR VDPWR a_15672_4585# w_14764_4500# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X710 VGND a_8785_5039# a_17346_5265# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=4514,209
X711 VGND VGND a_4183_2153# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X712 a_8596_5039# VDPWR a_7845_5295# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X713 VGND a_9290_1751# a_9238_1777# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X714 a_9875_13765# a_9597_13793# VDPWR w_9500_13979# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X715 a_18742_16187# a_18128_16189# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X716 a_7869_2145# a_6885_1783# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X717 a_8113_13753# a_7669_14003# VDPWR w_7604_13967# sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5930,268 d=10800,508
X718 a_6329_12927# a_5975_12927# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=5266,228 d=6760,364
X719 sky130_fd_sc_hd__mux4_1_0.A2 a_15185_2021# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X720 VDPWR VGND a_15936_1765# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X721 VGND VGND a_14066_2135# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X722 a_9725_5837# a_9671_5727# a_9332_5445# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X723 a_5945_2039# a_5069_1787# a_6362_1783# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X724 a_11455_4959# VDPWR a_11359_4959# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X725 sky130_fd_sc_hd__mux4_1_0.A0 a_22274_16171# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X726 a_10965_11919# a_9811_11277# VDPWR w_10868_12105# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X727 a_24318_14385# sky130_fd_sc_hd__mux4_1_0.A2 VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.10858 pd=1.36 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X728 a_11623_4593# a_11569_4849# a_11230_4567# w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X729 a_9801_12841# VDPWR a_9717_12841# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X730 VDPWR VDPWR a_4627_12141# w_4530_12327# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X731 a_6281_11907# a_6003_11935# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X732 a_10380_1777# VDPWR a_9629_2033# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X733 VGND VDPWR a_10046_2143# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X734 a_4915_10549# a_4637_10577# VDPWR w_4540_10763# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X735 a_2343_5417# a_2217_5025# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X736 a_9290_1751# a_8755_1779# a_9515_1777# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X737 a_12976_1743# a_12439_1773# a_13201_2135# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X738 a_5831_1783# VDPWR a_5735_1783# w_5454_1698# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X739 a_24318_14385# a_23731_14309# a_24234_14385# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.10858 pd=1.36 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=4318,272
X740 a_9549_13091# VDPWR a_9467_13091# w_9394_13055# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X741 a_9477_11527# VDPWR VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X742 a_3229_5051# a_2289_5307# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X743 a_6087_14735# a_5809_14763# VDPWR w_5712_14949# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X744 VDPWR VDPWR a_4637_10577# w_4540_10763# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X745 VGND VDPWR a_6029_5409# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X746 a_12481_5467# a_11541_5723# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X747 a_11499_2029# a_10569_1777# a_11916_1773# w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X748 a_13369_1769# a_13315_2025# a_12976_1743# w_12824_1684# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X749 a_11427_5467# VDPWR a_11331_5467# w_11050_5382# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X750 VGND VDPWR a_13369_2135# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X751 a_4753_16339# VGND VDPWR w_4430_16303# sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X752 a_2175_5051# VDPWR a_2079_5051# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X753 a_10450_4963# VDPWR a_9699_4853# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X754 VDPWR VDPWR a_9683_1777# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X755 a_4763_14775# VGND VDPWR w_4440_14739# sky130_fd_pr__pfet_01v8_hvt ad=0.17667 pd=1.68667 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X756 a_9360_4571# VDPWR a_9585_4963# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X757 a_18128_16189# a_17254_16187# VDPWR w_17940_16403# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X758 a_4910_5413# VDPWR a_4159_5303# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X759 a_13439_4955# a_13385_4845# a_13046_4563# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X760 VDPWR VGND a_8596_5039# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X761 a_10088_5837# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X762 a_15017_5825# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X763 a_7899_5405# a_7845_5295# a_7506_5013# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X764 a_10422_5471# VDPWR a_9671_5727# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X765 VGND VDPWR a_6362_2149# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X766 VDPWR VDPWR a_10116_4597# w_9208_4512# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X767 a_13046_4563# a_12509_4593# a_13271_4589# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X768 a_9332_5445# VGND a_9557_5471# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X769 a_9599_10561# VGND VDPWR w_9502_10747# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X770 a_11359_4593# VGND VDPWR w_11078_4508# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X771 a_8785_5039# a_7845_5295# VDPWR w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X772 VGND a_3820_5021# a_3768_5047# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=4094,199
X773 a_11595_5833# a_10611_5471# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X774 VDPWR VDPWR a_7869_1779# w_7324_1694# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X775 VDPWR VDPWR a_13439_4589# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X776 a_7506_5013# a_6915_5043# a_7731_5039# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X777 VGND VDPWR a_15281_5825# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X778 VGND VGND a_7869_2145# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X779 a_9717_12841# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X780 a_8262_5039# VGND VDPWR w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X781 VDPWR VGND a_9557_14759# w_9402_14723# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X782 a_9867_12097# a_9589_12125# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X783 VDPWR VDPWR a_9725_5471# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X784 VDPWR VGND a_10380_1777# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X785 a_4839_12857# VDPWR a_4755_12857# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X786 a_3199_1791# a_2259_2047# VDPWR w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X787 a_12439_1773# a_11499_2029# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X788 a_9799_16073# a_9465_16323# a_9715_16323# w_9392_16287# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X789 a_12809_13987# a_11243_11891# a_12713_13987# w_12566_13951# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X790 a_2313_2157# a_2259_2047# a_1920_1765# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X791 VDPWR ui_in[0] a_23731_14309# sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.1083 ps=1.36 w=0.42 l=0.15
**devattr s=4332,272 d=4316,272
X792 a_1920_1765# a_2187_1765# a_2145_1791# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X793 VDPWR VGND a_4585_16339# w_4430_16303# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X794 a_17053_4938# a_16871_4938# VDPWR w_16764_4814# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X795 a_12075_13379# a_11824_13629# VDPWR w_11718_13593# sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5830,267 d=13600,536
X796 VDPWR VGND a_4595_14775# w_4440_14739# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X797 a_7701_2145# VDPWR a_7605_2145# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X798 VGND VGND a_10450_4963# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X799 a_15281_5825# a_15227_5715# a_14888_5433# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X800 a_10046_1777# VGND VDPWR w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X801 a_9419_1777# VGND VDPWR w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X802 VDPWR VDPWR a_2313_1791# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X803 a_13105_2135# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X804 VGND VGND a_4910_5413# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=4094,199
X805 a_2706_5051# VGND VDPWR w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X806 a_15227_5715# a_14297_5463# a_15644_5459# w_14736_5374# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X807 a_17254_16187# a_16486_16197# VDPWR w_17066_16401# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X808 VGND VGND a_6029_5409# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X809 a_14846_1739# a_14255_1769# a_15071_1765# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=2772,150
X810 a_6635_15235# a_6087_14735# VDPWR w_6570_15449# sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X811 a_5975_5299# a_5099_5047# a_6392_5043# w_5484_4958# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X812 a_11553_1773# a_10569_1777# VDPWR w_11008_1688# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X813 ui_in[1] a_23731_14309# a_23511_14701# sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0742 pd=0.91333 as=0.1092 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X814 VDPWR VGND a_10422_5471# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2520,144 d=5914,269
X815 VDPWR VGND a_9683_1777# w_9138_1692# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X816 VDPWR VDPWR a_15239_1765# w_14694_1680# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X817 a_10116_4963# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0742 pd=0.91333 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X818 a_9489_4963# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X819 a_13385_4845# a_12509_4593# a_13802_4955# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X820 a_24962_14701# ui_in[1] ui_in[1] sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09209 pd=0.99 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=3683,198
X821 a_3919_1787# VGND VDPWR w_3638_1702# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X822 VDPWR a_13046_4563# a_12994_4589# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X823 VGND a_7113_13395# a_7669_14003# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.063 ps=0.72 w=0.42 l=0.15
**devattr s=2268,138 d=4075,198
X824 VGND a_9467_13091# a_9801_12841# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.25025 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X825 a_10611_5471# a_9671_5727# VDPWR w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.20702 ps=2.00005 w=1 l=0.15
**devattr s=5914,269 d=10400,504
X826 a_2049_2157# VGND VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=4094,199 d=2772,150
X827 a_9557_14759# VDPWR a_9475_14759# w_9402_14723# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X828 a_2343_5417# a_2289_5307# a_1950_5025# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X829 a_7845_5295# a_6915_5043# a_8262_5405# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X830 VDPWR a_9332_5445# a_9280_5471# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X831 VGND sky130_fd_sc_hd__mux4_1_0.A2 a_2187_1765# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.12891 pd=1.32823 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X832 a_14946_4905# VDPWR a_15309_4951# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.07384 pd=0.80236 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X833 VGND VGND a_9753_4963# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X834 VDPWR VDPWR a_9725_14759# w_9402_14723# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X835 a_13175_4589# VGND VDPWR w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X836 a_4849_11293# VDPWR a_4765_11293# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X837 a_13411_5829# a_12481_5467# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0833 ps=0.85824 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X838 a_7731_5405# VDPWR a_7635_5405# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X839 a_14297_5463# a_13357_5719# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X840 VDPWR VGND a_13439_4589# w_12894_4504# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X841 a_9461_5471# VGND VDPWR w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=5914,269 d=2772,150
X842 a_15239_2131# a_15185_2021# a_14846_1739# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X843 a_3010_2157# VDPWR a_2259_2047# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X844 a_7173_15235# a_6635_15235# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X845 a_13243_5463# VDPWR a_13147_5463# w_12866_5378# sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=1764,126
X846 a_5851_13769# a_4837_16089# VDPWR w_5786_13983# sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X847 a_4849_11293# a_4515_11543# a_4765_11543# w_4442_11507# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X848 VDPWR VGND a_9725_5471# w_9180_5386# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2478,143 d=2268,138
X849 a_14255_1769# a_13315_2025# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=4094,199 d=6760,364
X850 VGND a_4905_12113# a_6089_11935# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0833 pd=0.85824 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X851 a_4213_5047# a_3229_5051# VDPWR w_3668_4962# sky130_fd_pr__pfet_01v8_hvt ad=0.05932 pd=0.7025 as=0.08695 ps=0.84002 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X852 a_5999_2149# a_5945_2039# a_5606_1757# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.05932 pd=0.7025 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=2478,143
X853 a_4129_2043# a_3199_1791# a_4546_2153# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=2268,138 d=2268,138
X854 a_9811_11277# a_9477_11527# a_9727_11527# w_9404_11491# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.17667 ps=1.68667 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X855 a_20384_16179# a_19510_16177# VGND sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12891 ps=1.32823 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X856 a_6911_15235# a_6087_14735# a_6805_15235# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X857 VDPWR a_4839_12857# a_5851_13769# w_5786_13983# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.06615 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X858 VDPWR a_1950_5025# a_1898_5051# w_1798_4966# sky130_fd_pr__pfet_01v8_hvt ad=0.20702 pd=2.00005 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5914,269
X859 a_8566_2145# VDPWR a_7815_2035# sky130_fd_sc_hd__mux4_1_0.VNB sky130_fd_pr__nfet_01v8 ad=0.063 pd=0.72 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=2520,144
X860 VDPWR VDPWR a_2676_1791# w_1768_1706# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.0742 ps=0.91333 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X861 VDPWR VDPWR a_7899_5039# w_7354_4954# sky130_fd_pr__pfet_01v8_hvt ad=0.08695 pd=0.84002 as=0.05932 ps=0.7025 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
C0 a_12976_1743# a_12924_1769# 0.1439f
C1 a_15936_2131# sky130_fd_sc_hd__mux4_1_0.A2 0
C2 a_14946_4905# a_14325_4589# 0.58451f
C3 a_5975_5299# a_6029_5409# 0.03622f
C4 a_12509_4593# a_8785_5039# 0.02903f
C5 w_1768_1706# ua[7] 0
C6 ui_in[0] sky130_fd_sc_hd__mux4_1_0.VPB 0.35114f
C7 a_7899_5039# VGND 0.0165f
C8 a_9683_13793# a_9875_13765# 0.00222f
C9 VDPWR a_4587_13107# 0.02512f
C10 sky130_fd_sc_hd__mux4_1_0.A3 a_10611_5471# 0.0073f
C11 a_14794_1765# VGND 0.08635f
C12 w_5786_13983# a_4849_11293# 0.10705f
C13 a_4045_5047# VGND 0
C14 a_13385_4845# w_12866_5378# 0.00166f
C15 VGND a_5099_5047# 0.67875f
C16 a_15141_4951# a_15309_4951# 0
C17 a_10937_12911# w_10872_13125# 0.04996f
C18 a_9589_12125# w_9502_10747# 0
C19 a_3820_5021# w_3668_4962# 0.05213f
C20 a_4903_15345# a_6389_13769# 0
C21 a_5945_2039# VGND 1.20001f
C22 a_12250_2139# a_12439_1773# 0
C23 a_9360_4571# sky130_fd_sc_hd__mux4_1_0.A3 0
C24 a_9727_11277# VGND 0.00834f
C25 a_9629_2033# VGND 1.19975f
C26 w_11532_15433# a_12135_15219# 0.01567f
C27 a_6362_2149# w_5454_1698# 0.00139f
C28 a_10569_1777# w_11008_1688# 0.25055f
C29 a_4753_16339# a_6629_15387# 0
C30 a_6003_11935# a_4849_11293# 0.10332f
C31 ui_in[0] rst_n 0.03102f
C32 a_14916_4559# a_14297_5463# 0
C33 a_21506_16181# a_22274_16171# 0.1036f
C34 a_14836_5459# VDPWR 0.07614f
C35 w_9180_5386# a_8785_5039# 0.00671f
C36 VGND a_6389_13769# 0.25955f
C37 a_7701_1779# a_7869_1779# 0
C38 VGND a_4576_5047# 0.01333f
C39 a_11289_1773# a_11160_1747# 0.00758f
C40 a_4903_15345# a_4849_11293# 0.30844f
C41 uio_oe[4] uio_oe[3] 0.03102f
C42 a_15936_2131# VGND 0.00236f
C43 w_22086_16385# VDPWR 0.07223f
C44 ui_in[0] a_24318_14385# 0.00255f
C45 a_9801_12841# a_11091_12911# 0.00312f
C46 w_5786_13983# a_7669_14003# 0
C47 a_4763_14775# a_4513_14775# 0.02504f
C48 w_11078_4508# a_11178_4593# 0.01793f
C49 a_15602_2131# a_14255_1769# 0.03325f
C50 w_4530_12327# VDPWR 0.17848f
C51 a_13201_2135# a_13315_2025# 0
C52 a_4847_14525# w_6570_15449# 0.07233f
C53 a_9877_10533# a_9685_10561# 0
C54 w_9392_17212# VGND 0.01278f
C55 a_9599_10561# VDPWR 0.36832f
C56 a_7605_1779# a_7476_1753# 0.00758f
C57 VGND a_4849_11293# 1.26863f
C58 a_9673_15357# VGND 0.00661f
C59 a_6089_11935# a_4915_10549# 0
C60 a_10569_1777# a_11385_1773# 0
C61 w_7604_13967# a_7173_15235# 0.11864f
C62 a_5945_2039# a_5999_1783# 0.00386f
C63 VDPWR a_11906_13629# 0.0014f
C64 VDPWR a_11958_5833# 0.01821f
C65 a_4637_10577# a_4849_11293# 0
C66 a_14325_4589# VDPWR 1.12038f
C67 a_7845_5295# a_9308_4597# 0
C68 a_8596_5405# a_8785_5039# 0
C69 w_4430_16303# a_4513_14775# 0
C70 VGND a_9867_12097# 0.43935f
C71 a_12976_1743# a_13201_2135# 0.00559f
C72 a_6629_15387# w_5712_14949# 0
C73 VGND a_7669_14003# 0.24155f
C74 VDPWR a_10422_5471# 0
C75 a_8755_1779# a_9290_1751# 0.11411f
C76 a_5809_14763# a_7173_15235# 0
C77 a_2217_5025# a_6029_5043# 0
C78 VGND w_17066_16401# 0.01227f
C79 a_12631_13987# w_11718_13593# 0
C80 VDPWR a_5831_2149# 0
C81 a_14836_5459# a_15017_5825# 0
C82 a_5851_13769# a_6389_13769# 0.07901f
C83 sky130_fd_sc_hd__mux4_1_0.A3 a_11427_5467# 0
C84 a_15255_4841# a_16167_5459# 0
C85 a_4839_12857# a_6129_12927# 0.00312f
C86 a_9587_15357# w_9500_13979# 0
C87 VDPWR a_4515_11543# 0.3853f
C88 a_9683_1777# a_8755_1779# 0.08124f
C89 VDPWR a_9308_4597# 0.10729f
C90 a_14946_4905# a_15978_5459# 0
C91 a_5851_13769# a_4849_11293# 0.17627f
C92 a_9809_14509# a_9465_16323# 0
C93 a_9877_10533# a_12135_15219# 0.07807f
C94 VGND a_19510_16177# 0.26921f
C95 a_9811_11277# a_11019_12911# 0.00146f
C96 a_7113_13395# w_6756_13609# 0.03222f
C97 a_2343_5417# a_2079_5417# 0
C98 a_12631_13987# a_12809_13987# 0.00412f
C99 a_4837_16089# a_4913_13781# 0.01745f
C100 w_9394_13055# a_9801_12841# 0.02723f
C101 a_23511_14335# ui_in[1] 0.08552f
C102 a_13271_4955# VGND 0.00234f
C103 a_6805_15235# a_4847_14525# 0.00624f
C104 a_4763_14775# a_4503_16339# 0
C105 a_15255_4841# a_15309_4585# 0.00386f
C106 a_9629_2033# a_10046_2143# 0.06611f
C107 w_9138_1692# sky130_fd_sc_hd__mux4_1_0.A2 0.00331f
C108 a_9727_11527# a_9811_11277# 0.08177f
C109 sky130_fd_sc_hd__mux4_1_0.A2 sky130_fd_sc_hd__mux4_1_0.A3 0.91673f
C110 w_11078_4508# a_10639_4597# 0.25055f
C111 a_4849_11293# a_6057_12927# 0.00146f
C112 a_5851_13769# a_7669_14003# 0
C113 a_10965_11919# a_11243_11891# 0.11706f
C114 a_4837_16089# a_6717_15235# 0
C115 w_20196_16393# VGND 0.01236f
C116 a_5554_1783# a_2187_1765# 0.0012f
C117 a_2706_5417# VGND 0.18671f
C118 VGND a_15227_5715# 1.19394f
C119 a_4183_2153# VDPWR 0.00888f
C120 a_14946_4905# a_13802_4589# 0
C121 a_4503_16339# w_4430_16303# 0.06993f
C122 VDPWR a_11385_2139# 0
C123 a_21506_16181# sky130_fd_sc_hd__mux4_1_0.A0 0.04638f
C124 a_4159_5303# a_2217_5025# 0.00305f
C125 a_15978_5825# a_16167_5459# 0
C126 a_9671_5727# a_7845_5295# 0
C127 w_14764_4500# sky130_fd_sc_hd__mux4_1_0.A2 0.00111f
C128 VGND w_9138_1692# 0.2932f
C129 a_13046_4563# sky130_fd_sc_hd__mux4_1_0.A2 0
C130 a_9465_16323# VGND 0.28565f
C131 VDPWR a_11331_5467# 0.00136f
C132 VGND sky130_fd_sc_hd__mux4_1_0.A3 2.34296f
C133 a_7815_2035# a_7869_1779# 0.00386f
C134 a_5809_14763# a_4513_14775# 0
C135 a_7869_2145# a_7476_1753# 0.02301f
C136 a_9801_12841# a_9477_11527# 0
C137 a_11359_4959# VGND 0.00292f
C138 a_7113_13395# a_8113_13753# 0.02955f
C139 uio_oe[1] uio_oe[2] 0.03102f
C140 a_10937_12911# a_9875_13765# 0.08477f
C141 w_12866_5378# a_13411_5829# 0
C142 a_9865_15329# a_9587_15357# 0.12165f
C143 VGND w_4432_13071# 0.07276f
C144 a_21506_16181# a_20384_16179# 0.10186f
C145 VDPWR a_11553_1773# 0.17705f
C146 a_15978_5459# VDPWR 0
C147 a_8755_1779# a_9515_1777# 0
C148 a_11427_5467# a_10611_5471# 0
C149 a_6329_12927# a_7113_13395# 0
C150 a_2217_5025# a_3949_5047# 0
C151 a_6885_1783# a_8232_2145# 0.03325f
C152 a_9332_5445# a_9308_4597# 0
C153 a_9465_16323# a_9715_16323# 0.02504f
C154 w_1768_1706# a_3790_1761# 0
C155 a_9671_5727# VDPWR 0.35696f
C156 w_4430_16303# a_4753_16339# 0.01327f
C157 a_13201_1769# a_13315_2025# 0
C158 VDPWR a_15045_4585# 0.00135f
C159 VGND w_14764_4500# 0.00461f
C160 a_17254_16187# a_16486_16197# 0.1036f
C161 ui_in[1] sky130_fd_sc_hd__mux4_1_0.VPB 0.27196f
C162 VGND a_13046_4563# 0.41147f
C163 a_7424_1779# w_7324_1694# 0.01793f
C164 a_4837_16089# a_4585_16339# 0
C165 a_3949_5413# VGND 0.00305f
C166 a_11150_5467# a_11331_5833# 0
C167 a_2145_1791# a_2313_1791# 0
C168 a_9477_11527# w_9492_12311# 0
C169 a_11499_2029# VDPWR 0.3456f
C170 w_10868_12105# a_10937_12911# 0
C171 a_4837_16089# a_5895_14763# 0
C172 a_7899_5405# w_7354_4954# 0
C173 a_8232_1779# sky130_fd_sc_hd__mux4_1_0.A2 0
C174 a_9360_4571# sky130_fd_sc_hd__mux4_1_0.A2 0
C175 a_2343_5051# VDPWR 0.17446f
C176 VDPWR a_13802_4589# 0.2102f
C177 a_12976_1743# a_13201_1769# 0.00487f
C178 a_23677_14335# VGND 0.00194f
C179 a_14255_1769# a_15185_2021# 0.21188f
C180 a_15672_4951# a_14325_4589# 0.03325f
C181 a_4880_2153# a_5069_1787# 0
C182 a_7731_5405# a_7845_5295# 0
C183 w_9394_13055# a_9475_14759# 0
C184 a_7815_2035# a_8566_2145# 0.00696f
C185 a_24318_14385# ui_in[1] 0.04767f
C186 a_10569_1777# a_11108_1773# 0.0725f
C187 a_5554_1783# a_5606_1757# 0.1439f
C188 a_2343_5051# a_1950_5025# 0.02283f
C189 a_4045_5413# a_2217_5025# 0
C190 a_14836_5459# a_13357_5719# 0
C191 w_12894_4504# sky130_fd_sc_hd__mux4_1_0.A3 0
C192 a_2217_5025# a_5584_5043# 0.0012f
C193 a_13018_5437# a_12966_5463# 0.1439f
C194 a_1868_1791# a_2049_2157# 0
C195 a_15227_5715# a_8785_5039# 0
C196 a_9599_10561# a_4915_10549# 0
C197 a_11230_4567# a_11202_5441# 0
C198 VGND a_10611_5471# 0.69145f
C199 a_3040_5051# a_2289_5307# 0.00682f
C200 a_5975_5299# a_7454_5039# 0
C201 ui_in[4] ui_in[5] 0.03102f
C202 a_4913_13781# a_6389_13769# 0
C203 a_8232_1779# VGND 0.01329f
C204 a_9360_4571# VGND 0.41248f
C205 w_14736_5374# a_15281_5459# 0.01092f
C206 VGND a_11243_11891# 0.5959f
C207 a_7731_5405# VDPWR 0
C208 a_1898_5051# VGND 0.09486f
C209 w_9138_1692# a_10046_2143# 0.00139f
C210 a_11291_12911# a_11351_13753# 0.20048f
C211 sky130_fd_sc_hd__mux4_1_0.A3 a_8785_5039# 0.02419f
C212 a_9671_5727# a_9332_5445# 0.04737f
C213 a_4913_13781# a_4849_11293# 0.26616f
C214 a_13046_4563# w_12894_4504# 0.05213f
C215 VDPWR a_13175_4589# 0.00117f
C216 a_9753_4597# a_10116_4597# 0.00985f
C217 VGND a_10965_11919# 0.13487f
C218 a_9725_14759# w_9402_14723# 0.01327f
C219 a_7845_5295# a_7506_5013# 0.04737f
C220 w_11718_13593# a_12135_15219# 0
C221 VGND a_3010_2157# 0.00245f
C222 a_14946_4905# a_15281_5459# 0.00242f
C223 a_11597_15219# a_12135_15219# 0.08446f
C224 a_14916_4559# a_15227_5715# 0
C225 w_14764_4500# a_8785_5039# 0.0011f
C226 a_4763_14775# a_4839_12857# 0.00187f
C227 a_4515_11543# a_4915_10549# 0
C228 a_13046_4563# a_8785_5039# 0
C229 a_10450_4597# VDPWR 0
C230 a_10046_1777# a_9683_1777# 0.00985f
C231 a_13774_5463# a_13411_5463# 0.00985f
C232 w_10748_13967# a_9865_15329# 0.07513f
C233 w_4440_14739# a_4847_14525# 0.02435f
C234 a_14916_4559# sky130_fd_sc_hd__mux4_1_0.A3 0
C235 VDPWR a_7506_5013# 0.29452f
C236 VDPWR w_11008_1688# 0.5148f
C237 a_11499_2029# a_12439_1773# 0.1382f
C238 w_10748_13967# a_11351_13753# 0.01492f
C239 a_5861_5043# VDPWR 0
C240 VGND a_11427_5467# 0
C241 a_5809_14763# w_5712_14949# 0.05631f
C242 a_9809_14509# a_11767_15219# 0.00624f
C243 sky130_fd_sc_hd__mux4_1_0.A3 a_17346_5265# 0.00101f
C244 a_24152_14385# a_24774_14701# 0
C245 sky130_fd_sc_hd__mux4_1_0.A3 a_23677_14701# 0
C246 a_4159_5303# a_3820_5021# 0.04737f
C247 a_9597_13793# w_9402_14723# 0
C248 a_14916_4559# w_14764_4500# 0.05213f
C249 VDPWR a_11385_1773# 0
C250 a_4635_13809# w_4440_14739# 0
C251 a_12481_5467# a_14297_5463# 0
C252 VDPWR a_9419_1777# 0.00114f
C253 a_3229_5051# a_2217_5025# 0.00475f
C254 VGND a_2175_5051# 0
C255 a_9809_14509# VGND 0.43095f
C256 w_5786_13983# a_4903_15345# 0.07513f
C257 a_8785_5039# a_10611_5471# 0.04731f
C258 a_17254_16187# w_18554_16401# 0
C259 a_23511_14335# a_23511_14701# 0.00987f
C260 a_11499_2029# a_12250_2139# 0.00696f
C261 a_15281_5459# VDPWR 0.16927f
C262 a_5636_5017# w_3668_4962# 0
C263 a_9877_10533# w_10868_12105# 0
C264 a_9360_4571# a_8785_5039# 0
C265 a_9801_12841# a_11291_12911# 0.08252f
C266 a_15255_4841# w_16764_4814# 0.00175f
C267 a_9290_1751# a_9238_1777# 0.1439f
C268 a_3820_5021# a_3949_5047# 0.00758f
C269 w_5786_13983# VGND 0.01862f
C270 a_12481_5467# a_12509_4593# 0.00249f
C271 a_10639_4597# a_10116_4597# 0
C272 VDPWR w_4528_15559# 0.18191f
C273 VGND sky130_fd_sc_hd__mux4_1_0.A2 0.75219f
C274 w_5484_4958# a_7506_5013# 0
C275 a_10813_13753# a_11089_13753# 0.00119f
C276 a_14946_4905# a_14136_4955# 0
C277 w_4530_12327# a_4515_11543# 0
C278 VDPWR a_10380_1777# 0
C279 VGND a_6003_11935# 0.13487f
C280 a_14846_1739# a_15071_1765# 0.00487f
C281 a_12631_13987# a_11243_11891# 0.19153f
C282 a_9597_13793# a_9875_13765# 0.1205f
C283 a_5895_14763# a_4849_11293# 0.00121f
C284 a_4755_12857# a_4505_13107# 0.00723f
C285 a_4837_16089# a_7173_15235# 0.04819f
C286 a_15602_1765# a_15185_2021# 0.03016f
C287 a_6915_5043# a_7506_5013# 0.11887f
C288 a_14136_4589# sky130_fd_sc_hd__mux4_1_0.A2 0
C289 VGND a_11767_15219# 0.00334f
C290 VGND a_4903_15345# 0.98587f
C291 a_9332_5445# a_7506_5013# 0
C292 a_4213_5047# a_4045_5047# 0
C293 a_4913_13781# w_4432_13071# 0.00226f
C294 a_4576_5413# VDPWR 0.01963f
C295 w_7604_13967# a_4839_12857# 0
C296 a_9475_14759# a_9587_15357# 0
C297 sky130_fd_sc_hd__mux4_1_0.A1 a_8113_13753# 0.16034f
C298 a_9727_11527# a_9467_13091# 0
C299 a_16195_4585# a_15309_4951# 0
C300 a_7635_5039# VDPWR 0.00116f
C301 w_14736_5374# a_15281_5825# 0
C302 a_4213_5047# a_4576_5047# 0.00985f
C303 w_10748_13967# a_9801_12841# 0.08124f
C304 a_5999_1783# sky130_fd_sc_hd__mux4_1_0.A2 0
C305 a_14297_5463# a_15017_5459# 0
C306 a_12439_1773# w_11008_1688# 0.0197f
C307 a_9717_13091# VGND 0.02544f
C308 a_4045_5413# a_3820_5021# 0.00559f
C309 a_11541_5723# sky130_fd_sc_hd__mux4_1_0.A3 0.00769f
C310 VDPWR w_6756_13609# 0.08767f
C311 a_5809_14763# a_4839_12857# 0.21988f
C312 a_5851_13769# w_5786_13983# 0.08205f
C313 a_14136_4589# VGND 0
C314 a_8755_1779# a_9683_2143# 0.04534f
C315 a_4637_10577# VGND 0.2439f
C316 VGND a_9715_16323# 0.01705f
C317 VDPWR a_9675_12125# 0.00297f
C318 a_5069_1787# w_5454_1698# 0.24988f
C319 a_6281_11907# w_7604_13967# 0.03664f
C320 a_6862_13645# w_6756_13609# 0.06114f
C321 a_14946_4905# a_15281_5825# 0.00186f
C322 a_16486_16197# w_17940_16403# 0
C323 a_23511_14701# sky130_fd_sc_hd__mux4_1_0.VPB 0.02285f
C324 VDPWR a_2343_5417# 0.00857f
C325 a_14136_4955# VDPWR 0
C326 a_5851_13769# a_4903_15345# 0.16764f
C327 a_15239_2131# a_15071_2131# 0
C328 w_12894_4504# sky130_fd_sc_hd__mux4_1_0.A2 0.00104f
C329 w_10872_13125# a_9867_12097# 0
C330 w_1768_1706# a_2259_2047# 0.10454f
C331 a_18128_16189# a_16486_16197# 0
C332 a_11289_2139# sky130_fd_sc_hd__mux4_1_0.A2 0
C333 w_1768_1706# a_3199_1791# 0.02026f
C334 a_2343_5417# a_1950_5025# 0.02301f
C335 a_5999_1783# VGND 0.01528f
C336 a_7424_1779# w_5454_1698# 0.00188f
C337 a_5554_1783# VDPWR 0.07432f
C338 ui_in[7] ui_in[6] 0.03102f
C339 a_5851_13769# VGND 0.15513f
C340 a_4837_16089# a_4513_14775# 0
C341 a_9799_16073# a_8113_13753# 0.36356f
C342 a_11958_5467# a_11595_5467# 0.00985f
C343 sky130_fd_sc_hd__mux4_1_0.A2 a_10046_2143# 0
C344 VDPWR a_8113_13753# 2.11591f
C345 a_6915_5043# a_7635_5039# 0
C346 a_4847_14525# a_4625_15373# 0.00215f
C347 a_14066_2135# a_13315_2025# 0.00696f
C348 a_9753_4963# a_7845_5295# 0
C349 VGND w_12894_4504# 0.28722f
C350 a_9811_11277# a_9799_16073# 0.03118f
C351 a_17254_16187# sky130_fd_sc_hd__mux4_1_0.A0 0.05745f
C352 a_6329_12927# VDPWR 0.23898f
C353 a_11289_2139# VGND 0.00305f
C354 VGND a_10857_14747# 0.00618f
C355 VGND a_6057_12927# 0.00238f
C356 VDPWR a_14108_5463# 0
C357 a_14325_4589# a_15045_4585# 0
C358 a_13018_5437# a_13411_5829# 0.02301f
C359 VDPWR a_9811_11277# 0.42529f
C360 a_6329_12927# a_6862_13645# 0.10646f
C361 a_15936_1765# sky130_fd_sc_hd__mux4_1_0.A2 0
C362 a_9671_5727# a_10422_5471# 0.00682f
C363 w_22960_16387# a_22274_16171# 0.05645f
C364 a_9725_5471# a_9557_5471# 0
C365 VDPWR a_15281_5825# 0.00604f
C366 a_11541_5723# a_10611_5471# 0.21188f
C367 VGND a_8785_5039# 1.9195f
C368 a_15309_4951# a_14297_5463# 0
C369 VDPWR a_9753_4963# 0.05505f
C370 VGND a_10046_2143# 0.1864f
C371 a_4635_13809# a_4625_15373# 0
C372 a_14916_4559# sky130_fd_sc_hd__mux4_1_0.A2 0
C373 a_6629_15387# a_6087_14735# 0.09734f
C374 ua[4] a_14846_1739# 0
C375 a_5999_2149# w_5454_1698# 0
C376 a_6389_13769# a_7173_15235# 0.00152f
C377 a_12631_13987# VGND 0.24002f
C378 VDPWR a_6726_5043# 0
C379 a_4837_16089# w_5906_12121# 0
C380 VDPWR a_11108_1773# 0.07418f
C381 a_14325_4589# a_13802_4589# 0
C382 a_3229_5051# a_3820_5021# 0.11887f
C383 w_12866_5378# a_14888_5433# 0
C384 a_11986_4593# a_10639_4597# 0.08907f
C385 a_15936_1765# VGND 0
C386 a_9461_5837# a_9725_5837# 0
C387 a_4015_2153# a_2187_1765# 0
C388 a_4849_11293# a_7173_15235# 0
C389 a_4837_16089# a_4503_16339# 0.16891f
C390 a_11595_5833# sky130_fd_sc_hd__mux4_1_0.A3 0.00169f
C391 a_14916_4559# VGND 0
C392 a_13105_2135# sky130_fd_sc_hd__mux4_1_0.A2 0
C393 a_1920_1765# a_2259_2047# 0.04737f
C394 a_2313_1791# a_2187_1765# 0.08436f
C395 a_15017_5825# a_15281_5825# 0
C396 a_5945_2039# a_6885_1783# 0.13962f
C397 a_16195_4585# a_16167_5459# 0.39945f
C398 a_17125_4938# a_16167_5459# 0.06947f
C399 a_2217_5025# a_2079_5417# 0
C400 a_11824_13629# a_9799_16073# 0
C401 a_23731_14309# sky130_fd_sc_hd__mux4_1_0.A3 0.1036f
C402 a_7669_14003# a_7173_15235# 0.16709f
C403 a_4837_16089# a_4753_16339# 0.07445f
C404 VGND a_17346_5265# 0.00328f
C405 a_6635_15235# w_6756_13609# 0
C406 VGND a_23677_14701# 0.00402f
C407 a_13147_5463# sky130_fd_sc_hd__mux4_1_0.A3 0
C408 a_10813_13753# a_10937_12911# 0
C409 a_12135_15219# a_11243_11891# 0.09936f
C410 uio_out[3] uio_out[4] 0.03102f
C411 VDPWR a_11824_13629# 0.09661f
C412 a_11049_14719# w_11532_15433# 0.06196f
C413 w_12894_4504# a_8785_5039# 0.00112f
C414 a_11541_5723# a_11427_5467# 0
C415 a_24152_14385# a_24234_14385# 0.04662f
C416 a_11873_15219# a_9799_16073# 0.00241f
C417 a_13105_2135# VGND 0.00305f
C418 a_4913_13781# w_5786_13983# 0.00175f
C419 VDPWR a_11873_15219# 0
C420 a_11569_4849# a_10639_4597# 0.21188f
C421 a_9875_13765# a_9867_12097# 0.00627f
C422 a_4913_13781# a_6003_11935# 0
C423 a_11499_2029# a_11385_2139# 0
C424 a_9585_4963# sky130_fd_sc_hd__mux4_1_0.A3 0
C425 a_5636_5017# a_6029_5043# 0.02283f
C426 a_5945_2039# a_5831_1783# 0
C427 w_18554_16401# a_18128_16189# 0.05841f
C428 a_11569_4849# a_11595_5467# 0
C429 a_10813_13753# a_12075_13379# 0
C430 a_5975_5299# a_6029_5043# 0.00386f
C431 a_4913_13781# a_4903_15345# 0.1161f
C432 a_2049_2157# a_2187_1765# 0
C433 a_11499_2029# a_11553_1773# 0.00386f
C434 w_6756_13609# a_4915_10549# 0.00404f
C435 a_4849_11293# a_4513_14775# 0.00146f
C436 a_9675_12125# a_4915_10549# 0
C437 a_5861_5409# a_6029_5409# 0
C438 a_4913_13781# VGND 0.70497f
C439 a_12481_5467# sky130_fd_sc_hd__mux4_1_0.A3 0.00671f
C440 a_14916_4559# w_12894_4504# 0
C441 a_4837_16089# w_5712_14949# 0.00872f
C442 a_11595_5833# a_10611_5471# 0.04534f
C443 w_10872_13125# a_11243_11891# 0
C444 w_22960_16387# sky130_fd_sc_hd__mux4_1_0.A0 0.04283f
C445 a_4910_5047# VDPWR 0
C446 a_2175_5417# a_2289_5307# 0
C447 sky130_fd_sc_hd__mux4_1_0.A1 w_9490_15543# 0
C448 a_12966_5463# VDPWR 0.06838f
C449 a_9465_16323# w_9402_14723# 0
C450 w_22960_16387# a_20384_16179# 0
C451 w_10868_12105# a_9867_12097# 0.08119f
C452 a_18742_16187# w_19322_16391# 0.05681f
C453 a_14916_4559# a_8785_5039# 0
C454 a_10965_11919# w_10872_13125# 0
C455 VGND a_6717_15235# 0.00151f
C456 ui_in[0] a_24152_14385# 0.03464f
C457 a_5765_5409# a_6029_5409# 0
C458 VGND a_11541_5723# 1.23723f
C459 a_14325_4589# a_15281_5459# 0
C460 w_11078_4508# a_12994_4589# 0.00227f
C461 a_7815_2035# w_7324_1694# 0.10454f
C462 VDPWR a_4763_14525# 0.00474f
C463 a_9685_10561# VGND 0.00697f
C464 a_12481_5467# a_13046_4563# 0
C465 a_13243_5463# sky130_fd_sc_hd__mux4_1_0.A3 0
C466 a_24407_14651# a_24774_14701# 0
C467 a_9809_14509# a_12135_15219# 0
C468 a_10937_12911# a_10771_14747# 0
C469 a_14297_5463# a_16167_5459# 0
C470 a_14946_4905# a_13385_4845# 0.00318f
C471 a_14846_1739# a_15239_1765# 0.02283f
C472 a_8113_13753# a_4915_10549# 0.13594f
C473 a_5636_5017# a_4159_5303# 0.00492f
C474 a_9725_5837# VDPWR 0.00613f
C475 a_7869_1779# VDPWR 0.17565f
C476 a_5851_13769# a_4913_13781# 0.0094f
C477 w_5906_12121# a_4849_11293# 0.0984f
C478 a_13732_1769# a_14255_1769# 0
C479 a_1920_1765# a_2049_1791# 0.00758f
C480 a_16486_16197# w_17066_16401# 0.05681f
C481 a_14946_4905# a_15672_4585# 0.01208f
C482 a_9811_11277# a_4915_10549# 0
C483 a_9559_11527# VGND 0.00172f
C484 a_8262_5405# w_7354_4954# 0.00139f
C485 a_9799_16073# a_11679_15219# 0
C486 a_7899_5039# a_7731_5039# 0
C487 a_9360_4571# a_9585_4963# 0.00559f
C488 w_11078_4508# VDPWR 0.52719f
C489 sky130_fd_sc_hd__mux4_1_0.A3 a_15017_5459# 0
C490 a_14297_5463# a_15309_4585# 0
C491 VDPWR a_11679_15219# 0
C492 a_14108_5463# a_13357_5719# 0.00682f
C493 a_11289_1773# sky130_fd_sc_hd__mux4_1_0.A2 0
C494 a_11767_15219# a_12135_15219# 0
C495 a_9799_16073# w_9490_15543# 0.00251f
C496 a_11202_5441# w_11050_5382# 0.05213f
C497 a_12481_5467# a_10611_5471# 0
C498 a_9727_11527# a_9477_11527# 0.02504f
C499 a_2259_2047# a_2676_2157# 0.06611f
C500 w_11008_1688# a_11553_1773# 0.01092f
C501 a_4837_16089# a_4839_12857# 0.4639f
C502 a_4585_16339# VGND 0.00117f
C503 a_5895_14763# a_4903_15345# 0
C504 VDPWR w_9490_15543# 0.18191f
C505 a_3229_5051# a_2706_5051# 0
C506 a_9877_10533# a_10813_13753# 0.00193f
C507 sky130_fd_sc_hd__mux4_1_0.A0 w_17940_16403# 0.00546f
C508 VGND a_12135_15219# 0.32171f
C509 a_6362_1783# VDPWR 0.20684f
C510 w_12866_5378# a_13411_5463# 0.01092f
C511 a_5895_14763# VGND 0.00618f
C512 a_4905_12113# a_6129_12927# 0
C513 a_7751_14003# a_6389_13769# 0
C514 a_13385_4845# VDPWR 0.37941f
C515 a_18128_16189# sky130_fd_sc_hd__mux4_1_0.A0 0.03043f
C516 a_11289_1773# VGND 0
C517 w_4432_13071# a_4513_14775# 0
C518 a_14325_4589# a_14136_4955# 0
C519 a_11385_1773# a_11553_1773# 0
C520 a_5765_5043# VDPWR 0.00114f
C521 a_14946_4905# a_14864_4585# 0.07951f
C522 a_8566_2145# VDPWR 0
C523 a_12509_4593# a_13439_4955# 0.04534f
C524 a_5975_5299# a_6392_5043# 0.03016f
C525 VDPWR a_15672_4585# 0.21095f
C526 a_11499_2029# w_11008_1688# 0.10454f
C527 w_4538_13995# a_4625_15373# 0
C528 a_24407_14651# sky130_fd_sc_hd__mux4_1_0.A0 0
C529 a_11541_5723# a_8785_5039# 0
C530 a_11178_4593# a_11230_4567# 0.1439f
C531 a_9467_13091# VDPWR 0.38927f
C532 a_5636_5017# a_5584_5043# 0.1439f
C533 a_9725_5837# a_9332_5445# 0.02301f
C534 a_5809_14763# a_6087_14735# 0.1109f
C535 a_4847_14525# a_6629_15387# 0.29596f
C536 a_15071_1765# sky130_fd_sc_hd__mux4_1_0.A2 0
C537 a_23731_14309# sky130_fd_sc_hd__mux4_1_0.A2 0
C538 a_10088_5471# a_7845_5295# 0
C539 a_9599_10561# a_9811_11277# 0
C540 a_15113_5459# a_14888_5433# 0.00487f
C541 VGND w_10872_13125# 0.02002f
C542 a_2259_2047# a_2145_2157# 0
C543 a_9865_15329# a_11089_13753# 0
C544 a_11595_5833# VGND 0.20021f
C545 a_13315_2025# a_13369_2135# 0.03622f
C546 a_5975_12927# a_6129_12927# 0.00401f
C547 a_4213_5047# VGND 0.01521f
C548 a_11499_2029# a_11385_1773# 0
C549 a_13369_2135# w_12824_1684# 0
C550 a_4849_11293# w_5712_14949# 0.08584f
C551 a_15309_4951# sky130_fd_sc_hd__mux4_1_0.A3 0
C552 a_9811_11277# a_11906_13629# 0
C553 a_7751_14003# a_7669_14003# 0.00695f
C554 a_11351_13753# a_11089_13753# 0
C555 a_10813_13753# a_9597_13793# 0
C556 a_14946_4905# a_13439_4589# 0
C557 a_10088_5471# VDPWR 0.2062f
C558 a_8232_1779# a_6885_1783# 0.08907f
C559 a_9875_13765# a_10965_11919# 0
C560 a_7731_5405# a_7506_5013# 0.00559f
C561 a_15071_1765# VGND 0
C562 a_14325_4589# a_15281_5825# 0
C563 a_12135_15219# a_10857_14747# 0
C564 a_23731_14309# VGND 0.12065f
C565 w_1768_1706# a_1868_1791# 0.01793f
C566 a_14975_1765# VDPWR 0.00115f
C567 w_11078_4508# a_11986_4959# 0.00139f
C568 a_15309_4951# w_14764_4500# 0
C569 a_13147_5463# VGND 0
C570 a_3738_1787# w_3638_1702# 0.01793f
C571 a_12976_1743# a_13369_2135# 0.02301f
C572 a_14864_4585# VDPWR 0.09402f
C573 a_7899_5039# a_8262_5039# 0.00985f
C574 a_3040_5417# VGND 0.00244f
C575 w_10868_12105# a_11243_11891# 0.02153f
C576 a_9809_14509# a_9725_14509# 0.00206f
C577 a_9809_14509# w_9402_14723# 0.02435f
C578 a_16195_4585# w_16764_4814# 0.09504f
C579 a_17125_4938# w_16764_4814# 0.04809f
C580 a_11160_1747# ua[5] 0
C581 a_12631_13987# a_12135_15219# 0.16709f
C582 VGND a_9585_4963# 0.00223f
C583 a_7113_13395# a_7919_14003# 0.00207f
C584 a_4015_2153# VDPWR 0
C585 a_24152_14385# ui_in[1] 0.02237f
C586 a_15255_4841# a_15141_4585# 0
C587 a_11049_14719# w_11718_13593# 0
C588 w_10868_12105# a_10965_11919# 0.05631f
C589 w_5786_13983# a_7173_15235# 0
C590 a_7731_5039# sky130_fd_sc_hd__mux4_1_0.A3 0
C591 a_11049_14719# a_11597_15219# 0.08954f
C592 a_10639_4597# a_11230_4567# 0.11887f
C593 a_6389_13769# a_4839_12857# 0.04676f
C594 VDPWR a_2313_1791# 0.17194f
C595 a_3738_1787# a_3790_1761# 0.1439f
C596 a_11569_4849# a_11455_4593# 0
C597 a_13439_4589# VDPWR 0.17474f
C598 a_13369_1769# a_13315_2025# 0.00386f
C599 a_12481_5467# VGND 0.75065f
C600 a_10983_13753# a_9799_16073# 0.00246f
C601 a_2706_5417# a_2289_5307# 0.06611f
C602 w_18554_16401# a_19510_16177# 0
C603 a_9809_14509# a_9875_13765# 0.0012f
C604 a_13369_1769# w_12824_1684# 0.01092f
C605 a_4849_11293# a_4839_12857# 0.82158f
C606 a_11906_13629# a_11824_13629# 0.00477f
C607 a_4903_15345# a_7173_15235# 0
C608 VDPWR a_10983_13753# 0
C609 a_9801_12841# a_11089_13753# 0.00253f
C610 VGND a_9725_14509# 0.00834f
C611 w_19322_16391# VDPWR 0.07226f
C612 VGND w_9402_14723# 0.07437f
C613 a_2217_5025# VDPWR 1.29284f
C614 VGND a_7173_15235# 0.32171f
C615 a_6281_11907# a_6389_13769# 0.00255f
C616 VDPWR a_13411_5829# 0.00606f
C617 a_4763_14775# a_4847_14525# 0.07979f
C618 a_10813_13753# w_11718_13593# 0.00132f
C619 a_13243_5463# VGND 0
C620 a_13369_1769# a_12976_1743# 0.02283f
C621 a_2217_5025# a_1950_5025# 0.08244f
C622 a_4839_12857# a_7669_14003# 0
C623 a_4910_5413# a_5099_5047# 0
C624 a_4546_1787# VGND 0.01333f
C625 a_6281_11907# a_4849_11293# 0.00683f
C626 a_8755_1779# a_9629_2033# 0.21161f
C627 a_1920_1765# a_1868_1791# 0.1439f
C628 a_6885_1783# sky130_fd_sc_hd__mux4_1_0.A2 0.00266f
C629 a_14846_1739# w_14694_1680# 0.05213f
C630 a_24407_14651# a_24234_14385# 0.00222f
C631 a_4837_16089# a_6127_13769# 0.00702f
C632 VDPWR a_2049_2157# 0
C633 a_5945_2039# a_7476_1753# 0.00446f
C634 a_3229_5051# w_1798_4966# 0.02026f
C635 a_4880_2153# a_2187_1765# 0
C636 a_4763_14775# a_4635_13809# 0
C637 a_9875_13765# VGND 0.70497f
C638 a_9801_12841# a_9683_13793# 0
C639 VDPWR a_10116_4597# 0.30078f
C640 a_4765_11543# a_4849_11293# 0.08177f
C641 w_4430_16303# a_4847_14525# 0
C642 a_15227_5715# a_16167_5459# 0.13856f
C643 a_9877_10533# w_9404_11491# 0
C644 a_1920_1765# a_2145_1791# 0.00487f
C645 ua[4] VGND 0
C646 VGND a_15017_5459# 0
C647 a_6281_11907# a_7669_14003# 0.19153f
C648 a_2217_5025# a_3768_5047# 0.00167f
C649 a_12481_5467# w_12894_4504# 0
C650 a_7635_5039# a_7506_5013# 0.00758f
C651 a_5851_13769# a_7173_15235# 0
C652 w_5484_4958# a_2217_5025# 0.00152f
C653 VDPWR w_6074_6018# 0.06609f
C654 VGND a_6885_1783# 0.67804f
C655 a_13385_4845# a_13357_5719# 0.00177f
C656 VDPWR a_11091_12911# 0
C657 a_14794_1765# w_14694_1680# 0.01793f
C658 a_5099_5047# a_6029_5409# 0.04534f
C659 sky130_fd_sc_hd__mux4_1_0.A3 a_16167_5459# 0.00975f
C660 VDPWR a_17339_4938# 0.00182f
C661 a_5945_2039# a_6362_2149# 0.06611f
C662 a_4903_15345# a_4513_14775# 0.00566f
C663 a_9467_13091# a_4915_10549# 0.00237f
C664 a_4129_2043# VGND 1.20051f
C665 a_9877_10533# a_11051_11919# 0
C666 sky130_fd_sc_hd__mux4_1_0.A3 a_24774_14701# 0
C667 a_13439_4955# a_13271_4955# 0
C668 a_12481_5467# a_8785_5039# 0.04118f
C669 a_2313_1791# a_2676_1791# 0.00985f
C670 w_10868_12105# VGND 0.02048f
C671 VDPWR w_6570_15449# 0.08494f
C672 VGND a_4513_14775# 0.29736f
C673 w_17066_16401# sky130_fd_sc_hd__mux4_1_0.A0 0.00801f
C674 a_14846_1739# a_15239_2131# 0.02301f
C675 sky130_fd_sc_hd__mux4_1_0.A3 a_8262_5039# 0
C676 a_23731_14309# a_23677_14701# 0.09132f
C677 a_9699_4853# a_9585_4597# 0
C678 a_9865_15329# a_10937_12911# 0
C679 a_6862_13645# w_6570_15449# 0
C680 ui_in[0] a_24407_14651# 0.00112f
C681 a_11623_4959# a_10639_4597# 0.04534f
C682 VGND a_5735_2149# 0.00305f
C683 ena clk 0.03102f
C684 VDPWR a_24241_14651# 0.25337f
C685 a_9489_4963# sky130_fd_sc_hd__mux4_1_0.A3 0
C686 VGND a_5831_1783# 0
C687 a_7869_2145# a_7605_2145# 0
C688 a_4711_15373# a_4847_14525# 0
C689 a_12881_13987# a_12075_13379# 0.00207f
C690 w_4432_13071# a_4839_12857# 0.02723f
C691 VDPWR a_14255_1769# 1.04578f
C692 a_19510_16177# sky130_fd_sc_hd__mux4_1_0.A0 0.05714f
C693 a_9717_12841# VGND 0.00847f
C694 VDPWR w_21318_16395# 0.07403f
C695 VGND a_16486_16197# 0.25569f
C696 a_10639_4597# a_11623_4593# 0.08312f
C697 a_12509_4593# a_12320_4959# 0
C698 w_5906_12121# a_6003_11935# 0.05631f
C699 a_13439_4955# sky130_fd_sc_hd__mux4_1_0.A3 0
C700 a_9865_15329# a_12075_13379# 0
C701 w_14764_4500# a_15309_4585# 0.01092f
C702 a_19510_16177# a_20384_16179# 0.10121f
C703 VGND a_4015_1787# 0
C704 a_24962_14701# sky130_fd_sc_hd__mux4_1_0.VPB 0.07712f
C705 a_4213_5413# w_3668_4962# 0
C706 a_5809_14763# a_4847_14525# 0.00524f
C707 a_9597_13793# a_9589_12125# 0
C708 a_11958_5467# VDPWR 0.20395f
C709 a_11351_13753# a_12075_13379# 0.06159f
C710 a_7815_2035# a_9290_1751# 0.00511f
C711 a_15071_2131# a_15185_2021# 0
C712 w_9394_13055# VDPWR 0.16326f
C713 VGND a_15309_4951# 0.00129f
C714 a_7845_5295# w_7354_4954# 0.10454f
C715 w_20196_16393# sky130_fd_sc_hd__mux4_1_0.A0 0.00551f
C716 a_11595_5833# a_11541_5723# 0.03622f
C717 a_4503_16339# a_4903_15345# 0
C718 a_9865_15329# w_11532_15433# 0
C719 VGND w_5906_12121# 0.02048f
C720 a_13385_4845# a_14325_4589# 0.13962f
C721 a_5999_1783# a_5831_1783# 0
C722 VDPWR a_6805_15235# 0.00151f
C723 a_13439_4955# a_13046_4563# 0.02301f
C724 a_17254_16187# w_16298_16411# 0
C725 a_13018_5437# a_13411_5463# 0.02283f
C726 w_20196_16393# a_20384_16179# 0.02658f
C727 a_4503_16339# VGND 0.28566f
C728 a_8755_1779# w_9138_1692# 0.24998f
C729 VDPWR w_7354_4954# 0.51208f
C730 sky130_fd_sc_hd__mux4_1_0.A3 sky130_fd_sc_hd__mux4_1_0.A0 0.00455f
C731 a_14325_4589# a_15672_4585# 0.08907f
C732 a_6389_13769# a_6127_13769# 0
C733 a_4837_16089# a_6087_14735# 0.29394f
C734 a_5975_5299# a_6392_5409# 0.06611f
C735 a_15239_1765# sky130_fd_sc_hd__mux4_1_0.A2 0
C736 a_11108_1773# w_11008_1688# 0.01793f
C737 a_11150_5467# VDPWR 0.07689f
C738 a_6726_5409# VDPWR 0
C739 a_3820_5021# VDPWR 0.29445f
C740 a_9360_4571# a_8262_5039# 0
C741 a_2289_5307# a_2175_5051# 0
C742 a_9809_14509# a_9557_14759# 0
C743 a_2313_2157# a_2049_2157# 0
C744 VDPWR a_9477_11527# 0.3853f
C745 a_4849_11293# a_6127_13769# 0
C746 a_23511_14335# sky130_fd_sc_hd__mux4_1_0.A1 0.04403f
C747 VGND a_4753_16339# 0.01705f
C748 a_9489_4963# a_9360_4571# 0.00792f
C749 a_9801_12841# a_10937_12911# 0.30276f
C750 a_5851_13769# w_5906_12121# 0
C751 a_7731_5039# VGND 0
C752 a_7815_2035# a_7869_2145# 0.03622f
C753 a_11986_4593# VDPWR 0.20847f
C754 a_14297_5463# a_13774_5463# 0
C755 a_9725_5837# a_9671_5727# 0.03622f
C756 a_15239_1765# VGND 0.01387f
C757 a_4597_11543# a_4849_11293# 0
C758 a_6029_5409# sky130_fd_sc_hd__mux4_1_0.A3 0
C759 a_13411_5829# a_13357_5719# 0.03622f
C760 a_12439_1773# a_14255_1769# 0
C761 a_5809_14763# a_5975_12927# 0
C762 a_17125_5265# a_16195_4585# 0.00499f
C763 a_12881_13987# a_9877_10533# 0
C764 w_9180_5386# a_11202_5441# 0
C765 VGND a_7751_14003# 0
C766 VDPWR a_4753_16089# 0.00472f
C767 a_11230_4567# a_11455_4593# 0.00487f
C768 a_9801_12841# a_9549_13091# 0
C769 a_9597_13793# w_9500_13979# 0.05631f
C770 a_10046_1777# a_9629_2033# 0.03016f
C771 a_9801_12841# a_12075_13379# 0.00444f
C772 a_12481_5467# a_11541_5723# 0.13811f
C773 a_23677_14335# sky130_fd_sc_hd__mux4_1_0.A0 0
C774 a_14325_4589# a_14864_4585# 0.0725f
C775 a_2187_1765# w_5454_1698# 0.00152f
C776 a_11569_4849# a_12994_4589# 0
C777 a_3820_5021# a_3768_5047# 0.1439f
C778 a_2259_2047# a_3738_1787# 0
C779 VDPWR a_12320_4593# 0
C780 a_4903_15345# w_5712_14949# 0.00546f
C781 w_9208_4512# a_10116_4963# 0.00139f
C782 a_6635_15235# w_6570_15449# 0.08205f
C783 VDPWR a_12924_1769# 0.07449f
C784 a_2289_5307# VGND 1.20002f
C785 a_3199_1791# a_3738_1787# 0.0725f
C786 a_15309_4951# a_8785_5039# 0
C787 a_5809_14763# w_5910_13141# 0
C788 w_9208_4512# a_11178_4593# 0.00188f
C789 a_14916_4559# a_15045_4951# 0.00792f
C790 a_9557_14759# VGND 0.00172f
C791 a_9419_2143# VDPWR 0
C792 a_6915_5043# w_7354_4954# 0.25055f
C793 a_6329_12927# w_6756_13609# 0.04962f
C794 w_9208_4512# a_9753_4597# 0.01092f
C795 a_9865_15329# a_9725_14759# 0.00327f
C796 a_9877_10533# a_11351_13753# 0.00262f
C797 a_6717_15235# a_7173_15235# 0
C798 VGND w_5712_14949# 0.0161f
C799 w_12566_13951# a_12075_13379# 0.04664f
C800 a_6915_5043# a_6726_5409# 0
C801 a_9811_11277# a_9675_12125# 0
C802 a_8232_1779# a_8755_1779# 0
C803 VDPWR a_7919_14003# 0
C804 a_23511_14335# VDPWR 0.00214f
C805 a_15602_1765# VDPWR 0.2057f
C806 a_9699_4853# a_10116_4963# 0.06611f
C807 a_9699_4853# a_11178_4593# 0
C808 w_14736_5374# a_14888_5433# 0.05213f
C809 sky130_fd_sc_hd__mux4_1_0.A1 sky130_fd_sc_hd__mux4_1_0.VPB 0.08143f
C810 a_11569_4849# VDPWR 0.35466f
C811 VGND w_18554_16401# 0.01283f
C812 a_9699_4853# a_9753_4597# 0.00386f
C813 sky130_fd_sc_hd__mux4_1_0.A2 a_24774_14701# 0.00262f
C814 a_14846_1739# a_13315_2025# 0.00446f
C815 VGND a_22274_16171# 0.27907f
C816 VDPWR a_12250_1773# 0
C817 a_14846_1739# w_12824_1684# 0
C818 a_14916_4559# a_15309_4951# 0.02301f
C819 a_4837_16089# a_6021_13769# 0.00246f
C820 VDPWR w_7324_1694# 0.51443f
C821 w_1768_1706# a_2187_1765# 0.25031f
C822 a_9587_15357# a_9799_16073# 0
C823 a_14946_4905# a_14888_5433# 0.00485f
C824 sky130_fd_sc_hd__mux4_1_0.A2 a_15309_4585# 0
C825 VDPWR a_9587_15357# 0.38646f
C826 w_5786_13983# a_4839_12857# 0.08124f
C827 a_10813_13753# a_11243_11891# 0
C828 VGND a_16167_5459# 0.40622f
C829 a_9865_15329# a_9597_13793# 0.00159f
C830 a_13385_4845# a_13802_4589# 0.03016f
C831 a_4913_13781# a_4513_14775# 0
C832 ua[0] sky130_fd_sc_hd__mux4_1_0.A2 0
C833 uio_out[1] uio_out[0] 0.03102f
C834 a_6635_15235# a_6805_15235# 0.00167f
C835 a_6389_13769# a_6087_14735# 0.00427f
C836 a_14794_1765# a_13315_2025# 0
C837 VDPWR w_9502_10747# 0.166f
C838 a_6003_11935# a_4839_12857# 0
C839 VGND a_24774_14701# 0.06373f
C840 VDPWR a_13201_2135# 0
C841 a_14794_1765# w_12824_1684# 0.00188f
C842 a_10088_5471# a_9671_5727# 0.03016f
C843 a_4903_15345# a_4839_12857# 0.1369f
C844 a_14946_4905# a_15113_5825# 0
C845 a_5606_1757# w_5454_1698# 0.05213f
C846 VGND a_8262_5039# 0.01509f
C847 a_4849_11293# a_6087_14735# 0.00179f
C848 sky130_fd_sc_hd__mux4_1_0.A3 a_24234_14385# 0.07599f
C849 a_5895_14763# a_7173_15235# 0
C850 w_9208_4512# a_10639_4597# 0.02026f
C851 sky130_fd_sc_hd__mux4_1_0.A3 w_16764_4814# 0.03021f
C852 VGND a_15309_4585# 0
C853 a_9867_12097# w_9404_11491# 0.00119f
C854 w_9394_13055# a_4915_10549# 0.00179f
C855 a_6281_11907# w_5786_13983# 0
C856 a_4015_2153# a_4183_2153# 0
C857 VGND a_4839_12857# 1.32139f
C858 a_9809_14509# a_11049_14719# 0.3196f
C859 a_3919_1787# VGND 0
C860 a_9877_10533# a_9801_12841# 0.00243f
C861 ua[0] VGND 0.06916f
C862 a_9489_4963# VGND 0.00325f
C863 a_12439_1773# a_12924_1769# 0.07531f
C864 a_4880_2153# VDPWR 0
C865 VDPWR sky130_fd_sc_hd__mux4_1_0.VPB 0.22983f
C866 VDPWR w_4440_14739# 0.16205f
C867 a_6281_11907# a_6003_11935# 0.11706f
C868 a_9801_12841# a_9725_14759# 0.00187f
C869 a_9589_12125# a_9867_12097# 0.1206f
C870 a_9461_5471# a_9725_5471# 0
C871 a_11051_11919# a_9867_12097# 0
C872 a_9699_4853# a_10639_4597# 0.13962f
C873 a_13439_4955# VGND 0.19548f
C874 VDPWR a_14888_5433# 0.30504f
C875 a_9877_10533# w_12566_13951# 0.0566f
C876 a_10046_1777# w_9138_1692# 0.01154f
C877 a_8755_1779# sky130_fd_sc_hd__mux4_1_0.A2 0.00258f
C878 sky130_fd_sc_hd__mux4_1_0.A2 sky130_fd_sc_hd__mux4_1_0.A0 0
C879 a_7869_2145# a_7701_2145# 0
C880 a_4913_13781# w_5906_12121# 0
C881 a_9465_16323# w_9392_16287# 0.06993f
C882 VDPWR a_2706_5051# 0.20629f
C883 a_6281_11907# VGND 0.5959f
C884 a_11767_15219# a_11049_14719# 0.00366f
C885 a_11291_12911# VDPWR 0.23898f
C886 a_11455_4593# a_11623_4593# 0
C887 a_24318_14385# VDPWR 0
C888 sky130_fd_sc_hd__mux4_1_0.A2 a_7476_1753# 0.00206f
C889 a_15644_5459# a_14297_5463# 0.08907f
C890 a_9477_11527# a_4915_10549# 0.00232f
C891 a_11569_4849# a_11986_4959# 0.06611f
C892 a_1920_1765# a_2187_1765# 0.08244f
C893 a_12481_5467# a_13147_5463# 0
C894 a_9809_14509# a_10813_13753# 0
C895 a_15113_5825# VDPWR 0
C896 a_3919_2153# a_3738_1787# 0
C897 a_5851_13769# a_4839_12857# 0.13074f
C898 a_4765_11543# VGND 0.02702f
C899 a_11455_4959# a_11569_4849# 0
C900 VGND a_11049_14719# 0.35053f
C901 ui_in[0] sky130_fd_sc_hd__mux4_1_0.A3 0.08702f
C902 a_13147_5829# sky130_fd_sc_hd__mux4_1_0.A3 0
C903 a_16167_5459# a_8785_5039# 0.1717f
C904 a_9875_13765# w_10872_13125# 0.09336f
C905 uio_oe[0] uio_out[7] 0.03102f
C906 a_4910_5413# VGND 0.00246f
C907 a_8755_1779# VGND 0.67634f
C908 VGND sky130_fd_sc_hd__mux4_1_0.A0 0.51517f
C909 a_9801_12841# a_9597_13793# 0.00246f
C910 a_9811_11277# a_11824_13629# 0
C911 a_4765_11543# a_4637_10577# 0
C912 a_9865_15329# a_11597_15219# 0
C913 a_4849_11293# a_4505_13107# 0.00376f
C914 sky130_fd_sc_hd__mux4_1_0.A2 w_14694_1680# 0.02746f
C915 sky130_fd_sc_hd__mux4_1_0.A2 a_6362_2149# 0
C916 VGND a_7476_1753# 0.40126f
C917 a_15017_5825# a_14888_5433# 0.00792f
C918 VGND a_20384_16179# 0.26555f
C919 a_5099_5047# w_3668_4962# 0.02073f
C920 a_6021_13769# a_6389_13769# 0
C921 a_6057_12927# a_4839_12857# 0.00149f
C922 a_11351_13753# w_11718_13593# 0.06723f
C923 a_4837_16089# a_4847_14525# 0.46421f
C924 a_10639_4597# w_11050_5382# 0.00258f
C925 w_10748_13967# a_9799_16073# 0.06973f
C926 a_13439_4589# a_13802_4589# 0.00985f
C927 a_8785_5039# a_8262_5039# 0
C928 a_9699_4853# a_10450_4963# 0.00696f
C929 a_6281_11907# a_5851_13769# 0
C930 w_10748_13967# VDPWR 0.0898f
C931 w_4442_11507# a_4849_11293# 0.02399f
C932 w_11050_5382# a_11595_5467# 0.01092f
C933 w_9138_1692# a_9238_1777# 0.01793f
C934 a_13439_4955# w_12894_4504# 0
C935 a_12292_5467# sky130_fd_sc_hd__mux4_1_0.A3 0
C936 a_4576_5047# w_3668_4962# 0.01154f
C937 a_4849_11293# a_6021_13769# 0
C938 a_10813_13753# VGND 0.15513f
C939 ua[4] a_15071_1765# 0
C940 a_4159_5303# a_4213_5413# 0.03622f
C941 w_9500_13979# a_7669_14003# 0
C942 VGND a_10895_13753# 0.00382f
C943 VGND a_6029_5409# 0.20237f
C944 VGND w_14694_1680# 0.29099f
C945 a_2343_5051# a_2217_5025# 0.0842f
C946 a_11202_5441# sky130_fd_sc_hd__mux4_1_0.A3 0.00521f
C947 a_9597_13793# w_9492_12311# 0
C948 VGND a_6362_2149# 0.18643f
C949 a_11160_1747# a_11553_2139# 0.02301f
C950 a_11916_2139# sky130_fd_sc_hd__mux4_1_0.A2 0
C951 a_7919_14003# a_4915_10549# 0
C952 a_7454_5039# sky130_fd_sc_hd__mux4_1_0.A3 0.00118f
C953 VDPWR a_13201_1769# 0
C954 a_4837_16089# a_4905_12113# 0
C955 a_9599_10561# a_9477_11527# 0.00144f
C956 a_16167_5459# a_17346_5265# 0
C957 a_9475_14759# a_9725_14759# 0.02504f
C958 a_12481_5467# a_13243_5463# 0
C959 a_4585_16339# a_4503_16339# 0.00641f
C960 a_4913_13781# w_5712_14949# 0
C961 a_15239_2131# sky130_fd_sc_hd__mux4_1_0.A2 0.00137f
C962 a_5945_2039# a_5069_1787# 0.21148f
C963 a_11049_14719# a_10857_14747# 0
C964 a_14916_4559# a_15309_4585# 0.02283f
C965 a_7845_5295# a_9725_5471# 0
C966 a_14946_4905# a_13802_4955# 0
C967 a_4837_16089# a_6911_15235# 0.00241f
C968 a_9809_14509# a_10771_14747# 0.00524f
C969 a_13439_4589# a_13175_4589# 0
C970 sky130_fd_sc_hd__mux4_1_0.A3 a_13774_5463# 0
C971 a_9673_15357# a_9865_15329# 0.00101f
C972 a_11916_2139# VGND 0.1864f
C973 w_7354_4954# a_9308_4597# 0.00201f
C974 a_13774_5829# sky130_fd_sc_hd__mux4_1_0.A3 0.00188f
C975 a_5945_2039# a_7424_1779# 0
C976 VDPWR a_9725_5471# 0.16959f
C977 a_8755_1779# a_10046_2143# 0.03325f
C978 a_4915_10549# w_9502_10747# 0.00202f
C979 a_15239_2131# VGND 0.19769f
C980 a_4837_16089# a_5975_12927# 0
C981 VDPWR a_4625_15373# 0.38724f
C982 a_9875_13765# w_9402_14723# 0
C983 a_9801_12841# w_11718_13593# 0.00515f
C984 a_5636_5017# VDPWR 0.29499f
C985 a_4880_1787# VGND 0
C986 a_13385_4845# a_14136_4955# 0.00696f
C987 VGND w_3638_1702# 0.2935f
C988 a_15644_5825# w_14736_5374# 0.00139f
C989 a_5975_5299# VDPWR 0.34514f
C990 VDPWR a_11230_4567# 0.31788f
C991 a_4903_15345# a_6127_13769# 0
C992 a_9597_13793# a_9475_14759# 0.00144f
C993 a_4045_5413# a_4213_5413# 0
C994 a_17053_4938# VDPWR 0
C995 a_4837_16089# w_5910_13141# 0
C996 a_5765_5409# a_5584_5043# 0
C997 sky130_fd_sc_hd__mux4_1_0.A2 a_24234_14385# 0.04346f
C998 a_8113_13753# w_9490_15543# 0.00459f
C999 a_5945_2039# a_6696_2149# 0.00696f
C1000 a_9589_12125# a_11243_11891# 0
C1001 a_10771_14747# VGND 0.13243f
C1002 w_4432_13071# a_4505_13107# 0.06993f
C1003 VDPWR w_5454_1698# 0.5159f
C1004 a_11202_5441# a_10611_5471# 0.11887f
C1005 VGND a_6127_13769# 0.00413f
C1006 a_11051_11919# a_11243_11891# 0
C1007 a_14108_5829# VDPWR 0
C1008 VDPWR a_13802_4955# 0.02429f
C1009 a_12994_4589# a_13175_4955# 0
C1010 a_2676_2157# a_2187_1765# 0.03547f
C1011 a_14946_4905# a_15644_5825# 0.00336f
C1012 VDPWR a_4765_11293# 0.00377f
C1013 a_5861_5043# a_2217_5025# 0
C1014 a_9809_14509# w_9392_16287# 0
C1015 a_9589_12125# a_10965_11919# 0
C1016 VDPWR a_13411_5463# 0.1693f
C1017 a_12631_13987# a_10813_13753# 0
C1018 a_4913_13781# a_4839_12857# 0.44871f
C1019 a_5945_2039# a_5999_2149# 0.03622f
C1020 a_4597_11543# VGND 0.00172f
C1021 a_6389_13769# a_4847_14525# 0
C1022 a_11051_11919# a_10965_11919# 0.00658f
C1023 VGND a_3790_1761# 0.40141f
C1024 a_12439_1773# a_13201_1769# 0
C1025 VGND a_24234_14385# 0.05676f
C1026 VGND w_16764_4814# 0.01288f
C1027 a_4546_1787# a_4129_2043# 0.03016f
C1028 VDPWR w_1798_4966# 0.51758f
C1029 a_10046_1777# sky130_fd_sc_hd__mux4_1_0.A2 0
C1030 a_5636_5017# w_5484_4958# 0.05213f
C1031 a_13357_5719# a_14888_5433# 0.00446f
C1032 a_23677_14701# sky130_fd_sc_hd__mux4_1_0.A0 0.01449f
C1033 a_7815_2035# a_8232_2145# 0.06611f
C1034 a_7845_5295# a_8596_5039# 0.00682f
C1035 a_4755_12857# VDPWR 0.00415f
C1036 a_5975_5299# w_5484_4958# 0.10454f
C1037 a_4849_11293# a_4847_14525# 0.00506f
C1038 ui_in[1] sky130_fd_sc_hd__mux4_1_0.A3 0.07335f
C1039 a_9332_5445# a_9725_5471# 0.02283f
C1040 a_13018_5437# w_11050_5382# 0
C1041 VDPWR a_13175_4955# 0
C1042 a_1950_5025# w_1798_4966# 0.05213f
C1043 a_9599_10561# w_9502_10747# 0.05631f
C1044 a_11150_5467# a_9671_5727# 0
C1045 w_1768_1706# VDPWR 0.51727f
C1046 a_9467_13091# a_9811_11277# 0.00376f
C1047 a_5851_13769# a_6127_13769# 0.00119f
C1048 ui_in[0] sky130_fd_sc_hd__mux4_1_0.A2 0.03574f
C1049 a_5975_5299# a_6915_5043# 0.13962f
C1050 w_10868_12105# a_9875_13765# 0
C1051 a_17125_5265# sky130_fd_sc_hd__mux4_1_0.A3 0
C1052 VDPWR a_8596_5039# 0
C1053 a_15071_1765# a_15239_1765# 0
C1054 VDPWR a_7605_1779# 0.00115f
C1055 a_14946_4905# a_16006_4951# 0.0022f
C1056 a_9465_16323# a_9865_15329# 0
C1057 a_10088_5837# w_9180_5386# 0.00139f
C1058 a_10046_1777# VGND 0.01329f
C1059 a_2145_2157# a_2187_1765# 0
C1060 VGND w_9392_16287# 0.06272f
C1061 a_4635_13809# a_4849_11293# 0.00317f
C1062 w_12866_5378# a_14297_5463# 0.02026f
C1063 a_10771_14747# a_10857_14747# 0.00658f
C1064 a_15644_5825# VDPWR 0.01852f
C1065 a_12320_4959# VGND 0.00281f
C1066 a_11202_5441# a_11427_5467# 0.00487f
C1067 a_4905_12113# a_4849_11293# 0.25265f
C1068 a_14836_5459# a_14888_5433# 0.1439f
C1069 a_4576_5413# a_2217_5025# 0
C1070 w_1798_4966# a_3768_5047# 0.00188f
C1071 a_9801_12841# a_9867_12097# 0.04364f
C1072 a_9715_16323# w_9392_16287# 0.01327f
C1073 ui_in[0] VGND 0.11268f
C1074 a_12509_4593# w_12866_5378# 0.00258f
C1075 VGND w_4540_10763# 0.12086f
C1076 a_3229_5051# a_4213_5413# 0.04534f
C1077 w_5786_13983# a_6087_14735# 0
C1078 VGND a_13147_5829# 0.00333f
C1079 a_11916_1773# sky130_fd_sc_hd__mux4_1_0.A2 0
C1080 sky130_fd_sc_hd__mux4_1_0.A2 a_9238_1777# 0.00119f
C1081 a_15644_5459# a_15227_5715# 0.03016f
C1082 a_21506_16181# sky130_fd_sc_hd__mux4_1_0.A1 0
C1083 a_11455_4959# a_11230_4567# 0.00559f
C1084 a_23677_14335# ui_in[1] 0
C1085 a_9290_1751# VDPWR 0.29556f
C1086 a_11623_4959# VDPWR 0.00948f
C1087 a_4637_10577# w_4540_10763# 0.05631f
C1088 a_3040_5417# a_2289_5307# 0.00696f
C1089 VGND w_9404_11491# 0.07411f
C1090 a_2217_5025# a_2343_5417# 0.0517f
C1091 a_15255_4841# w_14736_5374# 0.00166f
C1092 a_14325_4589# a_14888_5433# 0
C1093 sky130_fd_sc_hd__mux4_1_0.A2 a_13315_2025# 0.00291f
C1094 a_5895_14763# a_4839_12857# 0
C1095 a_4903_15345# a_6087_14735# 0
C1096 a_14846_1739# a_15185_2021# 0.04737f
C1097 a_9683_1777# VDPWR 0.17495f
C1098 a_15644_5459# sky130_fd_sc_hd__mux4_1_0.A3 0
C1099 w_16764_4814# a_8785_5039# 0.17704f
C1100 a_5099_5047# a_6029_5043# 0.08101f
C1101 a_4849_11293# a_5975_12927# 0.18651f
C1102 sky130_fd_sc_hd__mux4_1_0.A2 w_12824_1684# 0.00315f
C1103 VDPWR a_16006_4951# 0
C1104 a_9867_12097# w_9492_12311# 0.0247f
C1105 a_11916_1773# VGND 0.01327f
C1106 VGND a_9589_12125# 0.24254f
C1107 a_12292_5467# VGND 0
C1108 a_11499_2029# a_12924_1769# 0
C1109 VGND a_9238_1777# 0.08667f
C1110 VDPWR a_11623_4593# 0.17434f
C1111 VGND a_6087_14735# 0.35053f
C1112 uo_out[5] uo_out[6] 0.03102f
C1113 a_4129_2043# a_4015_1787# 0
C1114 a_11051_11919# VGND 0.00568f
C1115 a_12881_13987# a_11243_11891# 0
C1116 w_5910_13141# a_4849_11293# 0.05304f
C1117 a_9717_13091# a_9589_12125# 0
C1118 VGND a_11202_5441# 0.40461f
C1119 a_15255_4841# a_14946_4905# 1.1874f
C1120 a_1920_1765# VDPWR 0.30549f
C1121 a_7454_5039# VGND 0.08651f
C1122 w_1768_1706# a_2676_1791# 0.01154f
C1123 VGND a_13315_2025# 1.19935f
C1124 a_12976_1743# sky130_fd_sc_hd__mux4_1_0.A2 0.00202f
C1125 w_4432_13071# a_4847_14525# 0
C1126 a_7506_5013# w_7354_4954# 0.05213f
C1127 VGND w_12824_1684# 0.29354f
C1128 a_2259_2047# a_3010_2157# 0.00696f
C1129 a_9811_11277# a_10983_13753# 0
C1130 a_11049_14719# a_12135_15219# 0.00425f
C1131 a_3199_1791# a_3010_2157# 0
C1132 a_11359_4593# a_11230_4567# 0.00758f
C1133 a_15045_4951# a_15309_4951# 0
C1134 a_23731_14309# a_24774_14701# 0.00253f
C1135 a_11351_13753# a_11243_11891# 0.00255f
C1136 a_7869_2145# VDPWR 0.00911f
C1137 sky130_fd_sc_hd__mux4_1_0.A2 a_14066_1769# 0
C1138 w_7604_13967# a_7113_13395# 0.04664f
C1139 a_11499_2029# a_12250_1773# 0.00682f
C1140 a_21506_16181# VDPWR 0.25743f
C1141 VGND a_13774_5463# 0.01425f
C1142 a_10937_12911# a_11019_12911# 0.00517f
C1143 a_15936_2131# a_15185_2021# 0.00696f
C1144 sky130_fd_sc_hd__mux4_1_0.A1 a_6629_15387# 0.10747f
C1145 a_4503_16339# a_4513_14775# 0.00102f
C1146 VDPWR a_6129_12927# 0
C1147 sky130_fd_sc_hd__mux4_1_0.A3 a_9557_5471# 0
C1148 a_13774_5829# VGND 0.1873f
C1149 a_4635_13809# w_4432_13071# 0.00101f
C1150 w_5712_14949# a_7173_15235# 0
C1151 a_5851_13769# a_6087_14735# 0
C1152 a_12976_1743# VGND 0.40116f
C1153 a_4159_5303# a_4045_5047# 0
C1154 a_4159_5303# a_5099_5047# 0.14245f
C1155 a_9515_1777# VDPWR 0
C1156 a_23731_14309# ua[0] 0
C1157 a_4905_12113# w_4432_13071# 0
C1158 w_1768_1706# a_2313_2157# 0
C1159 a_14066_2135# VDPWR 0
C1160 VGND a_14066_1769# 0
C1161 a_14108_5829# a_13357_5719# 0.00696f
C1162 a_9799_16073# a_9715_16073# 0.00234f
C1163 a_4159_5303# a_4576_5047# 0.03016f
C1164 a_10813_13753# a_12135_15219# 0
C1165 a_14946_4905# a_15978_5825# 0
C1166 a_4713_12141# a_4849_11293# 0
C1167 a_15255_4841# VDPWR 0.35508f
C1168 a_4913_13781# a_6127_13769# 0
C1169 a_11331_5833# sky130_fd_sc_hd__mux4_1_0.A3 0
C1170 VDPWR a_9715_16073# 0.00472f
C1171 a_13357_5719# a_13411_5463# 0.00386f
C1172 VGND a_4505_13107# 0.29689f
C1173 VGND w_9500_13979# 0.11975f
C1174 a_11623_4959# a_11986_4959# 0.00847f
C1175 a_15255_4841# a_16871_4938# 0
C1176 w_11008_1688# a_12924_1769# 0.00227f
C1177 a_11623_4959# a_11455_4959# 0
C1178 a_4903_15345# a_6021_13769# 0.00818f
C1179 a_15141_4951# a_14946_4905# 0.00207f
C1180 a_11091_12911# a_9811_11277# 0
C1181 a_7899_5405# sky130_fd_sc_hd__mux4_1_0.A3 0
C1182 VGND w_4442_11507# 0.07411f
C1183 sky130_fd_sc_hd__mux4_1_0.A2 ui_in[1] 0.24408f
C1184 a_9809_14509# a_9865_15329# 0.15229f
C1185 w_4432_13071# a_5975_12927# 0
C1186 VGND a_6021_13769# 0.00475f
C1187 a_11202_5441# a_8785_5039# 0
C1188 a_12509_4593# a_10639_4597# 0
C1189 uio_oe[1] uio_oe[0] 0.03102f
C1190 a_7847_14003# a_7669_14003# 0.00412f
C1191 VDPWR a_6629_15387# 1.38991f
C1192 ui_in[0] a_23677_14701# 0.02095f
C1193 a_9809_14509# a_11351_13753# 0
C1194 a_4637_10577# w_4442_11507# 0
C1195 a_23731_14309# sky130_fd_sc_hd__mux4_1_0.A0 0.09059f
C1196 a_9801_12841# a_11243_11891# 0.02336f
C1197 VGND w_3668_4962# 0.29364f
C1198 a_10813_13753# w_10872_13125# 0.00142f
C1199 a_6392_5043# a_5099_5047# 0.08907f
C1200 a_18742_16187# a_17254_16187# 0
C1201 a_13369_1769# a_13732_1769# 0.00985f
C1202 w_5712_14949# a_4513_14775# 0
C1203 sky130_fd_sc_hd__mux4_1_0.A3 a_6029_5043# 0
C1204 a_12481_5467# a_13439_4955# 0
C1205 a_23511_14701# sky130_fd_sc_hd__mux4_1_0.A3 0.00138f
C1206 VGND a_4721_13809# 0.00661f
C1207 a_4839_12857# a_7173_15235# 0.00685f
C1208 a_14946_4905# a_16006_4585# 0
C1209 a_5069_1787# sky130_fd_sc_hd__mux4_1_0.A2 0
C1210 VGND ui_in[1] 0.53405f
C1211 a_5099_5047# a_5584_5043# 0.07558f
C1212 a_2343_5051# a_2706_5051# 0.00985f
C1213 a_2259_2047# VGND 1.20011f
C1214 a_3199_1791# VGND 0.67808f
C1215 a_9465_16323# a_9475_14759# 0.00102f
C1216 a_9801_12841# a_10965_11919# 0
C1217 a_12881_13987# VGND 0
C1218 w_12566_13951# a_11243_11891# 0.03664f
C1219 a_4503_16339# a_4753_16339# 0.02504f
C1220 a_10088_5837# sky130_fd_sc_hd__mux4_1_0.A3 0.00192f
C1221 a_17125_5265# VGND 0.00352f
C1222 VDPWR a_2079_5051# 0.00123f
C1223 a_9865_15329# VGND 0.98587f
C1224 a_1920_1765# a_2313_2157# 0.02301f
C1225 a_7424_1779# sky130_fd_sc_hd__mux4_1_0.A2 0.00118f
C1226 a_5851_13769# a_6021_13769# 0.00167f
C1227 a_15141_4951# VDPWR 0
C1228 a_10771_14747# a_12135_15219# 0
C1229 a_15113_5459# a_14297_5463# 0
C1230 w_9394_13055# a_9811_11277# 0.00299f
C1231 VDPWR a_2676_2157# 0.02063f
C1232 a_2079_5051# a_1950_5025# 0.00758f
C1233 a_4910_5047# a_2217_5025# 0
C1234 a_5069_1787# VGND 0.67702f
C1235 a_11351_13753# VGND 0.25955f
C1236 a_6281_11907# a_7173_15235# 0.09936f
C1237 a_4849_11293# w_4538_13995# 0.00123f
C1238 a_15602_2131# sky130_fd_sc_hd__mux4_1_0.A2 0.00187f
C1239 a_11359_4593# a_11623_4593# 0
C1240 a_10569_1777# a_11160_1747# 0.11887f
C1241 w_18554_16401# a_16486_16197# 0
C1242 a_10965_11919# w_9492_12311# 0
C1243 a_9515_2143# VDPWR 0
C1244 a_4515_11543# a_4765_11293# 0.00723f
C1245 a_9360_4571# a_9585_4597# 0.00487f
C1246 a_6696_2149# sky130_fd_sc_hd__mux4_1_0.A2 0
C1247 VGND a_7424_1779# 0.08651f
C1248 a_11089_13753# a_9799_16073# 0.00702f
C1249 w_9208_4512# VDPWR 0.78497f
C1250 VDPWR a_16006_4585# 0
C1251 a_9699_4853# a_7845_5295# 0
C1252 a_13385_4845# a_14864_4585# 0
C1253 w_10674_14933# a_11597_15219# 0
C1254 w_12866_5378# sky130_fd_sc_hd__mux4_1_0.A3 0.00618f
C1255 a_9809_14509# a_9801_12841# 0.20053f
C1256 VDPWR a_11089_13753# 0.0014f
C1257 a_10771_14747# w_10872_13125# 0
C1258 VGND a_15644_5459# 0.01334f
C1259 a_4913_13781# a_6087_14735# 0
C1260 a_15602_2131# VGND 0.18859f
C1261 a_4839_12857# a_4513_14775# 0.00442f
C1262 a_15071_2131# VDPWR 0
C1263 a_9477_11527# a_9811_11277# 0.16782f
C1264 a_5069_1787# a_5999_1783# 0.08097f
C1265 a_5999_2149# sky130_fd_sc_hd__mux4_1_0.A2 0
C1266 a_9875_13765# a_11049_14719# 0
C1267 uo_out[0] uo_out[1] 0.03102f
C1268 a_9671_5727# a_9725_5471# 0.00386f
C1269 VDPWR a_2145_2157# 0
C1270 a_4903_15345# a_4847_14525# 0.15229f
C1271 a_12976_1743# a_13105_2135# 0.00792f
C1272 a_9699_4853# VDPWR 0.60063f
C1273 VGND a_6696_2149# 0.00244f
C1274 a_15672_4951# a_15255_4841# 0.06611f
C1275 w_5786_13983# a_4635_13809# 0
C1276 a_3229_5051# a_4045_5047# 0
C1277 a_9865_15329# a_10857_14747# 0
C1278 a_6717_15235# a_6087_14735# 0.00232f
C1279 a_12292_5467# a_11541_5723# 0.00682f
C1280 w_12866_5378# a_13046_4563# 0.00104f
C1281 a_4763_14775# VDPWR 0.32009f
C1282 a_3229_5051# a_5099_5047# 0.00117f
C1283 VGND a_4847_14525# 0.43095f
C1284 a_4627_12141# a_4849_11293# 0.0022f
C1285 a_13385_4845# a_13439_4589# 0.00386f
C1286 a_13271_4589# VDPWR 0
C1287 a_11202_5441# a_11541_5723# 0.04737f
C1288 VDPWR a_9557_5837# 0
C1289 a_9683_13793# VDPWR 0.003f
C1290 a_4905_12113# a_6003_11935# 0.18618f
C1291 a_5999_2149# VGND 0.20086f
C1292 a_12881_13987# a_12631_13987# 0.00876f
C1293 a_3229_5051# a_4576_5047# 0.08907f
C1294 a_8755_1779# a_6885_1783# 0
C1295 a_15281_5459# a_14888_5433# 0.02283f
C1296 a_4635_13809# a_4903_15345# 0.00159f
C1297 a_9801_12841# VGND 1.32139f
C1298 a_6635_15235# a_6629_15387# 0.1684f
C1299 a_3738_1787# a_2187_1765# 0.00167f
C1300 a_13018_5437# a_12509_4593# 0
C1301 a_6885_1783# a_7476_1753# 0.11887f
C1302 a_6392_5043# sky130_fd_sc_hd__mux4_1_0.A3 0
C1303 VGND a_2049_1791# 0
C1304 a_10813_13753# a_9875_13765# 0.0094f
C1305 a_7919_14003# a_8113_13753# 0
C1306 a_9717_13091# a_9801_12841# 0.08134f
C1307 sky130_fd_sc_hd__mux4_1_0.A3 a_10116_4963# 0
C1308 VGND w_16298_16411# 0.01283f
C1309 VDPWR w_4430_16303# 0.16502f
C1310 a_4635_13809# VGND 0.24546f
C1311 a_11359_4959# a_11178_4593# 0
C1312 a_11178_4593# sky130_fd_sc_hd__mux4_1_0.A3 0
C1313 a_9875_13765# a_10895_13753# 0
C1314 a_23731_14309# a_24234_14385# 0.12294f
C1315 w_5906_12121# a_4839_12857# 0.00131f
C1316 VGND a_9557_5471# 0
C1317 a_13385_4845# a_13411_5829# 0
C1318 a_4905_12113# VGND 0.43935f
C1319 a_17254_16187# sky130_fd_sc_hd__mux4_1_0.A1 0
C1320 w_9208_4512# a_9332_5445# 0
C1321 a_5765_5043# a_2217_5025# 0
C1322 w_12566_13951# VGND 0.00711f
C1323 a_12631_13987# a_11351_13753# 0.00196f
C1324 w_5786_13983# a_5975_12927# 0
C1325 a_3919_2153# VGND 0.00305f
C1326 VDPWR w_11050_5382# 0.51351f
C1327 a_3040_5051# VDPWR 0
C1328 VDPWR a_9683_2143# 0.00879f
C1329 a_5851_13769# a_4847_14525# 0
C1330 VDPWR a_24152_14385# 0.00352f
C1331 a_4913_13781# a_4505_13107# 0
C1332 VGND a_6911_15235# 0.00384f
C1333 a_9585_4597# sky130_fd_sc_hd__mux4_1_0.A2 0
C1334 w_22086_16385# a_21506_16181# 0.05681f
C1335 ui_in[1] a_23677_14701# 0.0594f
C1336 a_6003_11935# a_5975_12927# 0
C1337 VGND w_9492_12311# 0.11704f
C1338 a_9587_15357# a_8113_13753# 0.00113f
C1339 a_3010_1791# VGND 0
C1340 a_11331_5833# VGND 0.00311f
C1341 a_6281_11907# w_5906_12121# 0.02153f
C1342 a_4837_16089# a_5933_13769# 0
C1343 a_16486_16197# sky130_fd_sc_hd__mux4_1_0.A0 0.14964f
C1344 a_4903_15345# a_5975_12927# 0
C1345 a_9597_13793# a_7113_13395# 0
C1346 a_5895_14763# a_6087_14735# 0
C1347 a_2313_2157# a_2676_2157# 0.00847f
C1348 a_10813_13753# w_10868_12105# 0
C1349 w_5910_13141# a_6003_11935# 0
C1350 a_9809_14509# a_9475_14759# 0.1679f
C1351 a_10771_14747# w_9402_14723# 0
C1352 ui_in[4] ui_in[3] 0.03102f
C1353 a_4913_13781# a_6021_13769# 0.00104f
C1354 a_15141_4585# sky130_fd_sc_hd__mux4_1_0.A2 0
C1355 a_5851_13769# a_4635_13809# 0
C1356 VGND a_5975_12927# 0.14511f
C1357 a_4546_1787# w_3638_1702# 0.01154f
C1358 VGND a_7899_5405# 0.20211f
C1359 a_4903_15345# w_5910_13141# 0.00114f
C1360 a_2343_5051# w_1798_4966# 0.01092f
C1361 w_7604_13967# VDPWR 0.07722f
C1362 a_13018_5437# a_13243_5829# 0.00559f
C1363 a_9585_4597# VGND 0
C1364 a_9332_5445# a_9557_5837# 0.00559f
C1365 VDPWR a_4711_15373# 0.00333f
C1366 a_9801_12841# a_10857_14747# 0
C1367 a_23731_14309# ui_in[0] 0.48787f
C1368 a_4837_16089# a_7113_13395# 0
C1369 VGND w_5910_13141# 0.02002f
C1370 a_4913_13781# a_4721_13809# 0.00222f
C1371 a_17254_16187# VDPWR 0.26221f
C1372 VDPWR a_13369_2135# 0.00905f
C1373 a_18742_16187# w_17940_16403# 0
C1374 a_5809_14763# VDPWR 0.1486f
C1375 a_9875_13765# a_10771_14747# 0
C1376 sky130_fd_sc_hd__mux4_1_0.A2 a_15185_2021# 0.1531f
C1377 uio_in[6] uio_in[5] 0.03102f
C1378 VGND a_6029_5043# 0.01597f
C1379 a_4627_12141# w_4432_13071# 0
C1380 sky130_fd_sc_hd__mux4_1_0.A1 a_12075_13379# 0.03027f
C1381 a_10639_4597# sky130_fd_sc_hd__mux4_1_0.A3 0
C1382 a_10380_2143# a_9629_2033# 0.00696f
C1383 a_23511_14701# VGND 0.00202f
C1384 a_15255_4841# a_14325_4589# 0.21188f
C1385 a_5975_5299# a_7506_5013# 0.00446f
C1386 a_2313_2157# a_2145_2157# 0
C1387 a_18742_16187# a_18128_16189# 0.10376f
C1388 a_11595_5833# a_11202_5441# 0.02301f
C1389 a_13105_1769# a_13369_1769# 0
C1390 a_9360_4571# a_9753_4597# 0.02283f
C1391 a_12631_13987# a_9801_12841# 0
C1392 sky130_fd_sc_hd__mux4_1_0.A3 a_11595_5467# 0
C1393 a_9475_14759# VGND 0.29736f
C1394 a_4839_12857# w_5712_14949# 0.08813f
C1395 a_5636_5017# a_5861_5043# 0.00487f
C1396 a_4129_2043# a_4880_1787# 0.00682f
C1397 a_4129_2043# w_3638_1702# 0.10454f
C1398 a_5851_13769# a_5975_12927# 0
C1399 a_5975_5299# a_5861_5043# 0
C1400 a_10088_5837# VGND 0.22304f
C1401 a_6281_11907# a_7751_14003# 0.00373f
C1402 sky130_fd_sc_hd__mux4_1_0.A1 w_11532_15433# 0
C1403 a_9717_13091# a_9475_14759# 0
C1404 VGND a_15185_2021# 1.19592f
C1405 a_7635_5405# sky130_fd_sc_hd__mux4_1_0.A3 0
C1406 VDPWR a_8232_2145# 0.01966f
C1407 a_15281_5825# a_14888_5433# 0.02301f
C1408 a_12631_13987# w_12566_13951# 0.05168f
C1409 a_10937_12911# a_9799_16073# 0
C1410 a_5851_13769# w_5910_13141# 0.00142f
C1411 a_7815_2035# w_9138_1692# 0
C1412 a_11291_12911# a_9811_11277# 0.00976f
C1413 a_10937_12911# VDPWR 0.1592f
C1414 a_6057_12927# a_5975_12927# 0.00517f
C1415 w_4528_15559# a_4625_15373# 0.05631f
C1416 VGND a_4713_12141# 0.00662f
C1417 a_6392_5409# a_5099_5047# 0.03325f
C1418 a_4129_2043# a_3790_1761# 0.04737f
C1419 a_15113_5459# a_15227_5715# 0
C1420 VGND a_7847_14003# 0
C1421 sky130_fd_sc_hd__mux4_1_0.A2 a_11553_2139# 0
C1422 a_15113_5825# a_15281_5825# 0
C1423 a_9799_16073# a_12075_13379# 0
C1424 w_9394_13055# a_9467_13091# 0.06993f
C1425 a_13732_2135# a_13369_2135# 0.00847f
C1426 a_4159_5303# VGND 1.20044f
C1427 a_11986_4593# w_11078_4508# 0.01154f
C1428 a_9549_13091# VDPWR 0.02512f
C1429 a_13369_1769# VDPWR 0.17556f
C1430 VDPWR a_12075_13379# 0.24586f
C1431 w_12866_5378# VGND 0.31514f
C1432 w_10748_13967# a_8113_13753# 0
C1433 ua[0] a_24774_14701# 0.00406f
C1434 a_15113_5459# sky130_fd_sc_hd__mux4_1_0.A3 0
C1435 a_15239_1765# w_14694_1680# 0.01092f
C1436 a_5933_13769# a_6389_13769# 0
C1437 a_5861_5409# VDPWR 0
C1438 a_9683_13793# a_4915_10549# 0
C1439 a_10639_4597# a_10611_5471# 0.00251f
C1440 w_11532_15433# a_9799_16073# 0.09702f
C1441 a_12881_13987# a_12135_15219# 0
C1442 VGND a_3949_5047# 0
C1443 a_14975_1765# a_14255_1769# 0
C1444 a_10611_5471# a_11595_5467# 0.08312f
C1445 a_12439_1773# a_13369_2135# 0.04534f
C1446 w_10748_13967# a_9811_11277# 0.10705f
C1447 a_11160_1747# VDPWR 0.29475f
C1448 a_4913_13781# a_4847_14525# 0.0012f
C1449 VGND a_11553_2139# 0.20244f
C1450 VDPWR w_11532_15433# 0.08492f
C1451 w_18554_16401# sky130_fd_sc_hd__mux4_1_0.A0 0.00562f
C1452 a_4723_10577# VGND 0.00697f
C1453 a_9865_15329# a_12135_15219# 0
C1454 a_5933_13769# a_4849_11293# 0
C1455 a_5945_2039# a_2187_1765# 0
C1456 a_14946_4905# a_16195_4585# 0.08128f
C1457 a_14946_4905# a_17125_4938# 0.00161f
C1458 a_7173_15235# a_6087_14735# 0.00425f
C1459 a_22274_16171# sky130_fd_sc_hd__mux4_1_0.A0 0.15979f
C1460 uio_in[2] uio_in[1] 0.03102f
C1461 a_11178_4593# sky130_fd_sc_hd__mux4_1_0.A2 0
C1462 a_9877_10533# sky130_fd_sc_hd__mux4_1_0.A1 0.22585f
C1463 a_2217_5025# w_6074_6018# 0.02708f
C1464 a_5765_5409# VDPWR 0
C1465 a_9467_13091# a_9477_11527# 0.00102f
C1466 a_4015_1787# a_3790_1761# 0.00487f
C1467 a_7701_1779# sky130_fd_sc_hd__mux4_1_0.A2 0
C1468 a_9753_4597# sky130_fd_sc_hd__mux4_1_0.A2 0
C1469 a_11351_13753# a_12135_15219# 0.00152f
C1470 VDPWR a_4213_5413# 0.00874f
C1471 a_7113_13395# a_6389_13769# 0.06159f
C1472 a_4723_10577# a_4637_10577# 0.00658f
C1473 a_6717_15235# a_4847_14525# 0.00159f
C1474 a_22274_16171# a_20384_16179# 0
C1475 a_12481_5467# a_13774_5463# 0.08907f
C1476 a_1868_1791# VGND 0.09509f
C1477 a_11291_12911# a_11824_13629# 0.10646f
C1478 a_10569_1777# a_9629_2033# 0.13962f
C1479 a_4913_13781# a_4635_13809# 0.1205f
C1480 a_4213_5047# w_3668_4962# 0.01092f
C1481 VDPWR w_22960_16387# 0.06784f
C1482 a_7869_1779# w_7324_1694# 0.01092f
C1483 a_12481_5467# a_13774_5829# 0.03325f
C1484 a_4913_13781# a_4905_12113# 0.00627f
C1485 a_8232_1779# a_7815_2035# 0.03016f
C1486 a_15141_4585# a_14916_4559# 0.00487f
C1487 a_6281_11907# a_4839_12857# 0.02336f
C1488 a_11569_4849# w_11078_4508# 0.10454f
C1489 a_4903_15345# w_4538_13995# 0.00397f
C1490 a_10422_5837# sky130_fd_sc_hd__mux4_1_0.A3 0
C1491 a_7113_13395# a_4849_11293# 0.00118f
C1492 VGND a_6392_5043# 0.01331f
C1493 sky130_fd_sc_hd__mux4_1_0.A0 a_24774_14701# 0
C1494 VGND a_10116_4963# 0.1833f
C1495 a_11178_4593# VGND 0.07994f
C1496 sky130_fd_sc_hd__mux4_1_0.A2 a_7605_2145# 0
C1497 a_4045_5413# VGND 0.00231f
C1498 a_2145_1791# VGND 0
C1499 a_7701_1779# VGND 0
C1500 VGND w_4538_13995# 0.11975f
C1501 VGND a_5584_5043# 0.08665f
C1502 a_9865_15329# w_10872_13125# 0.00114f
C1503 a_9753_4597# VGND 0.01261f
C1504 a_15936_1765# a_15185_2021# 0.00682f
C1505 a_5554_1783# w_5454_1698# 0.01793f
C1506 a_13018_5437# sky130_fd_sc_hd__mux4_1_0.A3 0.00516f
C1507 w_9208_4512# a_9308_4597# 0.01793f
C1508 ui_in[5] ui_in[6] 0.03102f
C1509 w_7604_13967# a_4915_10549# 0.05671f
C1510 a_23731_14309# ui_in[1] 0.35239f
C1511 sky130_fd_sc_hd__mux4_1_0.A1 a_18128_16189# 0
C1512 a_9290_1751# a_9419_1777# 0.00758f
C1513 a_7113_13395# a_7669_14003# 0.28206f
C1514 a_23511_14701# a_23677_14701# 0.05551f
C1515 a_17125_4938# VDPWR 0.06504f
C1516 a_11427_5467# a_11595_5467# 0
C1517 a_16195_4585# VDPWR 0.2778f
C1518 w_12866_5378# a_8785_5039# 0.00344f
C1519 a_9877_10533# a_9799_16073# 0.01618f
C1520 a_13369_1769# a_12439_1773# 0.08096f
C1521 a_2343_5417# w_1798_4966# 0
C1522 w_14736_5374# a_14297_5463# 0.25055f
C1523 a_11289_2139# a_11553_2139# 0
C1524 a_9587_15357# w_9490_15543# 0.05631f
C1525 w_10868_12105# a_9589_12125# 0
C1526 a_9683_1777# a_9419_1777# 0
C1527 VGND a_7605_2145# 0.00305f
C1528 a_4913_13781# a_5975_12927# 0.08477f
C1529 a_9877_10533# VDPWR 0.59881f
C1530 a_16195_4585# a_16871_4938# 0.15182f
C1531 a_4513_14775# a_6087_14735# 0
C1532 uio_out[6] uio_out[7] 0.03102f
C1533 a_13018_5437# a_13046_4563# 0
C1534 w_9500_13979# a_7173_15235# 0
C1535 VDPWR a_9725_14759# 0.32009f
C1536 a_5945_2039# a_5606_1757# 0.04737f
C1537 a_8262_5405# sky130_fd_sc_hd__mux4_1_0.A3 0
C1538 a_4627_12141# a_6003_11935# 0
C1539 a_10639_4597# sky130_fd_sc_hd__mux4_1_0.A2 0
C1540 a_4913_13781# w_5910_13141# 0.09336f
C1541 a_6392_5409# sky130_fd_sc_hd__mux4_1_0.A3 0
C1542 a_5851_13769# w_4538_13995# 0
C1543 a_3738_1787# VDPWR 0.07401f
C1544 a_9801_12841# a_12135_15219# 0.00685f
C1545 a_14946_4905# a_14297_5463# 0.01842f
C1546 a_9809_14509# w_10674_14933# 0.00381f
C1547 a_5975_5299# a_6726_5043# 0.00682f
C1548 a_11958_5833# w_11050_5382# 0.00139f
C1549 a_8566_1779# sky130_fd_sc_hd__mux4_1_0.A2 0
C1550 a_10422_5837# a_10611_5471# 0
C1551 VDPWR w_17940_16403# 0.07531f
C1552 a_4627_12141# VGND 0.24254f
C1553 a_9875_13765# w_9500_13979# 0.01958f
C1554 a_12509_4593# a_14946_4905# 0
C1555 w_12566_13951# a_12135_15219# 0.11864f
C1556 a_3820_5021# a_2217_5025# 0.00242f
C1557 a_10639_4597# VGND 0.65621f
C1558 a_2343_5051# a_2079_5051# 0
C1559 VDPWR a_18128_16189# 0.25317f
C1560 a_12292_5833# sky130_fd_sc_hd__mux4_1_0.A3 0
C1561 w_9208_4512# a_9671_5727# 0
C1562 a_4627_12141# a_4637_10577# 0
C1563 a_7815_2035# sky130_fd_sc_hd__mux4_1_0.A2 0.00297f
C1564 VGND a_11595_5467# 0.01545f
C1565 a_20384_16179# sky130_fd_sc_hd__mux4_1_0.A0 0.07865f
C1566 a_9597_13793# VDPWR 0.37502f
C1567 a_3229_5051# VGND 0.67714f
C1568 a_8566_1779# VGND 0
C1569 a_4183_1787# VGND 0.0153f
C1570 a_9801_12841# w_10872_13125# 0.05199f
C1571 a_12509_4593# a_12994_4589# 0.07537f
C1572 a_10813_13753# a_11049_14719# 0
C1573 a_9865_15329# a_9725_14509# 0
C1574 VDPWR a_24407_14651# 0.00288f
C1575 a_9865_15329# w_9402_14723# 0.00599f
C1576 VGND w_10674_14933# 0.0161f
C1577 a_10569_1777# w_9138_1692# 0.02026f
C1578 VGND a_7635_5405# 0.00305f
C1579 a_3199_1791# a_4546_1787# 0.08907f
C1580 a_18742_16187# a_19510_16177# 0.1036f
C1581 a_9549_13091# a_4915_10549# 0
C1582 a_9699_4853# a_9671_5727# 0.00177f
C1583 a_4505_13107# a_4513_14775# 0
C1584 a_6944_13645# a_6389_13769# 0.00183f
C1585 VDPWR a_14297_5463# 1.06327f
C1586 a_7815_2035# VGND 1.2f
C1587 a_4837_16089# VDPWR 1.09775f
C1588 a_15255_4841# a_15281_5459# 0
C1589 a_15644_5825# a_15281_5825# 0.00847f
C1590 sky130_fd_sc_hd__mux4_1_0.A1 a_11597_15219# 0
C1591 w_16764_4814# a_16167_5459# 0.1118f
C1592 a_6944_13645# a_4849_11293# 0
C1593 a_4837_16089# a_6862_13645# 0
C1594 a_12509_4593# VDPWR 1.05267f
C1595 a_9671_5727# a_9557_5837# 0
C1596 a_7845_5295# w_9180_5386# 0
C1597 a_4839_12857# a_6127_13769# 0.00253f
C1598 a_18742_16187# w_20196_16393# 0
C1599 a_24234_14385# a_24774_14701# 0.17579f
C1600 a_4546_1787# a_5069_1787# 0
C1601 a_9865_15329# a_9875_13765# 0.1161f
C1602 a_9280_5471# w_9180_5386# 0.01793f
C1603 a_10450_4963# VGND 0.00221f
C1604 a_9467_13091# a_11291_12911# 0
C1605 a_2175_5417# VDPWR 0
C1606 a_10813_13753# a_10895_13753# 0.00578f
C1607 a_11331_5833# a_11595_5833# 0
C1608 VGND a_15113_5459# 0
C1609 a_11351_13753# a_9875_13765# 0
C1610 a_3199_1791# a_4129_2043# 0.21188f
C1611 a_3919_1787# a_3790_1761# 0.00758f
C1612 VDPWR w_9180_5386# 0.52056f
C1613 w_12866_5378# a_11541_5723# 0
C1614 a_2175_5417# a_1950_5025# 0.00559f
C1615 ua[0] a_24234_14385# 0
C1616 a_15672_4951# a_16195_4585# 0
C1617 a_1898_5051# a_2079_5417# 0
C1618 a_10639_4597# a_8785_5039# 0.03363f
C1619 w_4528_15559# a_6629_15387# 0
C1620 a_4595_14775# a_4903_15345# 0
C1621 a_5945_2039# a_6696_1783# 0.00682f
C1622 a_9671_5727# w_11050_5382# 0
C1623 a_5069_1787# a_6885_1783# 0
C1624 a_8596_5405# a_7845_5295# 0.00696f
C1625 a_10380_2143# sky130_fd_sc_hd__mux4_1_0.A2 0
C1626 a_14864_4585# a_14888_5433# 0
C1627 a_10771_14747# a_11049_14719# 0.1109f
C1628 w_11718_13593# a_9799_16073# 0
C1629 w_5712_14949# a_6087_14735# 0.02211f
C1630 a_5069_1787# a_4129_2043# 0.13724f
C1631 VGND a_4595_14775# 0.00172f
C1632 a_11597_15219# a_9799_16073# 0.232f
C1633 a_4847_14525# a_7173_15235# 0
C1634 VDPWR w_11718_13593# 0.08767f
C1635 a_13243_5829# VDPWR 0
C1636 VDPWR a_11597_15219# 0.3359f
C1637 ui_in[0] a_24774_14701# 0.02524f
C1638 a_7424_1779# a_6885_1783# 0.0725f
C1639 w_9392_17212# sky130_fd_sc_hd__mux4_1_0.A1 0.05602f
C1640 a_9801_12841# a_9725_14509# 0
C1641 a_11906_13629# a_12075_13379# 0
C1642 a_8596_5405# VDPWR 0
C1643 a_9801_12841# w_9402_14723# 0.00408f
C1644 a_4913_13781# w_4538_13995# 0.01958f
C1645 a_14846_1739# VDPWR 0.29469f
C1646 a_3010_2157# a_2187_1765# 0
C1647 VGND a_10422_5837# 0.00262f
C1648 a_7899_5039# a_7845_5295# 0.00386f
C1649 w_9394_13055# a_9477_11527# 0
C1650 a_3199_1791# a_4015_1787# 0
C1651 a_10380_2143# VGND 0.00244f
C1652 a_9877_10533# a_4915_10549# 0.00316f
C1653 a_15239_2131# w_14694_1680# 0
C1654 a_5069_1787# a_5831_1783# 0
C1655 a_9699_4853# a_10450_4597# 0.00682f
C1656 VDPWR a_12809_13987# 0
C1657 w_11078_4508# a_11230_4567# 0.05213f
C1658 VDPWR ua[6] 0
C1659 a_24234_14385# sky130_fd_sc_hd__mux4_1_0.A0 0
C1660 ui_in[0] ua[0] 0.32623f
C1661 a_13018_5437# VGND 0.42749f
C1662 a_23731_14309# a_23511_14701# 0.00549f
C1663 a_10813_13753# a_10771_14747# 0
C1664 a_7899_5039# VDPWR 0.1761f
C1665 a_6885_1783# a_6696_2149# 0
C1666 a_14794_1765# VDPWR 0.07423f
C1667 a_4045_5047# VDPWR 0
C1668 a_9332_5445# w_9180_5386# 0.05213f
C1669 a_9801_12841# a_9875_13765# 0.44871f
C1670 VDPWR a_5099_5047# 1.05308f
C1671 sky130_fd_sc_hd__mux4_1_0.A2 a_7701_2145# 0
C1672 a_5945_2039# VDPWR 0.34532f
C1673 a_9727_11277# VDPWR 0.00377f
C1674 a_9461_5471# sky130_fd_sc_hd__mux4_1_0.A3 0
C1675 VDPWR a_9629_2033# 0.34514f
C1676 a_9461_5837# sky130_fd_sc_hd__mux4_1_0.A3 0
C1677 a_6911_15235# a_7173_15235# 0
C1678 a_12713_13987# a_12075_13379# 0.00226f
C1679 VGND a_11019_12911# 0.00238f
C1680 VDPWR a_6389_13769# 0.38708f
C1681 a_15071_1765# a_15185_2021# 0
C1682 VDPWR a_4576_5047# 0.20634f
C1683 a_6362_1783# w_5454_1698# 0.01154f
C1684 sky130_fd_sc_hd__mux4_1_0.A1 a_19510_16177# 0
C1685 a_15602_1765# a_14255_1769# 0.08907f
C1686 a_2217_5025# a_2706_5051# 0.08994f
C1687 a_15255_4841# a_15281_5825# 0
C1688 a_5765_5043# a_5636_5017# 0.00758f
C1689 a_10046_1777# a_8755_1779# 0.08907f
C1690 a_15672_4951# a_14297_5463# 0
C1691 a_9727_11527# VGND 0.02702f
C1692 VGND a_8262_5405# 0.18713f
C1693 a_6862_13645# a_6389_13769# 0.24537f
C1694 a_4837_16089# a_6635_15235# 0.232f
C1695 a_4903_15345# a_5933_13769# 0.0035f
C1696 a_4847_14525# a_4513_14775# 0.1679f
C1697 a_4839_12857# a_6087_14735# 0.02474f
C1698 w_14736_5374# a_15227_5715# 0.10454f
C1699 w_9392_17212# VDPWR 0.0708f
C1700 a_6392_5409# VGND 0.18646f
C1701 VDPWR a_4849_11293# 0.42529f
C1702 a_9673_15357# VDPWR 0.00333f
C1703 a_14946_4905# a_13271_4955# 0
C1704 a_8113_13753# a_6629_15387# 0.03523f
C1705 a_13732_1769# sky130_fd_sc_hd__mux4_1_0.A2 0
C1706 a_4159_5303# a_4213_5047# 0.00386f
C1707 VGND a_7701_2145# 0.00231f
C1708 w_5786_13983# a_7113_13395# 0
C1709 a_9597_13793# a_4915_10549# 0.00124f
C1710 a_13385_4845# a_13802_4955# 0.06611f
C1711 a_7869_1779# a_7605_1779# 0
C1712 sky130_fd_sc_hd__mux4_1_0.A2 a_2187_1765# 0.11803f
C1713 VGND a_5933_13769# 0.00382f
C1714 a_9801_12841# w_10868_12105# 0.00131f
C1715 a_6862_13645# a_4849_11293# 0
C1716 a_9360_4571# a_9489_4597# 0.00758f
C1717 ui_in[0] sky130_fd_sc_hd__mux4_1_0.A0 0.02204f
C1718 w_14736_5374# sky130_fd_sc_hd__mux4_1_0.A3 0.00647f
C1719 a_11455_4593# sky130_fd_sc_hd__mux4_1_0.A2 0
C1720 a_9867_12097# a_9799_16073# 0
C1721 a_13385_4845# a_13411_5463# 0
C1722 a_9599_10561# a_9877_10533# 0.1296f
C1723 a_5999_2149# a_5735_2149# 0
C1724 w_5484_4958# a_5099_5047# 0.25047f
C1725 a_2289_5307# w_3668_4962# 0
C1726 a_10088_5471# a_9725_5471# 0.00985f
C1727 a_4213_5047# a_3949_5047# 0
C1728 a_4635_13809# a_4513_14775# 0.00144f
C1729 a_14946_4905# a_15227_5715# 0.04605f
C1730 VDPWR a_9867_12097# 0.28921f
C1731 a_16195_4585# a_14325_4589# 0.00122f
C1732 VGND a_2079_5417# 0.00311f
C1733 a_10569_1777# sky130_fd_sc_hd__mux4_1_0.A2 0.00267f
C1734 a_13018_5437# w_12894_4504# 0
C1735 VDPWR a_7669_14003# 0.082f
C1736 a_6915_5043# a_7899_5039# 0.08312f
C1737 a_7113_13395# a_4903_15345# 0
C1738 VDPWR w_17066_16401# 0.07225f
C1739 a_9465_16323# sky130_fd_sc_hd__mux4_1_0.A1 0
C1740 a_12292_5833# VGND 0.00291f
C1741 a_13732_1769# VGND 0.01325f
C1742 a_11160_1747# a_11385_2139# 0.00559f
C1743 sky130_fd_sc_hd__mux4_1_0.A1 sky130_fd_sc_hd__mux4_1_0.A3 0.00503f
C1744 a_6915_5043# a_5099_5047# 0
C1745 a_4837_16089# a_4915_10549# 0.01618f
C1746 a_9475_14759# a_9725_14509# 0.00723f
C1747 a_10639_4597# a_11541_5723# 0
C1748 a_9801_12841# a_9717_12841# 0.00208f
C1749 a_6862_13645# a_7669_14003# 0
C1750 a_9475_14759# w_9402_14723# 0.06993f
C1751 a_14297_5463# a_13357_5719# 0.13962f
C1752 VGND a_2187_1765# 1.11393f
C1753 a_14946_4905# sky130_fd_sc_hd__mux4_1_0.A3 0.01569f
C1754 a_7113_13395# VGND 0.35166f
C1755 a_4755_13107# a_4849_11293# 0
C1756 a_11541_5723# a_11595_5467# 0.00386f
C1757 a_11160_1747# a_11553_1773# 0.02283f
C1758 a_13018_5437# a_8785_5039# 0
C1759 a_24241_14651# sky130_fd_sc_hd__mux4_1_0.VPB 0.0237f
C1760 VDPWR a_19510_16177# 0.26197f
C1761 a_16486_16197# w_16298_16411# 0.02625f
C1762 w_3638_1702# a_3790_1761# 0.05213f
C1763 a_9557_14759# a_9865_15329# 0
C1764 a_8755_1779# a_9238_1777# 0.07352f
C1765 a_12509_4593# a_13357_5719# 0
C1766 a_5851_13769# a_5933_13769# 0.00578f
C1767 a_10569_1777# VGND 0.6772f
C1768 VDPWR a_13271_4955# 0
C1769 a_4503_16339# a_4847_14525# 0
C1770 a_12994_4589# sky130_fd_sc_hd__mux4_1_0.A3 0
C1771 a_14946_4905# w_14764_4500# 0.28173f
C1772 a_11623_4959# w_11078_4508# 0
C1773 a_14946_4905# a_13046_4563# 0
C1774 a_9475_14759# a_9875_13765# 0
C1775 a_11427_5833# sky130_fd_sc_hd__mux4_1_0.A3 0
C1776 a_9877_10533# a_12713_13987# 0
C1777 a_4839_12857# a_4505_13107# 0.16952f
C1778 a_11986_4593# a_11569_4849# 0.03016f
C1779 a_6089_11935# a_4849_11293# 0
C1780 a_7845_5295# sky130_fd_sc_hd__mux4_1_0.A3 0.00297f
C1781 w_20196_16393# VDPWR 0.07122f
C1782 a_12481_5467# w_12866_5378# 0.25012f
C1783 a_5999_1783# a_2187_1765# 0
C1784 a_14836_5459# a_14297_5463# 0.0725f
C1785 a_11499_2029# a_11160_1747# 0.04737f
C1786 a_9280_5471# sky130_fd_sc_hd__mux4_1_0.A3 0.00331f
C1787 a_24318_14385# a_24241_14651# 0.01352f
C1788 VDPWR a_15227_5715# 0.32967f
C1789 a_2706_5417# VDPWR 0.01961f
C1790 a_4905_12113# w_5906_12121# 0.08119f
C1791 w_11078_4508# a_11623_4593# 0.01092f
C1792 a_5851_13769# a_7113_13395# 0
C1793 a_24962_14701# sky130_fd_sc_hd__mux4_1_0.A2 0.00234f
C1794 a_14846_1739# a_14975_2131# 0.00792f
C1795 w_4442_11507# a_4839_12857# 0
C1796 a_9465_16323# a_9799_16073# 0.16891f
C1797 a_4546_2153# VGND 0.18648f
C1798 uio_in[5] uio_in[4] 0.03102f
C1799 a_9477_11527# w_9502_10747# 0.0035f
C1800 a_12994_4589# a_13046_4563# 0.1439f
C1801 VDPWR w_9138_1692# 0.51534f
C1802 a_6021_13769# a_4839_12857# 0
C1803 a_9465_16323# VDPWR 0.3941f
C1804 VDPWR sky130_fd_sc_hd__mux4_1_0.A3 0.3547f
C1805 a_9811_11277# a_11089_13753# 0
C1806 a_11359_4959# VDPWR 0
C1807 ui_in[1] a_24774_14701# 0.63083f
C1808 a_11569_4849# a_12320_4593# 0.00682f
C1809 a_18742_16187# VGND 0.25574f
C1810 a_17125_5265# a_16167_5459# 0.00576f
C1811 w_9208_4512# a_9753_4963# 0
C1812 VDPWR w_4432_13071# 0.16326f
C1813 a_9489_4597# sky130_fd_sc_hd__mux4_1_0.A2 0
C1814 a_16871_4938# sky130_fd_sc_hd__mux4_1_0.A3 0.00367f
C1815 a_5636_5017# a_2217_5025# 0.0021f
C1816 a_13243_5829# a_13357_5719# 0
C1817 a_13315_2025# w_14694_1680# 0
C1818 a_14794_1765# a_14975_2131# 0
C1819 sky130_fd_sc_hd__mux4_1_0.A1 a_11243_11891# 0.00295f
C1820 a_14325_4589# a_14297_5463# 0.00251f
C1821 a_5975_5299# a_2217_5025# 0
C1822 w_10674_14933# a_12135_15219# 0
C1823 VGND a_24962_14701# 0.18885f
C1824 w_6044_2758# sky130_fd_sc_hd__mux4_1_0.A2 0.05211f
C1825 a_4721_13809# a_4839_12857# 0
C1826 a_5606_1757# VGND 0.40141f
C1827 a_4765_11543# a_4505_13107# 0
C1828 ua[0] ui_in[1] 0.47781f
C1829 VDPWR w_14764_4500# 0.52659f
C1830 a_3199_1791# a_3919_1787# 0
C1831 w_5906_12121# a_5975_12927# 0
C1832 VDPWR a_13046_4563# 0.29743f
C1833 a_9699_4853# a_9753_4963# 0.03622f
C1834 a_3949_5413# VDPWR 0
C1835 a_12509_4593# a_14325_4589# 0
C1836 VGND a_9489_4597# 0
C1837 a_4765_11543# w_4442_11507# 0.01327f
C1838 a_4847_14525# w_5712_14949# 0.00381f
C1839 a_9557_14759# a_9801_12841# 0
C1840 a_9727_11277# a_4915_10549# 0
C1841 a_11595_5833# a_10639_4597# 0
C1842 a_4755_13107# w_4432_13071# 0.01327f
C1843 a_15017_5825# sky130_fd_sc_hd__mux4_1_0.A3 0
C1844 w_5484_4958# sky130_fd_sc_hd__mux4_1_0.A3 0.00188f
C1845 uio_oe[4] uio_oe[5] 0.03102f
C1846 VGND w_6044_2758# 0.02955f
C1847 w_1768_1706# a_2313_1791# 0.01092f
C1848 ui_in[0] a_24234_14385# 0.28579f
C1849 a_23677_14335# VDPWR 0
C1850 a_4915_10549# a_6389_13769# 0.00254f
C1851 a_9360_4571# a_7845_5295# 0
C1852 a_15644_5459# a_16167_5459# 0
C1853 a_2217_5025# w_1798_4966# 0.25023f
C1854 a_5606_1757# a_5999_1783# 0.02283f
C1855 a_6915_5043# sky130_fd_sc_hd__mux4_1_0.A3 0.00267f
C1856 a_11160_1747# w_11008_1688# 0.05213f
C1857 a_3229_5051# a_4213_5047# 0.08312f
C1858 a_10813_13753# w_9500_13979# 0
C1859 a_9332_5445# sky130_fd_sc_hd__mux4_1_0.A3 0.00451f
C1860 a_4849_11293# a_4915_10549# 0.00639f
C1861 VDPWR a_10611_5471# 1.06898f
C1862 a_6944_13645# VGND 0
C1863 a_13018_5437# a_11541_5723# 0.00492f
C1864 a_3949_5413# a_3768_5047# 0
C1865 a_8232_1779# VDPWR 0.20639f
C1866 a_9461_5471# VGND 0
C1867 ui_in[1] sky130_fd_sc_hd__mux4_1_0.A0 0.06787f
C1868 a_9360_4571# VDPWR 0.39467f
C1869 a_9461_5837# VGND 0.00346f
C1870 VDPWR a_11243_11891# 0.21318f
C1871 a_1898_5051# VDPWR 0.08401f
C1872 a_9865_15329# a_11049_14719# 0
C1873 a_23511_14335# sky130_fd_sc_hd__mux4_1_0.VPB 0.00324f
C1874 a_11160_1747# a_11385_1773# 0.00487f
C1875 a_10965_11919# a_9799_16073# 0
C1876 a_9867_12097# a_4915_10549# 0.00417f
C1877 a_1898_5051# a_1950_5025# 0.1439f
C1878 w_7604_13967# a_8113_13753# 0.01891f
C1879 a_4915_10549# a_7669_14003# 0.07457f
C1880 uo_out[5] uo_out[4] 0.03102f
C1881 sky130_fd_sc_hd__mux4_1_0.A3 a_11986_4959# 0
C1882 VDPWR a_10965_11919# 0.1599f
C1883 a_11351_13753# a_11049_14719# 0.00427f
C1884 a_4913_13781# a_5933_13769# 0
C1885 a_3229_5051# a_3040_5417# 0
C1886 VDPWR a_3010_2157# 0
C1887 a_11455_4959# sky130_fd_sc_hd__mux4_1_0.A3 0
C1888 a_15255_4841# a_15672_4585# 0.03016f
C1889 a_4587_13107# a_4849_11293# 0
C1890 a_6696_1783# sky130_fd_sc_hd__mux4_1_0.A2 0
C1891 a_14946_4905# sky130_fd_sc_hd__mux4_1_0.A2 0
C1892 a_7701_1779# a_6885_1783# 0
C1893 a_13105_1769# sky130_fd_sc_hd__mux4_1_0.A2 0
C1894 a_4839_12857# a_4847_14525# 0.20053f
C1895 a_9465_16323# a_9547_16323# 0.00641f
C1896 w_14736_5374# VGND 0.29321f
C1897 a_10813_13753# a_9865_15329# 0.16764f
C1898 a_15672_4951# sky130_fd_sc_hd__mux4_1_0.A3 0
C1899 w_4530_12327# a_4849_11293# 0.00145f
C1900 a_9865_15329# a_10895_13753# 0.0035f
C1901 a_15239_1765# a_15185_2021# 0.00386f
C1902 w_4538_13995# a_4513_14775# 0.0035f
C1903 VGND sky130_fd_sc_hd__mux4_1_0.A1 0.7644f
C1904 a_12994_4589# sky130_fd_sc_hd__mux4_1_0.A2 0
C1905 a_1920_1765# a_2313_1791# 0.02283f
C1906 VDPWR a_11427_5467# 0.00102f
C1907 VGND a_6696_1783# 0
C1908 a_4635_13809# a_4839_12857# 0.00246f
C1909 a_10813_13753# a_11351_13753# 0.07901f
C1910 a_7424_1779# a_7476_1753# 0.1439f
C1911 a_5945_2039# a_5831_2149# 0
C1912 a_14946_4905# VGND 0.17745f
C1913 a_9557_14759# a_9475_14759# 0.00641f
C1914 a_11351_13753# a_10895_13753# 0
C1915 a_13105_1769# VGND 0
C1916 a_12292_5833# a_11541_5723# 0.00696f
C1917 a_9809_14509# a_9799_16073# 0.46421f
C1918 uo_out[1] uo_out[2] 0.03102f
C1919 a_9360_4571# a_9332_5445# 0
C1920 a_4905_12113# a_4839_12857# 0.04364f
C1921 a_5069_1787# a_6362_2149# 0.03325f
C1922 a_9671_5727# w_9180_5386# 0.10454f
C1923 a_4576_5413# a_4213_5413# 0.00847f
C1924 a_9809_14509# VDPWR 0.3635f
C1925 VDPWR a_2175_5051# 0.00105f
C1926 a_5975_5299# w_7354_4954# 0
C1927 a_15672_4951# w_14764_4500# 0.00139f
C1928 a_12509_4593# a_13802_4589# 0.08907f
C1929 a_2175_5051# a_1950_5025# 0.00487f
C1930 w_5786_13983# VDPWR 0.0898f
C1931 a_9589_12125# w_9404_11491# 0.00155f
C1932 a_12994_4589# VGND 0.08826f
C1933 a_5975_5299# a_6726_5409# 0.00696f
C1934 a_4183_1787# a_4546_1787# 0.00985f
C1935 VDPWR sky130_fd_sc_hd__mux4_1_0.A2 0.2927f
C1936 a_10611_5471# a_11986_4959# 0
C1937 a_10937_12911# a_9811_11277# 0.18651f
C1938 a_11427_5833# VGND 0.00241f
C1939 a_9699_4853# a_9725_5837# 0
C1940 a_2259_2047# w_3638_1702# 0
C1941 a_9801_12841# a_11049_14719# 0.02474f
C1942 a_11767_15219# a_9799_16073# 0
C1943 VGND a_7845_5295# 1.20783f
C1944 a_6281_11907# a_4905_12113# 0.03573f
C1945 a_13357_5719# sky130_fd_sc_hd__mux4_1_0.A3 0.00759f
C1946 VDPWR a_6003_11935# 0.1599f
C1947 a_3199_1791# w_3638_1702# 0.25055f
C1948 a_4515_11543# a_4849_11293# 0.16782f
C1949 a_9280_5471# VGND 0.12844f
C1950 a_15602_2131# w_14694_1680# 0.00139f
C1951 VDPWR a_11767_15219# 0.00151f
C1952 a_24318_14385# sky130_fd_sc_hd__mux4_1_0.VPB 0.00426f
C1953 VDPWR a_4903_15345# 0.24554f
C1954 a_5975_12927# a_4839_12857# 0.30276f
C1955 a_9875_13765# w_10674_14933# 0
C1956 a_1920_1765# a_2049_2157# 0.00792f
C1957 a_9699_4853# w_11078_4508# 0
C1958 VGND a_9799_16073# 0.68227f
C1959 w_16298_16411# sky130_fd_sc_hd__mux4_1_0.A0 0.07239f
C1960 a_9811_11277# a_12075_13379# 0.00118f
C1961 a_9725_5837# a_9557_5837# 0
C1962 a_9549_13091# a_9811_11277# 0
C1963 a_6862_13645# a_4903_15345# 0
C1964 a_12966_5463# w_11050_5382# 0.00227f
C1965 VDPWR VGND 63.55989f
C1966 w_14736_5374# a_8785_5039# 0.00355f
C1967 w_11532_15433# a_8113_13753# 0.097f
C1968 w_5910_13141# a_4839_12857# 0.05199f
C1969 a_9865_15329# a_10771_14747# 0.0039f
C1970 a_13046_4563# a_13357_5719# 0
C1971 a_5069_1787# w_3638_1702# 0.01972f
C1972 a_15141_4585# a_15309_4585# 0
C1973 a_14946_4905# w_12894_4504# 0.00104f
C1974 a_9715_16323# a_9799_16073# 0.07445f
C1975 a_9717_13091# VDPWR 0.31944f
C1976 a_12509_4593# a_13175_4589# 0
C1977 a_13018_5437# a_13147_5463# 0.00758f
C1978 a_3820_5021# w_1798_4966# 0
C1979 a_2259_2047# a_3790_1761# 0.00446f
C1980 a_16871_4938# VGND 0.1106f
C1981 VGND a_6862_13645# 0.13594f
C1982 uio_in[3] uio_in[4] 0.03102f
C1983 VGND a_1950_5025# 0.40871f
C1984 a_15113_5825# a_14888_5433# 0.00559f
C1985 a_4183_1787# a_4129_2043# 0.00386f
C1986 ui_in[1] a_24234_14385# 0.34741f
C1987 a_3199_1791# a_3790_1761# 0.11887f
C1988 a_14136_4589# VDPWR 0
C1989 VDPWR a_4637_10577# 0.36832f
C1990 VDPWR a_9715_16323# 0.32305f
C1991 a_10813_13753# a_9801_12841# 0.13074f
C1992 a_6281_11907# a_5975_12927# 0
C1993 a_14836_5459# sky130_fd_sc_hd__mux4_1_0.A3 0.003f
C1994 a_9801_12841# a_10895_13753# 0
C1995 a_5999_2149# a_6362_2149# 0.00847f
C1996 a_7815_2035# a_6885_1783# 0.21188f
C1997 a_14946_4905# a_8785_5039# 0.56407f
C1998 a_13315_2025# w_12824_1684# 0.10454f
C1999 a_12994_4589# w_12894_4504# 0.01793f
C2000 a_13732_2135# sky130_fd_sc_hd__mux4_1_0.A2 0
C2001 a_5735_1783# VGND 0
C2002 a_15239_2131# a_15602_2131# 0.00847f
C2003 a_6281_11907# w_5910_13141# 0
C2004 a_12631_13987# sky130_fd_sc_hd__mux4_1_0.A1 0.10369f
C2005 a_14325_4589# a_15227_5715# 0
C2006 a_10813_13753# w_12566_13951# 0
C2007 w_14736_5374# a_14916_4559# 0.00104f
C2008 a_4755_13107# VGND 0.02544f
C2009 a_5999_1783# VDPWR 0.17397f
C2010 a_13385_4845# a_13271_4589# 0
C2011 a_11289_1773# a_10569_1777# 0
C2012 a_11160_1747# a_11108_1773# 0.1439f
C2013 VGND a_3768_5047# 0.08661f
C2014 a_10937_12911# a_11824_13629# 0
C2015 a_11569_4849# a_11230_4567# 0.04737f
C2016 a_5851_13769# VDPWR 0.3558f
C2017 a_15017_5825# VGND 0.00305f
C2018 a_11958_5833# sky130_fd_sc_hd__mux4_1_0.A3 0.00158f
C2019 w_5484_4958# VGND 0.29342f
C2020 a_6089_11935# a_6003_11935# 0.00658f
C2021 a_4627_12141# w_5906_12121# 0
C2022 a_12481_5467# a_13018_5437# 0.11552f
C2023 a_14325_4589# sky130_fd_sc_hd__mux4_1_0.A3 0
C2024 a_12976_1743# a_13315_2025# 0.04737f
C2025 a_15281_5459# a_14297_5463# 0.08312f
C2026 a_5851_13769# a_6862_13645# 0
C2027 a_12439_1773# sky130_fd_sc_hd__mux4_1_0.A2 0.0028f
C2028 a_12976_1743# w_12824_1684# 0.05213f
C2029 a_9799_16073# a_10857_14747# 0
C2030 a_4183_1787# a_4015_1787# 0
C2031 a_7845_5295# a_8785_5039# 0.13855f
C2032 a_9589_12125# w_9500_13979# 0
C2033 a_6915_5043# VGND 0.68138f
C2034 a_10422_5471# sky130_fd_sc_hd__mux4_1_0.A3 0
C2035 a_13732_2135# VGND 0.18636f
C2036 a_14946_4905# a_14916_4559# 0.38909f
C2037 VDPWR w_12894_4504# 0.52899f
C2038 a_9280_5471# a_8785_5039# 0
C2039 a_9332_5445# VGND 0.51815f
C2040 a_13315_2025# a_14066_1769# 0.00682f
C2041 ui_in[0] ui_in[1] 5.47082f
C2042 a_11289_2139# VDPWR 0
C2043 VDPWR a_10857_14747# 0
C2044 a_11824_13629# a_12075_13379# 0.10945f
C2045 a_9865_15329# w_9392_16287# 0
C2046 VDPWR a_6057_12927# 0
C2047 a_4837_16089# w_4528_15559# 0.00251f
C2048 a_6089_11935# VGND 0.00568f
C2049 a_5999_1783# a_5735_1783# 0
C2050 a_9475_14759# a_11049_14719# 0
C2051 a_23511_14701# sky130_fd_sc_hd__mux4_1_0.A0 0.09907f
C2052 a_14325_4589# w_14764_4500# 0.25055f
C2053 uio_in[2] uio_in[3] 0.03102f
C2054 sky130_fd_sc_hd__mux4_1_0.A3 a_9308_4597# 0
C2055 sky130_fd_sc_hd__mux4_1_0.A1 a_23677_14701# 0
C2056 a_13018_5437# a_13243_5463# 0.00487f
C2057 uo_out[7] uio_out[0] 0.03102f
C2058 a_4515_11543# w_4432_13071# 0
C2059 a_14946_4905# a_17346_5265# 0
C2060 a_21506_16181# w_21318_16395# 0.02625f
C2061 VDPWR a_8785_5039# 2.23739f
C2062 VDPWR a_10046_2143# 0.01966f
C2063 a_12439_1773# VGND 0.67525f
C2064 w_11532_15433# a_11824_13629# 0
C2065 a_12250_2139# sky130_fd_sc_hd__mux4_1_0.A2 0
C2066 VGND a_2676_1791# 0.01464f
C2067 a_9877_10533# a_9811_11277# 0.00639f
C2068 a_9801_12841# a_10771_14747# 0.21988f
C2069 a_16871_4938# a_8785_5039# 0.25154f
C2070 a_14066_2135# a_14255_1769# 0
C2071 a_12631_13987# VDPWR 0.07848f
C2072 VGND a_11986_4959# 0.18607f
C2073 w_4440_14739# a_4625_15373# 0.00155f
C2074 a_6281_11907# a_7847_14003# 0.00264f
C2075 a_9811_11277# a_9725_14759# 0
C2076 a_11455_4959# VGND 0.00209f
C2077 a_4595_14775# a_4513_14775# 0.00641f
C2078 a_15936_1765# VDPWR 0
C2079 a_14975_2131# sky130_fd_sc_hd__mux4_1_0.A2 0
C2080 a_6635_15235# a_4903_15345# 0
C2081 a_4837_16089# w_6756_13609# 0
C2082 VGND a_9547_16323# 0.00117f
C2083 a_11958_5833# a_10611_5471# 0.03325f
C2084 a_11986_4593# a_11623_4593# 0.00985f
C2085 a_6629_15387# w_6570_15449# 0.097f
C2086 a_14916_4559# VDPWR 0.31865f
C2087 a_9809_14509# a_4915_10549# 0
C2088 a_12481_5467# a_12292_5833# 0
C2089 a_12250_2139# VGND 0.00244f
C2090 a_7899_5039# a_7506_5013# 0.02283f
C2091 a_15978_5459# a_15227_5715# 0.00682f
C2092 a_9290_1751# a_9419_2143# 0.00792f
C2093 a_2313_2157# VGND 0.19866f
C2094 a_11906_13629# a_11243_11891# 0
C2095 a_11359_4593# sky130_fd_sc_hd__mux4_1_0.A2 0
C2096 VGND a_6635_15235# 0.13063f
C2097 uio_out[3] uio_out[2] 0.03102f
C2098 sky130_fd_sc_hd__mux4_1_0.A3 a_11331_5467# 0
C2099 a_9629_2033# w_11008_1688# 0
C2100 a_4159_5303# a_4910_5413# 0.00696f
C2101 a_9597_13793# a_8113_13753# 0.00382f
C2102 w_5786_13983# a_4915_10549# 0
C2103 a_15672_4951# VGND 0
C2104 a_15978_5459# sky130_fd_sc_hd__mux4_1_0.A3 0
C2105 VDPWR a_17346_5265# 0
C2106 a_15185_2021# w_14694_1680# 0.10454f
C2107 a_5861_5043# a_5099_5047# 0
C2108 a_3919_2153# a_3790_1761# 0.00792f
C2109 VDPWR a_23677_14701# 0.18463f
C2110 a_6003_11935# a_4915_10549# 0
C2111 a_14975_2131# VGND 0.00305f
C2112 a_13439_4589# a_13271_4589# 0
C2113 a_6915_5043# a_8785_5039# 0
C2114 a_4839_12857# w_4538_13995# 0.00445f
C2115 a_9671_5727# sky130_fd_sc_hd__mux4_1_0.A3 0.00739f
C2116 a_9597_13793# a_9811_11277# 0.00317f
C2117 a_3229_5051# a_2289_5307# 0.13962f
C2118 a_2175_5417# a_2343_5417# 0
C2119 a_7113_13395# a_7173_15235# 0.36868f
C2120 VDPWR a_13105_2135# 0
C2121 w_4442_11507# a_4505_13107# 0
C2122 a_9332_5445# a_8785_5039# 0
C2123 a_9360_4571# a_9308_4597# 0.1439f
C2124 a_11623_4959# a_11569_4849# 0.03622f
C2125 a_23731_14309# a_24962_14701# 0
C2126 w_9208_4512# a_10116_4597# 0.01154f
C2127 a_4546_1787# a_2187_1765# 0
C2128 a_9290_1751# w_7324_1694# 0
C2129 a_9877_10533# a_11824_13629# 0
C2130 a_12713_13987# a_11243_11891# 0.00373f
C2131 VGND a_4915_10549# 1.01177f
C2132 a_2706_5051# w_1798_4966# 0.01154f
C2133 a_11569_4849# a_11623_4593# 0.00386f
C2134 a_14297_5463# a_15281_5825# 0.04534f
C2135 a_9717_13091# a_4915_10549# 0
C2136 VGND a_13357_5719# 1.20852f
C2137 a_4637_10577# a_4915_10549# 0.1296f
C2138 uio_oe[6] uio_oe[5] 0.03102f
C2139 a_9699_4853# a_10116_4597# 0.03016f
C2140 a_11427_5833# a_11541_5723# 0
C2141 a_4913_13781# VDPWR 0.60287f
C2142 a_9629_2033# a_10380_1777# 0.00682f
C2143 a_15239_2131# a_15185_2021# 0.03622f
C2144 a_9475_14759# a_10771_14747# 0
C2145 a_9467_13091# a_10937_12911# 0
C2146 a_4913_13781# a_6862_13645# 0
C2147 a_7899_5039# a_7635_5039# 0
C2148 a_9801_12841# w_9404_11491# 0
C2149 a_11331_5467# a_10611_5471# 0
C2150 VGND a_4587_13107# 0.00171f
C2151 a_4847_14525# a_6087_14735# 0.3196f
C2152 sky130_fd_sc_hd__mux4_1_0.A1 a_12135_15219# 0.04463f
C2153 a_9865_15329# w_9500_13979# 0.00397f
C2154 a_3040_5051# a_2217_5025# 0
C2155 a_4129_2043# a_2187_1765# 0.00305f
C2156 w_4530_12327# a_6003_11935# 0
C2157 VDPWR a_6717_15235# 0
C2158 a_7731_5405# sky130_fd_sc_hd__mux4_1_0.A3 0
C2159 a_4627_12141# a_4839_12857# 0
C2160 VDPWR a_11541_5723# 0.33237f
C2161 a_5851_13769# a_4915_10549# 0.00193f
C2162 a_9801_12841# a_9589_12125# 0
C2163 a_7701_1779# a_7476_1753# 0.00487f
C2164 a_9685_10561# VDPWR 0.00176f
C2165 a_15672_4951# a_8785_5039# 0
C2166 a_14836_5459# VGND 0.08665f
C2167 a_9671_5727# a_10611_5471# 0.13962f
C2168 a_7869_2145# w_7324_1694# 0
C2169 a_9467_13091# a_9549_13091# 0.00641f
C2170 a_14325_4589# sky130_fd_sc_hd__mux4_1_0.A2 0
C2171 a_9360_4571# a_9671_5727# 0
C2172 w_22086_16385# VGND 0.01425f
C2173 a_5735_2149# a_2187_1765# 0
C2174 a_11597_15219# a_8113_13753# 0.1684f
C2175 w_4530_12327# VGND 0.11704f
C2176 w_6756_13609# a_6389_13769# 0.06723f
C2177 a_5831_1783# a_2187_1765# 0
C2178 a_11916_2139# a_11553_2139# 0.00847f
C2179 a_3199_1791# a_2259_2047# 0.13962f
C2180 a_9599_10561# VGND 0.24388f
C2181 a_4183_1787# a_3919_1787# 0
C2182 a_9811_11277# w_11718_13593# 0
C2183 a_7605_2145# a_7476_1753# 0.00792f
C2184 a_9559_11527# VDPWR 0.02511f
C2185 a_4627_12141# a_6281_11907# 0
C2186 w_12894_4504# a_13357_5719# 0
C2187 sky130_fd_sc_hd__mux4_1_0.A2 a_9308_4597# 0
C2188 VGND a_11958_5833# 0.1907f
C2189 w_6756_13609# a_4849_11293# 0
C2190 VGND a_11906_13629# 0
C2191 a_6911_15235# a_6087_14735# 0.00651f
C2192 a_14325_4589# VGND 0.07198f
C2193 a_17254_16187# w_19322_16391# 0
C2194 a_5975_5299# a_5636_5017# 0.04737f
C2195 a_9589_12125# w_9492_12311# 0.05631f
C2196 a_7506_5013# sky130_fd_sc_hd__mux4_1_0.A3 0.00206f
C2197 a_13046_4563# a_13175_4589# 0.00758f
C2198 a_4015_1787# a_2187_1765# 0
C2199 a_4129_2043# a_4546_2153# 0.06611f
C2200 a_9475_14759# w_9392_16287# 0
C2201 a_12135_15219# a_9799_16073# 0.04819f
C2202 a_4627_12141# a_4765_11543# 0
C2203 a_4585_16339# VDPWR 0.0251f
C2204 a_13357_5719# a_8785_5039# 0
C2205 a_3199_1791# a_5069_1787# 0
C2206 VGND a_10422_5471# 0
C2207 a_5831_2149# VGND 0.00231f
C2208 VDPWR a_12135_15219# 0.55326f
C2209 ui_in[0] a_23511_14701# 0.00322f
C2210 a_11331_5833# a_11202_5441# 0.00792f
C2211 w_6756_13609# a_7669_14003# 0
C2212 a_5895_14763# VDPWR 0
C2213 a_4515_11543# VGND 0.29765f
C2214 a_4847_14525# a_4505_13107# 0
C2215 a_9867_12097# a_9675_12125# 0
C2216 a_15281_5459# a_15227_5715# 0.00386f
C2217 a_9865_15329# a_11351_13753# 0
C2218 VGND a_9308_4597# 0.08793f
C2219 a_11289_1773# VDPWR 0.00117f
C2220 uio_in[7] uo_out[0] 0.03102f
C2221 a_9727_11277# a_9811_11277# 0.00206f
C2222 a_6329_12927# a_6389_13769# 0.20048f
C2223 a_4129_2043# a_5606_1757# 0.00492f
C2224 a_12713_13987# VGND 0
C2225 a_11427_5833# a_11595_5833# 0
C2226 a_11049_14719# w_10674_14933# 0.02211f
C2227 a_4515_11543# a_4637_10577# 0.00144f
C2228 a_9801_12841# w_9500_13979# 0.00445f
C2229 a_15281_5459# sky130_fd_sc_hd__mux4_1_0.A3 0
C2230 w_9392_17212# a_8113_13753# 0.00457f
C2231 a_11385_2139# sky130_fd_sc_hd__mux4_1_0.A2 0
C2232 w_10872_13125# a_9799_16073# 0
C2233 a_4635_13809# a_4505_13107# 0.00115f
C2234 a_16195_4585# a_15672_4585# 0
C2235 a_6329_12927# a_4849_11293# 0.00976f
C2236 a_5606_1757# a_5735_2149# 0.00792f
C2237 sky130_fd_sc_hd__mux4_1_0.A2 a_11553_1773# 0
C2238 a_4905_12113# a_4505_13107# 0
C2239 VDPWR w_10872_13125# 0.0888f
C2240 a_9629_2033# a_11108_1773# 0
C2241 w_11718_13593# a_11824_13629# 0.06114f
C2242 a_8755_1779# a_7815_2035# 0.13781f
C2243 a_5606_1757# a_5831_1783# 0.00487f
C2244 a_11595_5833# VDPWR 0.00668f
C2245 a_11597_15219# a_11824_13629# 0
C2246 a_4595_14775# a_4839_12857# 0
C2247 a_11958_5467# w_11050_5382# 0.01154f
C2248 a_14325_4589# w_12894_4504# 0.02026f
C2249 a_4183_2153# VGND 0.20098f
C2250 a_4213_5047# VDPWR 0.17485f
C2251 a_8113_13753# a_7669_14003# 0.10318f
C2252 a_15045_4585# sky130_fd_sc_hd__mux4_1_0.A2 0
C2253 a_4905_12113# w_4442_11507# 0.00119f
C2254 a_7815_2035# a_7476_1753# 0.04737f
C2255 a_11385_2139# VGND 0.00231f
C2256 VGND a_11331_5467# 0
C2257 a_11873_15219# a_11597_15219# 0.00119f
C2258 a_7635_5039# sky130_fd_sc_hd__mux4_1_0.A3 0
C2259 a_9360_4571# a_7506_5013# 0
C2260 a_9811_11277# a_9867_12097# 0.25265f
C2261 a_15071_1765# VDPWR 0
C2262 a_2343_5051# a_2175_5051# 0
C2263 a_7113_13395# a_7751_14003# 0.00226f
C2264 a_6717_15235# a_6635_15235# 0.00578f
C2265 a_14325_4589# a_8785_5039# 0.03312f
C2266 a_23731_14309# VDPWR 0.15203f
C2267 VGND a_11553_1773# 0.01595f
C2268 a_5861_5409# a_2217_5025# 0
C2269 a_15978_5459# VGND 0
C2270 a_2706_5417# a_2343_5417# 0.00847f
C2271 a_11499_2029# sky130_fd_sc_hd__mux4_1_0.A2 0.00294f
C2272 a_13147_5463# VDPWR 0.00103f
C2273 a_4635_13809# a_4721_13809# 0.00658f
C2274 a_9671_5727# VGND 1.46609f
C2275 a_5975_12927# a_4505_13107# 0
C2276 sky130_fd_sc_hd__mux4_1_0.A2 a_13802_4589# 0
C2277 a_11150_5467# w_11050_5382# 0.01793f
C2278 a_3040_5417# VDPWR 0
C2279 a_10937_12911# a_11091_12911# 0.00401f
C2280 a_9801_12841# a_9865_15329# 0.1369f
C2281 a_12509_4593# w_11078_4508# 0.01988f
C2282 a_9308_4597# a_8785_5039# 0
C2283 a_5069_1787# a_5999_2149# 0.04534f
C2284 a_2217_5025# a_5765_5409# 0
C2285 w_5910_13141# a_4505_13107# 0
C2286 a_9801_12841# a_11351_13753# 0.04676f
C2287 VDPWR a_9585_4963# 0
C2288 a_9725_5837# w_9180_5386# 0
C2289 a_2217_5025# a_4213_5413# 0
C2290 a_11623_4959# a_11230_4567# 0.02301f
C2291 a_11499_2029# VGND 1.19976f
C2292 a_14325_4589# a_14916_4559# 0.11887f
C2293 a_9467_13091# a_9597_13793# 0.00115f
C2294 a_13385_4845# a_14297_5463# 0
C2295 a_2343_5051# VGND 0.01592f
C2296 a_2259_2047# a_3010_1791# 0.00682f
C2297 VGND a_13802_4589# 0.01131f
C2298 a_12631_13987# a_12713_13987# 0.00695f
C2299 a_12481_5467# VDPWR 1.01592f
C2300 a_9465_16323# a_8113_13753# 0.0062f
C2301 w_12566_13951# a_11351_13753# 0
C2302 a_14946_4905# a_15017_5459# 0
C2303 a_11230_4567# a_11623_4593# 0.02283f
C2304 a_14297_5463# a_15672_4585# 0
C2305 a_9475_14759# w_9500_13979# 0.0035f
C2306 a_4183_1787# w_3638_1702# 0.01092f
C2307 a_12509_4593# a_13385_4845# 0.21149f
C2308 a_9799_16073# w_9402_14723# 0
C2309 sky130_fd_sc_hd__mux4_1_0.A2 a_13175_4589# 0
C2310 a_15227_5715# a_15281_5825# 0.03622f
C2311 VDPWR a_9725_14509# 0.00474f
C2312 a_5933_13769# a_4839_12857# 0
C2313 VDPWR w_9402_14723# 0.16205f
C2314 a_14108_5463# sky130_fd_sc_hd__mux4_1_0.A3 0
C2315 w_12866_5378# a_13774_5463# 0.01154f
C2316 a_9559_11527# a_4915_10549# 0
C2317 VDPWR a_7173_15235# 0.55471f
C2318 a_10771_14747# w_10674_14933# 0.05631f
C2319 a_9419_2143# a_9683_2143# 0
C2320 a_7731_5405# VGND 0.00235f
C2321 a_15281_5825# sky130_fd_sc_hd__mux4_1_0.A3 0.00135f
C2322 a_10450_4597# sky130_fd_sc_hd__mux4_1_0.A2 0
C2323 a_13774_5829# w_12866_5378# 0.00139f
C2324 a_13243_5463# VDPWR 0
C2325 a_9753_4963# sky130_fd_sc_hd__mux4_1_0.A3 0
C2326 w_9394_13055# a_10937_12911# 0
C2327 a_11597_15219# a_11679_15219# 0.00578f
C2328 a_4546_1787# VDPWR 0.20643f
C2329 w_11008_1688# sky130_fd_sc_hd__mux4_1_0.A2 0.00321f
C2330 a_4183_1787# a_3790_1761# 0.02283f
C2331 a_11108_1773# w_9138_1692# 0.00188f
C2332 a_9875_13765# a_9799_16073# 0.01745f
C2333 a_14946_4905# a_15045_4951# 0.0029f
C2334 a_23511_14701# ui_in[1] 0.05408f
C2335 VGND a_13175_4589# 0
C2336 a_9671_5727# a_8785_5039# 0
C2337 a_11569_4849# w_11050_5382# 0.00166f
C2338 sky130_fd_sc_hd__mux4_1_0.A3 a_6726_5043# 0
C2339 a_7113_13395# a_4839_12857# 0.00444f
C2340 a_3919_1787# a_2187_1765# 0
C2341 VDPWR a_9875_13765# 0.60287f
C2342 a_18742_16187# w_18554_16401# 0.02625f
C2343 a_11178_4593# a_11202_5441# 0
C2344 a_4635_13809# a_4847_14525# 0
C2345 sky130_fd_sc_hd__mux4_1_0.A1 a_16486_16197# 0
C2346 a_10450_4597# VGND 0
C2347 w_12894_4504# a_13802_4589# 0.01154f
C2348 VDPWR a_15017_5459# 0.00132f
C2349 ua[4] VDPWR 0.00186f
C2350 a_9599_10561# a_9685_10561# 0.00658f
C2351 a_11385_1773# sky130_fd_sc_hd__mux4_1_0.A2 0
C2352 a_4763_14775# w_4440_14739# 0.01327f
C2353 VGND a_7506_5013# 0.40201f
C2354 VGND w_11008_1688# 0.29328f
C2355 sky130_fd_sc_hd__mux4_1_0.A2 a_9419_1777# 0
C2356 a_9865_15329# a_9475_14759# 0.00566f
C2357 VDPWR a_6885_1783# 1.0518f
C2358 w_1768_1706# a_1920_1765# 0.05213f
C2359 a_11958_5833# a_11541_5723# 0.06611f
C2360 a_4627_12141# w_4540_10763# 0
C2361 a_7701_2145# a_7476_1753# 0.00559f
C2362 a_14946_4905# a_15309_4951# 0.19411f
C2363 a_6281_11907# a_7113_13395# 0.19825f
C2364 w_19322_16391# a_18128_16189# 0
C2365 a_10088_5471# w_9180_5386# 0.01154f
C2366 a_9801_12841# w_12566_13951# 0
C2367 a_4129_2043# VDPWR 0.34561f
C2368 a_5861_5043# VGND 0
C2369 w_10868_12105# a_9799_16073# 0
C2370 a_16195_4585# a_17339_4938# 0
C2371 a_4159_5303# w_3668_4962# 0.10454f
C2372 a_17125_4938# a_17339_4938# 0.00557f
C2373 a_5945_2039# a_6362_1783# 0.03016f
C2374 a_14916_4559# a_15045_4585# 0.00758f
C2375 w_10868_12105# VDPWR 0.07869f
C2376 VDPWR a_4513_14775# 0.38904f
C2377 a_10380_1777# sky130_fd_sc_hd__mux4_1_0.A2 0
C2378 VGND a_11385_1773# 0
C2379 a_6629_15387# a_4625_15373# 0
C2380 a_9683_1777# a_9290_1751# 0.02283f
C2381 VGND a_9419_1777# 0
C2382 VDPWR a_15045_4951# 0
C2383 a_9811_11277# a_11243_11891# 0.00683f
C2384 VDPWR a_5735_2149# 0
C2385 a_24962_14701# a_24774_14701# 0.10432f
C2386 a_4903_15345# w_4528_15559# 0.01828f
C2387 a_6392_5409# a_6029_5409# 0.00847f
C2388 VDPWR a_5831_1783# 0
C2389 a_15281_5459# VGND 0.01492f
C2390 a_5765_5043# a_5099_5047# 0
C2391 a_9360_4571# a_9753_4963# 0.02301f
C2392 a_12509_4593# a_13439_4589# 0.08101f
C2393 a_24152_14385# sky130_fd_sc_hd__mux4_1_0.VPB 0.00146f
C2394 a_9717_12841# VDPWR 0.00415f
C2395 VGND w_4528_15559# 0.11947f
C2396 a_9811_11277# a_10965_11919# 0.10332f
C2397 a_8755_1779# a_10569_1777# 0
C2398 VDPWR a_16486_16197# 0.25987f
C2399 VGND a_10380_1777# 0
C2400 w_4538_13995# a_4505_13107# 0
C2401 ua[0] a_24962_14701# 0.13397f
C2402 VDPWR a_4015_1787# 0
C2403 a_10639_4597# a_11202_5441# 0
C2404 a_14846_1739# a_14975_1765# 0.00758f
C2405 a_4755_13107# a_4513_14775# 0
C2406 a_3820_5021# a_4213_5413# 0.02301f
C2407 a_15602_2131# a_15185_2021# 0.06611f
C2408 VDPWR a_15309_4951# 0.00889f
C2409 a_4905_12113# a_5975_12927# 0
C2410 a_13201_2135# a_13369_2135# 0
C2411 a_12509_4593# a_13411_5829# 0
C2412 a_4576_5413# VGND 0.18649f
C2413 a_11202_5441# a_11595_5467# 0.02283f
C2414 a_24318_14385# a_24152_14385# 0.05583f
C2415 VDPWR w_5906_12121# 0.07869f
C2416 a_7635_5039# VGND 0
C2417 a_2175_5417# a_2217_5025# 0
C2418 a_12966_5463# sky130_fd_sc_hd__mux4_1_0.A3 0.00303f
C2419 a_8232_2145# w_7324_1694# 0.00139f
C2420 a_6635_15235# a_7173_15235# 0.08446f
C2421 a_4905_12113# w_5910_13141# 0
C2422 a_4503_16339# VDPWR 0.39579f
C2423 a_7815_2035# a_9238_1777# 0
C2424 a_5584_5043# w_3668_4962# 0.00227f
C2425 a_9801_12841# a_9475_14759# 0.00442f
C2426 VGND w_6756_13609# 0.01919f
C2427 a_9809_14509# a_8113_13753# 0.30331f
C2428 a_9515_1777# a_9290_1751# 0.00487f
C2429 a_7454_5039# a_7635_5405# 0
C2430 a_18742_16187# sky130_fd_sc_hd__mux4_1_0.A0 0.04617f
C2431 VGND a_9675_12125# 0.00662f
C2432 a_7731_5039# a_7845_5295# 0
C2433 a_5809_14763# w_4440_14739# 0
C2434 a_2145_1791# a_2259_2047# 0
C2435 a_11824_13629# a_11243_11891# 0.00248f
C2436 a_9467_13091# a_9867_12097# 0
C2437 a_9683_1777# a_9515_1777# 0
C2438 VGND a_2343_5417# 0.20137f
C2439 a_9809_14509# a_9811_11277# 0.00506f
C2440 a_9725_5837# sky130_fd_sc_hd__mux4_1_0.A3 0.0014f
C2441 a_18742_16187# a_20384_16179# 0
C2442 a_11595_5833# a_11958_5833# 0.00847f
C2443 a_14136_4955# VGND 0.00215f
C2444 a_12481_5467# a_13357_5719# 0.21149f
C2445 a_24962_14701# sky130_fd_sc_hd__mux4_1_0.A0 0
C2446 a_6944_13645# a_4839_12857# 0
C2447 w_9208_4512# a_11230_4567# 0
C2448 a_9725_14509# a_4915_10549# 0
C2449 VDPWR a_4753_16339# 0.32314f
C2450 a_9699_4853# a_9725_5471# 0
C2451 a_13385_4845# a_13271_4955# 0
C2452 a_4627_12141# a_4505_13107# 0.00144f
C2453 a_5554_1783# VGND 0.08664f
C2454 a_24241_14651# a_24407_14651# 0.00988f
C2455 a_4915_10549# a_7173_15235# 0.07716f
C2456 VDPWR a_7731_5039# 0
C2457 w_14736_5374# a_16167_5459# 0.02073f
C2458 sky130_fd_sc_hd__mux4_1_0.A1 a_22274_16171# 0
C2459 a_4837_16089# w_6570_15449# 0.09702f
C2460 w_11078_4508# sky130_fd_sc_hd__mux4_1_0.A3 0
C2461 a_13243_5829# a_13411_5829# 0
C2462 w_5910_13141# a_5975_12927# 0.04996f
C2463 a_10569_1777# a_11916_2139# 0.03325f
C2464 a_15239_1765# VDPWR 0.17252f
C2465 a_9877_10533# a_9477_11527# 0
C2466 uio_in[0] uio_in[1] 0.03102f
C2467 uo_out[7] uo_out[6] 0.03102f
C2468 a_15255_4841# a_16006_4951# 0.00696f
C2469 a_4880_1787# a_2187_1765# 0
C2470 w_3638_1702# a_2187_1765# 0.00351f
C2471 a_4627_12141# w_4442_11507# 0.00155f
C2472 a_4763_14775# a_4625_15373# 0
C2473 VGND a_8113_13753# 0.15767f
C2474 a_5851_13769# w_6756_13609# 0.00132f
C2475 a_9699_4853# a_11230_4567# 0.00446f
C2476 a_13243_5463# a_13357_5719# 0
C2477 a_9465_16323# w_9490_15543# 0.0035f
C2478 VDPWR a_7751_14003# 0
C2479 w_9394_13055# a_9597_13793# 0.00101f
C2480 w_1768_1706# a_2676_2157# 0.00139f
C2481 a_6281_11907# a_6944_13645# 0
C2482 a_4905_12113# a_4713_12141# 0
C2483 a_6329_12927# VGND 0.19423f
C2484 a_14946_4905# a_16167_5459# 0.01594f
C2485 a_9875_13765# a_4915_10549# 0.00401f
C2486 a_11108_1773# sky130_fd_sc_hd__mux4_1_0.A2 0.00117f
C2487 VGND a_14108_5463# 0
C2488 a_2289_5307# VDPWR 0.34431f
C2489 a_9811_11277# VGND 1.26863f
C2490 w_11078_4508# a_13046_4563# 0
C2491 a_9557_14759# VDPWR 0.02511f
C2492 a_9715_16323# a_8113_13753# 0
C2493 a_13018_5437# a_13147_5829# 0.00792f
C2494 a_13385_4845# sky130_fd_sc_hd__mux4_1_0.A3 0
C2495 a_2217_5025# a_4045_5047# 0
C2496 a_2217_5025# a_5099_5047# 0.00185f
C2497 VGND a_15281_5825# 0.20007f
C2498 VDPWR w_5712_14949# 0.0786f
C2499 a_9717_13091# a_9811_11277# 0
C2500 a_2289_5307# a_1950_5025# 0.04737f
C2501 a_9753_4963# VGND 0.19554f
C2502 w_4430_16303# a_4625_15373# 0
C2503 a_11289_1773# a_11553_1773# 0
C2504 a_2187_1765# a_3790_1761# 0.00242f
C2505 a_11291_12911# a_10937_12911# 0.09582f
C2506 a_14946_4905# a_15309_4585# 0.01182f
C2507 a_2217_5025# a_4576_5047# 0
C2508 a_3229_5051# w_3668_4962# 0.25055f
C2509 VGND a_11108_1773# 0.08645f
C2510 VGND a_6726_5043# 0
C2511 a_7424_1779# a_7605_2145# 0
C2512 a_4546_2153# w_3638_1702# 0.00139f
C2513 VDPWR w_18554_16401# 0.0754f
C2514 a_13385_4845# w_14764_4500# 0
C2515 a_6915_5043# a_7731_5039# 0
C2516 a_4837_16089# a_6805_15235# 0
C2517 a_13385_4845# a_13046_4563# 0.04737f
C2518 VDPWR a_22274_16171# 0.26198f
C2519 a_8232_1779# a_7869_1779# 0.00985f
C2520 a_11230_4567# w_11050_5382# 0.00104f
C2521 a_6329_12927# a_5851_13769# 0
C2522 a_11291_12911# a_12075_13379# 0
C2523 a_2289_5307# a_3768_5047# 0
C2524 w_11078_4508# a_10611_5471# 0
C2525 a_4183_1787# a_3199_1791# 0.08312f
C2526 w_14764_4500# a_15672_4585# 0.01154f
C2527 a_13439_4955# a_14946_4905# 0
C2528 a_15672_4951# a_15309_4951# 0.00847f
C2529 a_9727_11527# w_9404_11491# 0.01327f
C2530 a_7845_5295# a_8262_5039# 0.03016f
C2531 VDPWR a_16167_5459# 0.13683f
C2532 a_5099_5047# w_6074_6018# 0
C2533 a_10088_5471# sky130_fd_sc_hd__mux4_1_0.A3 0
C2534 a_9515_2143# a_9290_1751# 0.00559f
C2535 a_5606_1757# w_3638_1702# 0
C2536 a_9717_12841# a_4915_10549# 0
C2537 VDPWR a_24774_14701# 0.0823f
C2538 a_9865_15329# w_10674_14933# 0.00546f
C2539 w_10748_13967# a_10937_12911# 0
C2540 a_16871_4938# a_16167_5459# 0.08041f
C2541 a_9727_11527# a_9589_12125# 0
C2542 uo_out[3] uo_out[2] 0.03102f
C2543 a_4635_13809# w_4538_13995# 0.05631f
C2544 a_4711_15373# a_4625_15373# 0.00658f
C2545 a_14846_1739# a_14255_1769# 0.11887f
C2546 a_9811_11277# a_10857_14747# 0.00121f
C2547 a_10046_1777# a_10569_1777# 0
C2548 VGND a_11824_13629# 0.13594f
C2549 a_14864_4585# sky130_fd_sc_hd__mux4_1_0.A3 0
C2550 VDPWR a_8262_5039# 0.2064f
C2551 uio_oe[6] uio_oe[7] 0.03102f
C2552 sky130_fd_sc_hd__mux4_1_0.A1 sky130_fd_sc_hd__mux4_1_0.A0 0.34711f
C2553 a_9587_15357# a_9725_14759# 0
C2554 a_9877_10533# w_9502_10747# 0.0204f
C2555 VDPWR a_15309_4585# 0.17334f
C2556 w_19322_16391# a_19510_16177# 0.02727f
C2557 VDPWR a_4839_12857# 0.75065f
C2558 a_11986_4593# a_12509_4593# 0
C2559 a_11150_5467# w_9180_5386# 0.00188f
C2560 a_3919_1787# VDPWR 0.00117f
C2561 VGND a_11873_15219# 0.00384f
C2562 VDPWR ua[0] 0.07056f
C2563 a_9489_4963# VDPWR 0
C2564 w_10748_13967# a_12075_13379# 0
C2565 sky130_fd_sc_hd__mux4_1_0.A1 a_20384_16179# 0
C2566 a_4837_16089# a_4753_16089# 0.00234f
C2567 w_5906_12121# a_4915_10549# 0
C2568 a_6862_13645# a_4839_12857# 0.00327f
C2569 a_24962_14701# a_24234_14385# 0.1456f
C2570 a_11289_2139# a_11108_1773# 0
C2571 a_14794_1765# a_14255_1769# 0.0725f
C2572 a_14864_4585# w_14764_4500# 0.01793f
C2573 a_13439_4955# VDPWR 0.00924f
C2574 a_13369_1769# a_13201_1769# 0
C2575 a_11091_12911# a_9867_12097# 0
C2576 a_6281_11907# VDPWR 0.2162f
C2577 a_4910_5047# VGND 0
C2578 a_2706_5417# a_2217_5025# 0.0357f
C2579 uio_out[5] uio_out[6] 0.03102f
C2580 a_9585_4597# a_9753_4597# 0
C2581 a_11049_14719# a_9799_16073# 0.29394f
C2582 VDPWR ua[7] 0
C2583 a_4755_13107# a_4839_12857# 0.08134f
C2584 a_13732_1769# a_13315_2025# 0.03016f
C2585 a_6281_11907# a_6862_13645# 0.00248f
C2586 a_9597_13793# a_9587_15357# 0
C2587 a_10088_5471# a_10611_5471# 0
C2588 a_1920_1765# a_2145_2157# 0.00559f
C2589 a_11916_1773# a_10569_1777# 0.08907f
C2590 a_15141_4951# a_15255_4841# 0
C2591 a_4763_14525# a_4903_15345# 0
C2592 a_12966_5463# VGND 0.10729f
C2593 a_13732_1769# w_12824_1684# 0.01154f
C2594 a_7869_1779# sky130_fd_sc_hd__mux4_1_0.A2 0
C2595 a_9809_14509# a_11679_15219# 0.00159f
C2596 a_4627_12141# a_4635_13809# 0
C2597 VDPWR a_11049_14719# 0.36334f
C2598 a_4765_11543# VDPWR 0.31817f
C2599 a_2217_5025# sky130_fd_sc_hd__mux4_1_0.A3 0.11807f
C2600 a_6392_5043# a_6029_5043# 0.00985f
C2601 a_6915_5043# a_8262_5039# 0.08907f
C2602 a_13411_5829# sky130_fd_sc_hd__mux4_1_0.A3 0.00117f
C2603 a_13439_4589# a_13046_4563# 0.02283f
C2604 a_6635_15235# w_5712_14949# 0
C2605 a_4627_12141# a_4905_12113# 0.1206f
C2606 a_7899_5039# w_7354_4954# 0.01092f
C2607 a_8755_1779# VDPWR 1.04258f
C2608 a_4763_14525# VGND 0.00834f
C2609 a_12509_4593# a_11569_4849# 0.13738f
C2610 a_4910_5413# VDPWR 0
C2611 VDPWR sky130_fd_sc_hd__mux4_1_0.A0 2.02287f
C2612 w_11078_4508# sky130_fd_sc_hd__mux4_1_0.A2 0
C2613 a_9290_1751# a_9683_2143# 0.02301f
C2614 ui_in[0] a_24962_14701# 0.02517f
C2615 VDPWR a_7476_1753# 0.29442f
C2616 a_7751_14003# a_4915_10549# 0
C2617 VDPWR a_20384_16179# 0.25715f
C2618 a_9801_12841# w_10674_14933# 0.08813f
C2619 a_3820_5021# a_4045_5047# 0.00487f
C2620 a_9725_5837# VGND 0.25449f
C2621 a_7869_1779# VGND 0.01554f
C2622 a_15255_4841# a_16006_4585# 0.00682f
C2623 a_12481_5467# a_13802_4589# 0
C2624 a_6362_1783# sky130_fd_sc_hd__mux4_1_0.A2 0
C2625 a_10813_13753# a_9799_16073# 0.08387f
C2626 a_3949_5413# a_2217_5025# 0
C2627 a_9727_11277# a_9477_11527# 0.00723f
C2628 a_14325_4589# a_15309_4951# 0.04534f
C2629 a_5636_5017# a_5861_5409# 0.00559f
C2630 a_10895_13753# a_9799_16073# 0
C2631 a_12631_13987# a_11824_13629# 0
C2632 a_5975_5299# a_5861_5409# 0
C2633 a_10813_13753# VDPWR 0.3558f
C2634 w_11078_4508# VGND 0.2898f
C2635 w_9394_13055# a_9867_12097# 0
C2636 a_13385_4845# sky130_fd_sc_hd__mux4_1_0.A2 0
C2637 VDPWR a_10895_13753# 0
C2638 VGND a_11679_15219# 0.00151f
C2639 a_4129_2043# a_4183_2153# 0.03622f
C2640 a_9809_14509# a_9467_13091# 0
C2641 VDPWR a_6029_5409# 0.00962f
C2642 sky130_fd_sc_hd__mux4_1_0.A3 w_6074_6018# 0.05211f
C2643 VDPWR w_14694_1680# 0.50762f
C2644 a_6329_12927# a_4913_13781# 0.0204f
C2645 VDPWR a_6362_2149# 0.01976f
C2646 w_10748_13967# a_9877_10533# 0
C2647 a_19510_16177# w_21318_16395# 0
C2648 a_8566_2145# sky130_fd_sc_hd__mux4_1_0.A2 0
C2649 a_6281_11907# a_6089_11935# 0
C2650 VGND w_9490_15543# 0.11947f
C2651 a_17339_4938# sky130_fd_sc_hd__mux4_1_0.A3 0.0023f
C2652 sky130_fd_sc_hd__mux4_1_0.A2 a_15672_4585# 0
C2653 a_7113_13395# w_9500_13979# 0
C2654 a_6362_1783# VGND 0.01331f
C2655 a_4837_16089# w_4440_14739# 0
C2656 a_5636_5017# a_5765_5409# 0.00792f
C2657 a_14297_5463# a_14888_5433# 0.11887f
C2658 a_4045_5413# a_4159_5303# 0
C2659 a_24318_14385# a_24407_14651# 0
C2660 a_4159_5303# a_5584_5043# 0
C2661 a_13385_4845# VGND 1.17207f
C2662 a_4595_14775# a_4847_14525# 0
C2663 a_5765_5043# VGND 0
C2664 a_1898_5051# a_2217_5025# 0.0073f
C2665 a_11916_2139# VDPWR 0.01968f
C2666 a_9477_11527# a_9867_12097# 0
C2667 a_8566_2145# VGND 0.00244f
C2668 a_7635_5405# a_7899_5405# 0
C2669 a_24241_14651# sky130_fd_sc_hd__mux4_1_0.A3 0.03341f
C2670 a_14946_4905# w_16764_4814# 0.00424f
C2671 VGND a_15672_4585# 0
C2672 a_14136_4589# a_13385_4845# 0.00682f
C2673 a_9467_13091# VGND 0.29689f
C2674 w_5484_4958# a_6029_5409# 0
C2675 a_15239_2131# VDPWR 0.00775f
C2676 ua[6] w_7324_1694# 0
C2677 a_6362_1783# a_5999_1783# 0.00985f
C2678 a_2259_2047# a_2187_1765# 0.25757f
C2679 a_9717_13091# a_9467_13091# 0.02504f
C2680 a_4880_1787# VDPWR 0
C2681 VDPWR w_3638_1702# 0.51485f
C2682 a_3199_1791# a_2187_1765# 0.0046f
C2683 a_14975_1765# sky130_fd_sc_hd__mux4_1_0.A2 0
C2684 w_10748_13967# a_9597_13793# 0
C2685 a_9559_11527# a_9811_11277# 0
C2686 a_10771_14747# a_9799_16073# 0.03093f
C2687 a_14864_4585# sky130_fd_sc_hd__mux4_1_0.A2 0
C2688 a_11958_5467# sky130_fd_sc_hd__mux4_1_0.A3 0
C2689 a_5945_2039# w_7324_1694# 0
C2690 VDPWR a_10771_14747# 0.1486f
C2691 a_4915_10549# a_4839_12857# 0.00243f
C2692 sky130_fd_sc_hd__mux4_1_0.A1 w_9392_16287# 0
C2693 a_9475_14759# w_10674_14933# 0
C2694 a_12135_15219# a_8113_13753# 0.002f
C2695 a_17053_4938# a_16195_4585# 0.00136f
C2696 a_17053_4938# a_17125_4938# 0
C2697 VDPWR a_6127_13769# 0.0014f
C2698 a_10088_5471# VGND 0.10448f
C2699 w_4430_16303# a_6629_15387# 0
C2700 a_4627_12141# a_4713_12141# 0.00658f
C2701 w_11078_4508# a_8785_5039# 0.00114f
C2702 w_22086_16385# a_22274_16171# 0.02727f
C2703 a_5069_1787# a_2187_1765# 0.0019f
C2704 a_9811_11277# a_12135_15219# 0
C2705 a_14975_1765# VGND 0
C2706 ui_in[0] sky130_fd_sc_hd__mux4_1_0.A1 0.00242f
C2707 a_13385_4845# w_12894_4504# 0.10454f
C2708 sky130_fd_sc_hd__mux4_1_0.A3 w_7354_4954# 0.00328f
C2709 a_14864_4585# VGND 0
C2710 VDPWR a_3790_1761# 0.29465f
C2711 a_4597_11543# VDPWR 0.02511f
C2712 VDPWR a_24234_14385# 0.22976f
C2713 VDPWR w_16764_4814# 0.1138f
C2714 a_13439_4589# sky130_fd_sc_hd__mux4_1_0.A2 0
C2715 a_9801_12841# a_11019_12911# 0.00149f
C2716 a_7919_14003# a_7669_14003# 0.00876f
C2717 a_6281_11907# a_4915_10549# 0.43285f
C2718 a_11150_5467# sky130_fd_sc_hd__mux4_1_0.A3 0.00306f
C2719 a_6726_5409# sky130_fd_sc_hd__mux4_1_0.A3 0
C2720 a_11291_12911# w_11718_13593# 0.04962f
C2721 a_9673_15357# a_9587_15357# 0.00658f
C2722 a_3199_1791# a_4546_2153# 0.03325f
C2723 a_4587_13107# a_4839_12857# 0
C2724 a_16871_4938# w_16764_4814# 0.07806f
C2725 a_13385_4845# a_8785_5039# 0
C2726 a_3229_5051# a_4159_5303# 0.21188f
C2727 w_9208_4512# a_9699_4853# 0.10454f
C2728 a_7869_2145# a_8232_2145# 0.00847f
C2729 a_4015_2153# VGND 0.00231f
C2730 w_9392_16287# a_9799_16073# 0.02445f
C2731 a_2313_1791# VGND 0.01474f
C2732 a_9811_11277# w_10872_13125# 0.05304f
C2733 a_13439_4589# VGND 0.01261f
C2734 a_24962_14701# ui_in[1] 0.12867f
C2735 a_3229_5051# a_3949_5047# 0
C2736 a_10046_1777# VDPWR 0.20638f
C2737 VDPWR w_9392_16287# 0.16528f
C2738 a_11958_5467# a_10611_5471# 0.08907f
C2739 a_3820_5021# a_3949_5413# 0.00792f
C2740 a_12320_4959# VDPWR 0
C2741 VGND a_10983_13753# 0.00475f
C2742 w_19322_16391# VGND 0.01227f
C2743 a_13385_4845# a_14916_4559# 0.00446f
C2744 w_4440_14739# a_4849_11293# 0.00324f
C2745 a_5809_14763# a_6629_15387# 0
C2746 ui_in[0] VDPWR 0.40754f
C2747 w_1768_1706# a_3738_1787# 0.00188f
C2748 a_14325_4589# a_15309_4585# 0.08312f
C2749 a_15281_5459# a_15017_5459# 0
C2750 a_2217_5025# VGND 1.11075f
C2751 a_4837_16089# a_4625_15373# 0
C2752 a_10116_4597# sky130_fd_sc_hd__mux4_1_0.A2 0
C2753 VDPWR w_4540_10763# 0.166f
C2754 VGND a_13411_5829# 0.20231f
C2755 a_14864_4585# w_12894_4504# 0.00188f
C2756 a_5999_2149# a_2187_1765# 0
C2757 a_12966_5463# a_11541_5723# 0
C2758 VDPWR a_13147_5829# 0
C2759 a_4627_12141# w_4538_13995# 0
C2760 a_9515_2143# a_9683_2143# 0
C2761 a_11178_4593# a_10639_4597# 0.0725f
C2762 a_5069_1787# a_5606_1757# 0.11545f
C2763 VDPWR ua[5] 0.00178f
C2764 w_6756_13609# a_7173_15235# 0
C2765 a_9360_4571# w_7354_4954# 0
C2766 uo_out[3] uo_out[4] 0.03102f
C2767 a_11873_15219# a_12135_15219# 0
C2768 VDPWR w_9404_11491# 0.16044f
C2769 a_14108_5829# a_14297_5463# 0
C2770 a_23511_14335# sky130_fd_sc_hd__mux4_1_0.A3 0.00544f
C2771 a_11150_5467# a_10611_5471# 0.0725f
C2772 a_11427_5833# a_11202_5441# 0.00559f
C2773 w_9180_5386# a_9725_5471# 0.01092f
C2774 a_11569_4849# sky130_fd_sc_hd__mux4_1_0.A3 0
C2775 a_8262_5405# a_7899_5405# 0.00847f
C2776 VGND a_2049_2157# 0.00311f
C2777 a_4515_11543# a_4839_12857# 0
C2778 a_13105_1769# a_12976_1743# 0.00758f
C2779 a_9489_4963# a_9308_4597# 0
C2780 VGND a_10116_4597# 0.01145f
C2781 w_22086_16385# sky130_fd_sc_hd__mux4_1_0.A0 0.00709f
C2782 a_11916_1773# VDPWR 0.20655f
C2783 a_3919_2153# a_2187_1765# 0
C2784 a_12292_5467# VDPWR 0
C2785 VDPWR a_9589_12125# 0.38028f
C2786 VDPWR a_9238_1777# 0.07483f
C2787 w_4528_15559# a_4513_14775# 0
C2788 VDPWR a_6087_14735# 0.36336f
C2789 a_12509_4593# a_13802_4955# 0.03325f
C2790 a_16195_4585# a_16006_4951# 0
C2791 a_5069_1787# w_6044_2758# 0
C2792 a_15239_2131# a_14975_2131# 0
C2793 a_13439_4589# w_12894_4504# 0.01092f
C2794 VDPWR a_11051_11919# 0
C2795 a_11986_4593# a_10611_5471# 0
C2796 a_9753_4963# a_9585_4963# 0
C2797 a_9465_16323# a_9587_15357# 0.00144f
C2798 a_2343_5051# a_2289_5307# 0.00386f
C2799 w_22086_16385# a_20384_16179# 0
C2800 VGND w_6074_6018# 0.0297f
C2801 a_21506_16181# w_22960_16387# 0
C2802 a_12509_4593# a_13411_5463# 0
C2803 VDPWR a_11202_5441# 0.30708f
C2804 a_6862_13645# a_6087_14735# 0
C2805 w_11078_4508# a_11541_5723# 0
C2806 a_11091_12911# VGND 0.00291f
C2807 a_3010_1791# a_2187_1765# 0
C2808 a_7701_1779# a_7815_2035# 0
C2809 a_11569_4849# a_13046_4563# 0.00492f
C2810 a_7454_5039# VDPWR 0.07407f
C2811 a_8113_13753# w_9402_14723# 0.00353f
C2812 VGND a_17339_4938# 0
C2813 a_24241_14651# sky130_fd_sc_hd__mux4_1_0.A2 0.03575f
C2814 a_4903_15345# w_6570_15449# 0
C2815 VDPWR a_13315_2025# 0.34547f
C2816 VDPWR w_12824_1684# 0.51496f
C2817 a_8113_13753# a_7173_15235# 0.00434f
C2818 a_15978_5459# a_16167_5459# 0
C2819 a_14864_4585# a_14916_4559# 0.1439f
C2820 sky130_fd_sc_hd__mux4_1_0.A2 a_14255_1769# 0.00715f
C2821 a_9809_14509# w_9394_13055# 0
C2822 VGND w_6570_15449# 0.00665f
C2823 a_7113_13395# a_5975_12927# 0
C2824 a_9811_11277# w_9402_14723# 0.00324f
C2825 a_23511_14335# a_23677_14335# 0.00648f
C2826 a_4765_11543# a_4515_11543# 0.02504f
C2827 VDPWR a_13774_5463# 0.20622f
C2828 a_15644_5825# a_14297_5463# 0.03325f
C2829 a_5606_1757# a_5999_2149# 0.02301f
C2830 a_13774_5829# VDPWR 0.01982f
C2831 a_13018_5437# w_12866_5378# 0.05213f
C2832 a_12976_1743# VDPWR 0.29521f
C2833 a_15227_5715# a_14888_5433# 0.04737f
C2834 sky130_fd_sc_hd__mux4_1_0.A3 sky130_fd_sc_hd__mux4_1_0.VPB 0.08221f
C2835 a_7731_5039# a_7506_5013# 0.00487f
C2836 VGND a_14255_1769# 0.67529f
C2837 a_10639_4597# a_11595_5467# 0
C2838 sky130_fd_sc_hd__mux4_1_0.A1 ui_in[1] 0.00113f
C2839 a_11569_4849# a_10611_5471# 0
C2840 VGND w_21318_16395# 0.01283f
C2841 a_15045_4585# a_15309_4585# 0
C2842 a_5554_1783# a_4129_2043# 0
C2843 a_7454_5039# w_5484_4958# 0.00188f
C2844 VDPWR a_14066_1769# 0
C2845 a_12881_13987# sky130_fd_sc_hd__mux4_1_0.A1 0
C2846 a_9875_13765# a_9811_11277# 0.26616f
C2847 a_4503_16339# w_4528_15559# 0.0035f
C2848 sky130_fd_sc_hd__mux4_1_0.A3 a_14888_5433# 0.00509f
C2849 a_5636_5017# a_5099_5047# 0.11566f
C2850 a_12135_15219# a_11679_15219# 0
C2851 a_11958_5467# VGND 0.01767f
C2852 a_15113_5825# a_15227_5715# 0
C2853 w_9394_13055# VGND 0.07276f
C2854 VDPWR a_4505_13107# 0.38927f
C2855 VDPWR w_9500_13979# 0.17935f
C2856 a_5975_5299# a_5099_5047# 0.2115f
C2857 a_6915_5043# a_7454_5039# 0.0725f
C2858 a_15255_4841# a_16195_4585# 0.14436f
C2859 a_15255_4841# a_17125_4938# 0
C2860 a_14946_4905# a_17125_5265# 0
C2861 a_8232_1779# w_7324_1694# 0.01154f
C2862 a_24318_14385# sky130_fd_sc_hd__mux4_1_0.A3 0.04268f
C2863 a_5554_1783# a_5735_2149# 0
C2864 a_13732_2135# a_13315_2025# 0.06611f
C2865 w_9394_13055# a_9717_13091# 0.01327f
C2866 a_11916_1773# a_12439_1773# 0
C2867 a_13732_2135# w_12824_1684# 0.00139f
C2868 a_5945_2039# w_5454_1698# 0.10454f
C2869 VGND a_6805_15235# 0.00334f
C2870 VDPWR w_4442_11507# 0.16044f
C2871 a_15113_5825# sky130_fd_sc_hd__mux4_1_0.A3 0
C2872 w_14764_4500# a_14888_5433# 0
C2873 VDPWR a_6021_13769# 0
C2874 VGND w_7354_4954# 0.29951f
C2875 a_17339_4938# a_8785_5039# 0.00688f
C2876 a_11986_4593# sky130_fd_sc_hd__mux4_1_0.A2 0
C2877 a_8566_1779# a_7815_2035# 0.00682f
C2878 w_10868_12105# a_9811_11277# 0.0984f
C2879 w_14736_5374# a_15644_5459# 0.01154f
C2880 a_12439_1773# a_13315_2025# 0.21148f
C2881 a_10450_4963# a_10639_4597# 0
C2882 VDPWR w_3668_4962# 0.51463f
C2883 a_12439_1773# w_12824_1684# 0.24987f
C2884 a_11150_5467# VGND 0.08811f
C2885 a_3820_5021# VGND 0.40141f
C2886 a_6726_5409# VGND 0.00245f
C2887 a_7113_13395# a_7847_14003# 0.00121f
C2888 a_4755_13107# a_4505_13107# 0.02504f
C2889 a_9477_11527# VGND 0.29765f
C2890 VDPWR a_4721_13809# 0.003f
C2891 a_2259_2047# VDPWR 0.3445f
C2892 VDPWR ui_in[1] 0.10597f
C2893 a_3199_1791# VDPWR 1.05386f
C2894 a_12881_13987# VDPWR 0
C2895 sky130_fd_sc_hd__mux4_1_0.A2 a_12320_4593# 0
C2896 a_4849_11293# a_4765_11293# 0.00206f
C2897 a_6635_15235# a_6087_14735# 0.08954f
C2898 sky130_fd_sc_hd__mux4_1_0.A2 a_12924_1769# 0.00116f
C2899 a_9717_12841# a_9811_11277# 0
C2900 a_14946_4905# a_15644_5459# 0.00474f
C2901 w_4540_10763# a_4915_10549# 0.0204f
C2902 a_9419_2143# sky130_fd_sc_hd__mux4_1_0.A2 0
C2903 a_9865_15329# a_9799_16073# 0.50561f
C2904 a_11986_4593# VGND 0.01315f
C2905 a_17125_5265# VDPWR 0
C2906 a_12976_1743# a_12439_1773# 0.11543f
C2907 a_9875_13765# a_11824_13629# 0
C2908 a_9865_15329# VDPWR 0.24549f
C2909 a_11351_13753# a_9799_16073# 0.00515f
C2910 a_12481_5467# a_12966_5463# 0.0754f
C2911 a_4915_10549# w_9404_11491# 0.00173f
C2912 VGND a_4753_16089# 0.00773f
C2913 a_15602_1765# sky130_fd_sc_hd__mux4_1_0.A2 0
C2914 a_5069_1787# VDPWR 1.04264f
C2915 w_3668_4962# a_3768_5047# 0.01793f
C2916 a_11351_13753# VDPWR 0.38708f
C2917 a_15141_4951# a_16195_4585# 0
C2918 a_6329_12927# w_5906_12121# 0
C2919 a_4755_12857# a_4849_11293# 0
C2920 a_11569_4849# sky130_fd_sc_hd__mux4_1_0.A2 0
C2921 a_11291_12911# a_11243_11891# 0.00298f
C2922 VGND a_12320_4593# 0
C2923 VGND a_12924_1769# 0.08648f
C2924 a_10569_1777# a_11553_2139# 0.04534f
C2925 a_9467_13091# w_10872_13125# 0
C2926 a_9419_2143# VGND 0.00305f
C2927 a_9589_12125# a_4915_10549# 0.00128f
C2928 a_12250_1773# sky130_fd_sc_hd__mux4_1_0.A2 0
C2929 a_9809_14509# a_9587_15357# 0.00215f
C2930 a_15255_4841# a_14297_5463# 0
C2931 a_1868_1791# a_2187_1765# 0.0073f
C2932 sky130_fd_sc_hd__mux4_1_0.A2 w_7324_1694# 0.00331f
C2933 VDPWR a_7424_1779# 0.07407f
C2934 ui_in[2] ui_in[1] 0.03102f
C2935 a_4597_11543# a_4515_11543# 0.00641f
C2936 VGND a_7919_14003# 0
C2937 a_15602_1765# VGND 0.01439f
C2938 a_23511_14335# VGND 0.23646f
C2939 w_7354_4954# a_8785_5039# 0.0206f
C2940 sky130_fd_sc_hd__mux4_1_0.A3 a_9725_5471# 0
C2941 a_4183_2153# w_3638_1702# 0
C2942 a_5069_1787# a_5735_1783# 0
C2943 w_12566_13951# sky130_fd_sc_hd__mux4_1_0.A1 0.02092f
C2944 a_2289_5307# a_2343_5417# 0.03622f
C2945 a_9290_1751# a_9629_2033# 0.04737f
C2946 a_11569_4849# VGND 1.20507f
C2947 VDPWR a_15644_5459# 0.2042f
C2948 a_15602_2131# VDPWR 0.01894f
C2949 a_13201_2135# sky130_fd_sc_hd__mux4_1_0.A2 0
C2950 VGND a_12250_1773# 0
C2951 a_9683_1777# a_9629_2033# 0.00386f
C2952 VGND w_7324_1694# 0.29306f
C2953 VDPWR a_6696_2149# 0
C2954 a_5975_5299# sky130_fd_sc_hd__mux4_1_0.A3 0.00228f
C2955 a_11230_4567# sky130_fd_sc_hd__mux4_1_0.A3 0
C2956 a_11359_4959# a_11230_4567# 0.00792f
C2957 w_10748_13967# a_11243_11891# 0
C2958 a_17053_4938# sky130_fd_sc_hd__mux4_1_0.A3 0
C2959 a_4837_16089# a_6629_15387# 0.27498f
C2960 VGND a_9587_15357# 0.24327f
C2961 a_2259_2047# a_2676_1791# 0.03016f
C2962 VDPWR a_4847_14525# 0.36398f
C2963 a_3199_1791# a_2676_1791# 0
C2964 a_13357_5719# a_13774_5463# 0.03016f
C2965 a_11499_2029# a_11916_2139# 0.06611f
C2966 a_9599_10561# w_9404_11491# 0
C2967 a_14108_5829# sky130_fd_sc_hd__mux4_1_0.A3 0
C2968 sky130_fd_sc_hd__mux4_1_0.A3 a_13802_4955# 0
C2969 a_4183_2153# a_3790_1761# 0.02301f
C2970 a_9801_12841# a_9799_16073# 0.4639f
C2971 sky130_fd_sc_hd__mux4_1_0.A2 sky130_fd_sc_hd__mux4_1_0.VPB 0.08268f
C2972 VGND w_9502_10747# 0.12086f
C2973 a_12481_5467# a_13385_4845# 0
C2974 a_13774_5829# a_13357_5719# 0.06611f
C2975 a_5999_2149# VDPWR 0.00848f
C2976 VGND a_13201_2135# 0.00231f
C2977 a_2706_5417# w_1798_4966# 0.00139f
C2978 a_9715_16323# a_9587_15357# 0
C2979 a_9801_12841# VDPWR 0.75043f
C2980 sky130_fd_sc_hd__mux4_1_0.A3 a_13411_5463# 0
C2981 a_9599_10561# a_9589_12125# 0
C2982 VDPWR a_2049_1791# 0.00125f
C2983 a_4635_13809# VDPWR 0.37531f
C2984 a_4515_11543# w_4540_10763# 0.0035f
C2985 VDPWR w_16298_16411# 0.07652f
C2986 a_4903_15345# w_4440_14739# 0.00599f
C2987 w_12566_13951# a_9799_16073# 0
C2988 VDPWR a_9557_5471# 0
C2989 w_9500_13979# a_4915_10549# 0.00206f
C2990 a_7869_1779# a_6885_1783# 0.08312f
C2991 a_4763_14525# a_4513_14775# 0.00723f
C2992 a_4905_12113# VDPWR 0.28921f
C2993 a_2259_2047# a_2313_2157# 0.03622f
C2994 a_4880_2153# VGND 0.00245f
C2995 w_12566_13951# VDPWR 0.07508f
C2996 VGND sky130_fd_sc_hd__mux4_1_0.VPB 0.01738f
C2997 a_24318_14385# sky130_fd_sc_hd__mux4_1_0.A2 0.05111f
C2998 VGND w_4440_14739# 0.07437f
C2999 a_11569_4849# w_12894_4504# 0
C3000 a_8755_1779# a_9419_1777# 0
C3001 a_3919_2153# VDPWR 0
C3002 a_23511_14701# sky130_fd_sc_hd__mux4_1_0.A1 0.04613f
C3003 w_6756_13609# a_4839_12857# 0.00515f
C3004 w_4442_11507# a_4915_10549# 0
C3005 VDPWR a_6911_15235# 0
C3006 a_9515_1777# a_9629_2033# 0
C3007 a_7815_2035# a_7701_2145# 0
C3008 VGND a_14888_5433# 0.40147f
C3009 a_15644_5825# a_15227_5715# 0.06611f
C3010 a_10639_4597# a_11455_4593# 0
C3011 a_7845_5295# a_7899_5405# 0.03622f
C3012 VDPWR w_9492_12311# 0.17848f
C3013 sky130_fd_sc_hd__mux4_1_0.A3 a_8596_5039# 0
C3014 a_11331_5833# VDPWR 0
C3015 a_3010_1791# VDPWR 0
C3016 a_11569_4849# a_8785_5039# 0
C3017 VGND a_2706_5051# 0.01359f
C3018 a_11230_4567# a_10611_5471# 0
C3019 a_4587_13107# a_4505_13107# 0.00641f
C3020 a_6362_1783# a_6885_1783# 0
C3021 a_4849_11293# a_6129_12927# 0
C3022 a_11291_12911# VGND 0.19423f
C3023 a_4183_1787# a_2187_1765# 0
C3024 a_4755_13107# a_4635_13809# 0
C3025 a_10937_12911# a_12075_13379# 0
C3026 a_4213_5047# a_2217_5025# 0
C3027 a_24318_14385# VGND 0.09477f
C3028 a_15644_5825# sky130_fd_sc_hd__mux4_1_0.A3 0.00186f
C3029 a_13175_4955# a_13046_4563# 0.00792f
C3030 a_11958_5467# a_11541_5723# 0.03016f
C3031 a_9753_4597# a_9489_4597# 0
C3032 VDPWR a_5975_12927# 0.1592f
C3033 a_6281_11907# w_6756_13609# 0.00315f
C3034 a_9467_13091# a_9875_13765# 0
C3035 a_15113_5825# VGND 0.00231f
C3036 VDPWR a_7899_5405# 0.00948f
C3037 a_9585_4597# VDPWR 0.00132f
C3038 uio_in[0] ui_in[7] 0.03102f
C3039 a_11916_2139# w_11008_1688# 0.00139f
C3040 a_6862_13645# a_5975_12927# 0
C3041 a_9597_13793# a_9683_13793# 0.00658f
C3042 a_9290_1751# w_9138_1692# 0.05213f
C3043 VDPWR w_5910_13141# 0.0888f
C3044 w_4530_12327# a_4505_13107# 0.0035f
C3045 a_6329_12927# a_4839_12857# 0.08252f
C3046 a_13105_2135# a_12924_1769# 0
C3047 a_11623_4959# sky130_fd_sc_hd__mux4_1_0.A3 0
C3048 a_15141_4585# VDPWR 0
C3049 a_9332_5445# a_9557_5471# 0.00487f
C3050 a_11623_4959# a_11359_4959# 0
C3051 VDPWR a_6029_5043# 0.17684f
C3052 a_2217_5025# a_3040_5417# 0
C3053 a_9683_1777# w_9138_1692# 0.01092f
C3054 a_13201_1769# sky130_fd_sc_hd__mux4_1_0.A2 0
C3055 a_6089_11935# a_4905_12113# 0
C3056 a_9475_14759# a_9799_16073# 0
C3057 a_23511_14701# VDPWR 0.07721f
C3058 a_21506_16181# a_19510_16177# 0
C3059 a_6389_13769# a_6629_15387# 0
C3060 a_1898_5051# w_1798_4966# 0.01793f
C3061 a_14946_4905# w_12866_5378# 0
C3062 a_16006_4951# sky130_fd_sc_hd__mux4_1_0.A3 0
C3063 w_10748_13967# VGND 0.01862f
C3064 a_12481_5467# a_13439_4589# 0
C3065 a_9475_14759# VDPWR 0.3877f
C3066 a_12509_4593# a_13271_4589# 0
C3067 a_9489_4963# a_9753_4963# 0
C3068 a_10088_5837# VDPWR 0.01964f
C3069 a_6281_11907# a_8113_13753# 0.00287f
C3070 a_11916_1773# a_11553_1773# 0.00985f
C3071 w_9392_17212# a_6629_15387# 0.02743f
C3072 a_9699_4853# w_9180_5386# 0.00166f
C3073 a_11202_5441# a_11331_5467# 0.00758f
C3074 a_4837_16089# w_4430_16303# 0.02445f
C3075 a_6635_15235# a_4847_14525# 0.17824f
C3076 a_6281_11907# a_6329_12927# 0.00298f
C3077 ua[4] a_14975_1765# 0
C3078 VDPWR a_15185_2021# 0.33214f
C3079 VGND a_13201_1769# 0
C3080 w_20196_16393# a_21506_16181# 0
C3081 a_4515_11543# a_4505_13107# 0.00102f
C3082 a_12481_5467# a_13411_5829# 0.04534f
C3083 a_14888_5433# a_8785_5039# 0
C3084 a_11049_14719# a_8113_13753# 0.09735f
C3085 a_6915_5043# a_7899_5405# 0.04534f
C3086 a_9467_13091# a_9717_12841# 0.00723f
C3087 a_9559_11527# a_9477_11527# 0.00641f
C3088 a_9671_5727# a_11202_5441# 0.00446f
C3089 a_9332_5445# a_7899_5405# 0
C3090 a_17254_16187# w_17940_16403# 0.05645f
C3091 w_5484_4958# a_6029_5043# 0.01092f
C3092 a_14846_1739# a_15071_2131# 0.00559f
C3093 VDPWR a_4713_12141# 0.00297f
C3094 a_9811_11277# a_11049_14719# 0.00179f
C3095 a_4515_11543# w_4442_11507# 0.06993f
C3096 w_7604_13967# a_9597_13793# 0
C3097 a_11499_2029# a_11916_1773# 0.03016f
C3098 VDPWR a_7847_14003# 0
C3099 a_11230_4567# sky130_fd_sc_hd__mux4_1_0.A2 0
C3100 a_17254_16187# a_18128_16189# 0.10467f
C3101 a_4159_5303# VDPWR 0.34523f
C3102 a_9515_2143# a_9629_2033# 0
C3103 a_4903_15345# a_4625_15373# 0.12165f
C3104 sky130_fd_sc_hd__mux4_1_0.A2 w_5454_1698# 0.00165f
C3105 w_12866_5378# VDPWR 0.51437f
C3106 VGND a_9725_5471# 0.10237f
C3107 a_11623_4959# a_10611_5471# 0
C3108 a_23731_14309# a_24241_14651# 0.02645f
C3109 a_15255_4841# a_15227_5715# 0.00177f
C3110 a_14864_4585# a_15045_4951# 0
C3111 a_9875_13765# a_10983_13753# 0.00104f
C3112 a_15071_1765# a_14255_1769# 0
C3113 a_14916_4559# a_14888_5433# 0
C3114 a_6635_15235# a_6911_15235# 0.00119f
C3115 a_4015_2153# a_4129_2043# 0
C3116 VGND a_4625_15373# 0.24327f
C3117 a_11499_2029# w_12824_1684# 0
C3118 a_4837_16089# w_7604_13967# 0
C3119 a_23677_14701# sky130_fd_sc_hd__mux4_1_0.VPB 0.01733f
C3120 a_9801_12841# a_4915_10549# 0
C3121 VDPWR a_3949_5047# 0.00114f
C3122 a_5636_5017# VGND 0.40145f
C3123 a_11351_13753# a_11906_13629# 0.00183f
C3124 a_11569_4849# a_11541_5723# 0.00177f
C3125 a_10380_2143# a_10569_1777# 0
C3126 a_9877_10533# a_12075_13379# 0.16207f
C3127 a_5975_5299# VGND 1.20008f
C3128 a_15255_4841# sky130_fd_sc_hd__mux4_1_0.A3 0
C3129 a_9465_16323# a_9715_16073# 0.00723f
C3130 a_11230_4567# VGND 0.38979f
C3131 VDPWR a_11553_2139# 0.00968f
C3132 a_11623_4593# a_10611_5471# 0
C3133 a_4723_10577# VDPWR 0.00176f
C3134 a_17053_4938# VGND 0
C3135 a_10813_13753# a_9811_11277# 0.17627f
C3136 a_9811_11277# a_10895_13753# 0
C3137 a_4905_12113# a_4915_10549# 0.0298f
C3138 VGND w_5454_1698# 0.29362f
C3139 a_5809_14763# a_4837_16089# 0.03093f
C3140 a_7845_5295# a_10116_4963# 0
C3141 a_14108_5829# VGND 0.00248f
C3142 a_11499_2029# a_12976_1743# 0.00492f
C3143 VGND a_13802_4955# 0.18285f
C3144 w_5484_4958# a_4159_5303# 0
C3145 a_1868_1791# VDPWR 0.08418f
C3146 VGND a_4765_11293# 0.00834f
C3147 w_10748_13967# a_12631_13987# 0
C3148 ua[5] w_11008_1688# 0
C3149 a_15255_4841# w_14764_4500# 0.10454f
C3150 VGND a_13411_5463# 0.01681f
C3151 a_3820_5021# a_4213_5047# 0.02283f
C3152 w_9492_12311# a_4915_10549# 0.00193f
C3153 VDPWR a_6392_5043# 0.20634f
C3154 a_11049_14719# a_11824_13629# 0
C3155 sky130_fd_sc_hd__mux4_1_0.A2 a_7605_1779# 0
C3156 w_6570_15449# a_7173_15235# 0.01567f
C3157 a_12713_13987# a_11351_13753# 0
C3158 a_4913_13781# w_4440_14739# 0
C3159 VDPWR a_10116_4963# 0.05672f
C3160 a_5554_1783# w_3638_1702# 0.00227f
C3161 a_11178_4593# VDPWR 0.09319f
C3162 a_15978_5825# a_15227_5715# 0.00696f
C3163 VGND w_1798_4966# 0.29762f
C3164 a_4045_5413# VDPWR 0
C3165 a_3199_1791# a_4183_2153# 0.04534f
C3166 a_4763_14775# a_4849_11293# 0
C3167 a_2145_1791# VDPWR 0.00107f
C3168 a_7701_1779# VDPWR 0
C3169 VDPWR w_4538_13995# 0.17926f
C3170 a_9753_4597# VDPWR 0.26479f
C3171 a_11091_12911# a_9875_13765# 0
C3172 VDPWR a_5584_5043# 0.07424f
C3173 a_4755_12857# VGND 0.00847f
C3174 a_11916_1773# w_11008_1688# 0.01154f
C3175 a_11049_14719# a_11873_15219# 0.00651f
C3176 a_5999_1783# w_5454_1698# 0.01092f
C3177 a_13175_4955# VGND 0.00329f
C3178 a_15978_5825# sky130_fd_sc_hd__mux4_1_0.A3 0
C3179 a_4763_14525# a_4839_12857# 0
C3180 w_1768_1706# VGND 0.29741f
C3181 a_12481_5467# a_11958_5467# 0
C3182 a_10771_14747# a_8113_13753# 0
C3183 VGND a_8596_5039# 0
C3184 VGND a_7605_1779# 0
C3185 a_9629_2033# a_9683_2143# 0.03622f
C3186 a_7454_5039# a_7506_5013# 0.1439f
C3187 w_4530_12327# a_4635_13809# 0
C3188 VDPWR a_7605_2145# 0
C3189 a_16195_4585# a_17125_4938# 0.19521f
C3190 a_15141_4951# sky130_fd_sc_hd__mux4_1_0.A3 0
C3191 a_15239_1765# a_14975_1765# 0
C3192 a_9801_12841# a_11906_13629# 0
C3193 w_4530_12327# a_4905_12113# 0.0247f
C3194 a_9290_1751# sky130_fd_sc_hd__mux4_1_0.A2 0.00208f
C3195 a_10813_13753# a_11824_13629# 0
C3196 a_15644_5825# VGND 0.18635f
C3197 a_9811_11277# a_10771_14747# 0.10553f
C3198 w_5484_4958# a_6392_5043# 0.01154f
C3199 w_12894_4504# a_13802_4955# 0.00139f
C3200 a_11230_4567# a_8785_5039# 0
C3201 a_5999_2149# a_5831_2149# 0
C3202 a_17053_4938# a_8785_5039# 0.00526f
C3203 a_9683_1777# sky130_fd_sc_hd__mux4_1_0.A2 0
C3204 uio_in[6] uio_in[7] 0.03102f
C3205 a_9475_14759# a_4915_10549# 0
C3206 w_5484_4958# a_5584_5043# 0.01793f
C3207 a_6805_15235# a_7173_15235# 0
C3208 a_6915_5043# a_6392_5043# 0
C3209 sky130_fd_sc_hd__mux4_1_0.A2 a_11623_4593# 0
C3210 a_11569_4849# a_11595_5833# 0
C3211 a_12976_1743# w_11008_1688# 0
C3212 a_9290_1751# VGND 0.40141f
C3213 w_9208_4512# sky130_fd_sc_hd__mux4_1_0.A3 0
C3214 a_4627_12141# VDPWR 0.38028f
C3215 w_9394_13055# a_9875_13765# 0.00226f
C3216 w_7604_13967# a_6389_13769# 0
C3217 a_11623_4959# VGND 0.19557f
C3218 a_10639_4597# VDPWR 1.11949f
C3219 a_9683_1777# VGND 0.01556f
C3220 a_23731_14309# a_23511_14335# 0.0457f
C3221 a_4905_12113# a_4515_11543# 0
C3222 a_4546_2153# a_2187_1765# 0
C3223 a_16006_4951# VGND 0
C3224 VDPWR a_11595_5467# 0.17063f
C3225 a_14946_4905# a_15113_5459# 0
C3226 VGND a_11623_4593# 0.01251f
C3227 w_9392_16287# a_8113_13753# 0.00656f
C3228 a_9699_4853# sky130_fd_sc_hd__mux4_1_0.A3 0
C3229 a_15672_4585# a_15309_4585# 0.00985f
C3230 w_10674_14933# a_9799_16073# 0.00872f
C3231 a_8566_1779# VDPWR 0
C3232 a_7869_2145# sky130_fd_sc_hd__mux4_1_0.A2 0
C3233 a_3229_5051# VDPWR 1.05177f
C3234 a_7847_14003# a_4915_10549# 0
C3235 a_4183_1787# VDPWR 0.17525f
C3236 VDPWR w_10674_14933# 0.07858f
C3237 a_11049_14719# a_11679_15219# 0.00232f
C3238 a_13439_4955# a_13385_4845# 0.03622f
C3239 a_7869_1779# a_7476_1753# 0.02283f
C3240 VDPWR a_7635_5405# 0
C3241 w_6756_13609# a_6087_14735# 0
C3242 a_1920_1765# VGND 0.40886f
C3243 w_11718_13593# a_12075_13379# 0.03222f
C3244 a_9589_12125# a_9675_12125# 0.00658f
C3245 a_5809_14763# a_4849_11293# 0.10553f
C3246 a_4627_12141# a_4755_13107# 0
C3247 a_11597_15219# a_12075_13379# 0
C3248 a_5606_1757# a_2187_1765# 0.0021f
C3249 a_9515_1777# sky130_fd_sc_hd__mux4_1_0.A2 0
C3250 w_7604_13967# a_7669_14003# 0.05168f
C3251 a_9557_5837# sky130_fd_sc_hd__mux4_1_0.A3 0
C3252 a_7815_2035# VDPWR 0.34502f
C3253 a_14066_2135# sky130_fd_sc_hd__mux4_1_0.A2 0
C3254 a_9597_13793# a_9725_14759# 0
C3255 w_12866_5378# a_13357_5719# 0.10454f
C3256 a_7869_2145# VGND 0.20146f
C3257 a_14325_4589# a_15141_4585# 0
C3258 a_2217_5025# a_2289_5307# 0.25757f
C3259 a_21506_16181# VGND 0.25659f
C3260 a_12809_13987# a_12075_13379# 0.00121f
C3261 a_15255_4841# sky130_fd_sc_hd__mux4_1_0.A2 0
C3262 w_11532_15433# a_11597_15219# 0.08205f
C3263 a_4723_10577# a_4915_10549# 0
C3264 a_18128_16189# w_17940_16403# 0.02697f
C3265 a_17254_16187# w_17066_16401# 0.02727f
C3266 a_3919_2153# a_4183_2153# 0
C3267 VGND a_6129_12927# 0.00291f
C3268 a_12481_5467# a_11569_4849# 0
C3269 a_10450_4963# VDPWR 0
C3270 a_3229_5051# a_3768_5047# 0.0725f
C3271 a_13271_4589# a_13046_4563# 0.00487f
C3272 w_6044_2758# a_2187_1765# 0.02708f
C3273 a_9515_1777# VGND 0
C3274 w_9138_1692# a_9683_2143# 0
C3275 VDPWR a_15113_5459# 0
C3276 w_9208_4512# a_9360_4571# 0.05213f
C3277 a_11291_12911# w_10872_13125# 0.02303f
C3278 a_7919_14003# a_7173_15235# 0
C3279 a_23731_14309# sky130_fd_sc_hd__mux4_1_0.VPB 0.22258f
C3280 a_9811_11277# w_9404_11491# 0.02399f
C3281 a_14066_2135# VGND 0.00244f
C3282 w_11050_5382# sky130_fd_sc_hd__mux4_1_0.A3 0.00615f
C3283 a_9671_5727# a_9557_5471# 0
C3284 a_8755_1779# a_8566_2145# 0
C3285 w_10748_13967# a_12135_15219# 0
C3286 a_24152_14385# sky130_fd_sc_hd__mux4_1_0.A3 0.01336f
C3287 a_17254_16187# a_19510_16177# 0
C3288 a_6329_12927# a_6087_14735# 0
C3289 w_5786_13983# a_6629_15387# 0
C3290 a_14836_5459# w_12866_5378# 0.00188f
C3291 a_15255_4841# VGND 0.00379f
C3292 a_9811_11277# a_9589_12125# 0.0022f
C3293 VGND a_9715_16073# 0.00773f
C3294 a_11108_1773# ua[5] 0
C3295 a_9699_4853# a_10611_5471# 0
C3296 a_6944_13645# a_7113_13395# 0
C3297 a_11051_11919# a_9811_11277# 0
C3298 a_11160_1747# a_9629_2033# 0.00446f
C3299 a_9699_4853# a_9360_4571# 0.04737f
C3300 a_11230_4567# a_11541_5723# 0
C3301 a_9587_15357# w_9402_14723# 0.00155f
C3302 a_10937_12911# a_9867_12097# 0
C3303 VDPWR a_4595_14775# 0.02511f
C3304 a_10639_4597# a_11986_4959# 0.03325f
C3305 a_23731_14309# a_24318_14385# 0.02707f
C3306 a_4903_15345# a_6629_15387# 0
C3307 a_13018_5437# a_12994_4589# 0
C3308 a_4576_5413# w_3668_4962# 0.00139f
C3309 a_15239_1765# a_14255_1769# 0.08312f
C3310 VGND a_6629_15387# 0.40404f
C3311 VDPWR a_10422_5837# 0
C3312 a_10380_2143# VDPWR 0
C3313 a_9877_10533# w_11718_13593# 0.00404f
C3314 a_13018_5437# VDPWR 0.28377f
C3315 VGND a_15978_5825# 0.00228f
C3316 a_6885_1783# w_7324_1694# 0.25055f
C3317 w_11050_5382# a_10611_5471# 0.25055f
C3318 a_8262_5405# a_7845_5295# 0.06611f
C3319 a_9877_10533# a_12809_13987# 0
C3320 a_8113_13753# w_9500_13979# 0.00438f
C3321 a_9515_2143# sky130_fd_sc_hd__mux4_1_0.A2 0
C3322 VDPWR a_11019_12911# 0
C3323 VGND a_2079_5051# 0
C3324 a_6329_12927# a_4505_13107# 0
C3325 a_11359_4593# a_10639_4597# 0
C3326 w_9208_4512# sky130_fd_sc_hd__mux4_1_0.A2 0.00107f
C3327 a_15281_5459# a_15644_5459# 0.00985f
C3328 a_16006_4585# sky130_fd_sc_hd__mux4_1_0.A2 0
C3329 VGND a_2676_2157# 0.18903f
C3330 a_9671_5727# a_10088_5837# 0.06611f
C3331 a_9811_11277# w_9500_13979# 0.00123f
C3332 a_15255_4841# a_8785_5039# 0.00102f
C3333 a_9727_11527# VDPWR 0.31817f
C3334 VDPWR a_8262_5405# 0.01999f
C3335 a_4503_16339# a_4753_16089# 0.00723f
C3336 a_15071_2131# sky130_fd_sc_hd__mux4_1_0.A2 0
C3337 a_6392_5409# VDPWR 0.01964f
C3338 VDPWR a_7701_2145# 0
C3339 a_12966_5463# a_13147_5829# 0
C3340 a_22274_16171# w_21318_16395# 0
C3341 a_9515_2143# VGND 0.00231f
C3342 a_7731_5405# a_7899_5405# 0
C3343 w_19322_16391# sky130_fd_sc_hd__mux4_1_0.A0 0.00534f
C3344 VDPWR a_5933_13769# 0
C3345 a_9699_4853# sky130_fd_sc_hd__mux4_1_0.A2 0
C3346 a_4910_5413# a_2217_5025# 0
C3347 w_9208_4512# VGND 0.28745f
C3348 VGND a_16006_4585# 0
C3349 a_14888_5433# a_15017_5459# 0.00758f
C3350 a_11291_12911# a_9875_13765# 0.0204f
C3351 a_4880_2153# a_4129_2043# 0.00696f
C3352 VGND a_11089_13753# 0.00413f
C3353 w_19322_16391# a_20384_16179# 0
C3354 a_24241_14651# a_24774_14701# 0.0098f
C3355 a_3820_5021# a_2289_5307# 0.00446f
C3356 VDPWR a_2079_5417# 0
C3357 a_13271_4589# sky130_fd_sc_hd__mux4_1_0.A2 0
C3358 a_15071_2131# VGND 0.00231f
C3359 a_15255_4841# a_14916_4559# 0.04737f
C3360 a_5554_1783# a_5069_1787# 0.07531f
C3361 VDPWR a_13732_1769# 0.20646f
C3362 uio_out[5] uio_out[4] 0.03102f
C3363 a_11385_2139# a_11553_2139# 0
C3364 a_11160_1747# w_9138_1692# 0
C3365 a_4763_14775# a_4903_15345# 0.00327f
C3366 a_18742_16187# sky130_fd_sc_hd__mux4_1_0.A1 0
C3367 a_1950_5025# a_2079_5417# 0.00792f
C3368 w_4440_14739# a_4513_14775# 0.06993f
C3369 a_9865_15329# a_8113_13753# 0.00176f
C3370 a_10813_13753# a_10983_13753# 0.00167f
C3371 VDPWR a_2187_1765# 1.34565f
C3372 VGND a_2145_2157# 0.0024f
C3373 a_7113_13395# VDPWR 0.24839f
C3374 a_9699_4853# VGND 1.17357f
C3375 a_9877_10533# a_9867_12097# 0.0298f
C3376 VDPWR a_11455_4593# 0.00101f
C3377 w_4530_12327# a_4627_12141# 0.05631f
C3378 a_6392_5409# w_5484_4958# 0.00139f
C3379 a_11351_13753# a_8113_13753# 0
C3380 a_7113_13395# a_6862_13645# 0.10945f
C3381 a_4763_14775# VGND 0.02642f
C3382 a_7899_5405# a_7506_5013# 0.02301f
C3383 a_9865_15329# a_9811_11277# 0.30844f
C3384 a_2217_5025# a_6029_5409# 0
C3385 a_10569_1777# VDPWR 1.05227f
C3386 a_6915_5043# a_8262_5405# 0.03325f
C3387 a_13271_4589# VGND 0
C3388 a_11291_12911# w_10868_12105# 0
C3389 VGND a_9557_5837# 0.00294f
C3390 a_9683_13793# VGND 0.00661f
C3391 a_9332_5445# a_8262_5405# 0
C3392 a_11351_13753# a_9811_11277# 0.00488f
C3393 a_4903_15345# w_4430_16303# 0
C3394 w_6756_13609# a_4847_14525# 0
C3395 a_15602_1765# a_15239_1765# 0.00985f
C3396 a_4913_13781# a_6129_12927# 0
C3397 a_9683_2143# sky130_fd_sc_hd__mux4_1_0.A2 0
C3398 w_10748_13967# a_9875_13765# 0.00175f
C3399 a_5735_1783# a_2187_1765# 0
C3400 a_10937_12911# a_11243_11891# 0
C3401 VGND w_4430_16303# 0.06271f
C3402 a_13147_5463# a_13411_5463# 0
C3403 a_11499_2029# a_11553_2139# 0.03622f
C3404 a_4837_16089# a_6389_13769# 0.00515f
C3405 w_7354_4954# a_8262_5039# 0.01154f
C3406 VDPWR a_4546_2153# 0.01963f
C3407 a_5861_5043# a_6029_5043# 0
C3408 a_3949_5413# a_4213_5413# 0
C3409 a_4627_12141# a_4515_11543# 0
C3410 a_18128_16189# w_17066_16401# 0
C3411 a_10937_12911# a_10965_11919# 0
C3412 VGND w_11050_5382# 0.31672f
C3413 w_11078_4508# a_11202_5441# 0
C3414 a_3040_5051# VGND 0
C3415 VGND a_9683_2143# 0.20145f
C3416 a_18742_16187# VDPWR 0.25742f
C3417 a_11243_11891# a_12075_13379# 0.19825f
C3418 w_11718_13593# a_11597_15219# 0
C3419 w_9208_4512# a_8785_5039# 0.00202f
C3420 a_24152_14385# VGND 0.22746f
C3421 a_24241_14651# sky130_fd_sc_hd__mux4_1_0.A0 0
C3422 a_4503_16339# w_4440_14739# 0
C3423 a_9597_13793# a_7669_14003# 0
C3424 a_4837_16089# a_4849_11293# 0.03118f
C3425 a_15141_4951# a_14916_4559# 0.00559f
C3426 a_16195_4585# sky130_fd_sc_hd__mux4_1_0.A3 0.01978f
C3427 a_17125_4938# sky130_fd_sc_hd__mux4_1_0.A3 0.1015f
C3428 a_4015_2153# a_3790_1761# 0.00559f
C3429 w_21318_16395# sky130_fd_sc_hd__mux4_1_0.A0 0.00562f
C3430 a_12481_5467# a_13802_4955# 0
C3431 a_19510_16177# a_18128_16189# 0
C3432 VDPWR a_24962_14701# 0.21151f
C3433 a_5606_1757# VDPWR 0.29517f
C3434 a_5809_14763# w_5786_13983# 0
C3435 sky130_fd_sc_hd__mux4_1_0.A2 a_13369_2135# 0
C3436 a_12439_1773# a_13732_1769# 0.08907f
C3437 a_9467_13091# w_9404_11491# 0
C3438 a_4903_15345# a_4711_15373# 0.00101f
C3439 a_12481_5467# a_13411_5463# 0.08099f
C3440 a_9465_16323# a_9725_14759# 0
C3441 a_9699_4853# a_8785_5039# 0
C3442 a_9865_15329# a_11824_13629# 0
C3443 a_20384_16179# w_21318_16395# 0.05549f
C3444 ui_in[2] ui_in[3] 0.03102f
C3445 a_9801_12841# a_8113_13753# 0.00389f
C3446 a_2187_1765# a_2676_1791# 0.08982f
C3447 a_16195_4585# w_14764_4500# 0.02202f
C3448 w_7604_13967# VGND 0.00757f
C3449 VDPWR a_9489_4597# 0.0015f
C3450 VGND a_4711_15373# 0.00661f
C3451 a_11351_13753# a_11824_13629# 0.24537f
C3452 a_9467_13091# a_9589_12125# 0.00144f
C3453 a_13018_5437# a_13357_5719# 0.04737f
C3454 a_5809_14763# a_4903_15345# 0.0039f
C3455 a_9801_12841# a_9811_11277# 0.82158f
C3456 w_20196_16393# a_18128_16189# 0
C3457 a_14846_1739# a_14794_1765# 0.1439f
C3458 a_10569_1777# a_12439_1773# 0
C3459 VDPWR w_6044_2758# 0.06793f
C3460 a_14255_1769# w_14694_1680# 0.25055f
C3461 a_17254_16187# VGND 0.26932f
C3462 VGND a_13369_2135# 0.20063f
C3463 a_13243_5463# a_13411_5463# 0
C3464 a_5606_1757# a_5735_1783# 0.00758f
C3465 a_5809_14763# VGND 0.13243f
C3466 a_8232_2145# sky130_fd_sc_hd__mux4_1_0.A2 0
C3467 a_14946_4905# w_14736_5374# 0.02228f
C3468 a_9461_5837# a_9280_5471# 0
C3469 a_9727_11527# a_4915_10549# 0
C3470 a_11331_5467# a_11595_5467# 0
C3471 w_11008_1688# a_11553_2139# 0
C3472 a_2313_2157# a_2187_1765# 0.05199f
C3473 a_7113_13395# a_6635_15235# 0
C3474 a_6944_13645# VDPWR 0.0014f
C3475 a_9461_5471# VDPWR 0.00116f
C3476 a_4513_14775# a_4625_15373# 0
C3477 a_9461_5837# VDPWR 0
C3478 a_15227_5715# a_14297_5463# 0.21188f
C3479 w_7604_13967# a_5851_13769# 0
C3480 a_6885_1783# w_5454_1698# 0.02026f
C3481 a_24407_14651# sky130_fd_sc_hd__mux4_1_0.A3 0
C3482 w_11050_5382# a_8785_5039# 0.00342f
C3483 a_9811_11277# w_9492_12311# 0.00145f
C3484 a_6944_13645# a_6862_13645# 0.00477f
C3485 a_9683_2143# a_10046_2143# 0.00847f
C3486 a_4129_2043# w_5454_1698# 0
C3487 VGND a_8232_2145# 0.18643f
C3488 a_2289_5307# a_2706_5051# 0.03016f
C3489 uio_oe[3] uio_oe[2] 0.03102f
C3490 a_13369_1769# sky130_fd_sc_hd__mux4_1_0.A2 0
C3491 a_14297_5463# sky130_fd_sc_hd__mux4_1_0.A3 0.00709f
C3492 a_5099_5047# a_4576_5047# 0
C3493 a_6329_12927# a_5975_12927# 0.09582f
C3494 a_9809_14509# w_11532_15433# 0.07233f
C3495 a_9877_10533# a_11243_11891# 0.44698f
C3496 a_10937_12911# VGND 0.14511f
C3497 a_15239_2131# a_14255_1769# 0.04534f
C3498 a_5809_14763# a_5851_13769# 0
C3499 a_7113_13395# a_4915_10549# 0.16058f
C3500 a_6281_11907# a_7919_14003# 0
C3501 a_4576_5413# a_4159_5303# 0.06611f
C3502 a_11160_1747# sky130_fd_sc_hd__mux4_1_0.A2 0.00203f
C3503 a_12509_4593# sky130_fd_sc_hd__mux4_1_0.A3 0
C3504 a_6329_12927# w_5910_13141# 0.02303f
C3505 a_9877_10533# a_10965_11919# 0
C3506 a_9801_12841# a_11824_13629# 0.00327f
C3507 w_14736_5374# VDPWR 0.5114f
C3508 a_9467_13091# w_9500_13979# 0
C3509 a_13411_5829# a_13147_5829# 0
C3510 w_14764_4500# a_14297_5463# 0
C3511 a_9549_13091# VGND 0.00171f
C3512 a_13369_1769# VGND 0.01514f
C3513 a_4849_11293# a_6389_13769# 0.00488f
C3514 VGND a_12075_13379# 0.34868f
C3515 a_9475_14759# a_8113_13753# 0.0055f
C3516 sky130_fd_sc_hd__mux4_1_0.A1 a_9799_16073# 0
C3517 a_9599_10561# a_9727_11527# 0
C3518 sky130_fd_sc_hd__mux4_1_0.VPB a_24774_14701# 0.14223f
C3519 a_5861_5409# VGND 0.00233f
C3520 a_6885_1783# a_7605_1779# 0
C3521 w_9180_5386# sky130_fd_sc_hd__mux4_1_0.A3 0.0065f
C3522 VDPWR sky130_fd_sc_hd__mux4_1_0.A1 0.93097f
C3523 a_24241_14651# a_24234_14385# 0.13413f
C3524 a_23511_14335# sky130_fd_sc_hd__mux4_1_0.A0 0.05256f
C3525 VDPWR a_6696_1783# 0
C3526 a_12509_4593# a_13046_4563# 0.11554f
C3527 a_14946_4905# VDPWR 1.2932f
C3528 a_11160_1747# VGND 0.40116f
C3529 a_9475_14759# a_9811_11277# 0.00146f
C3530 a_13105_1769# VDPWR 0.00117f
C3531 a_9865_15329# w_9490_15543# 0.01828f
C3532 VGND w_11532_15433# 0.00665f
C3533 a_4503_16339# a_4625_15373# 0.00144f
C3534 a_9461_5471# a_9332_5445# 0.00758f
C3535 a_9461_5837# a_9332_5445# 0.00792f
C3536 a_6389_13769# a_7669_14003# 0.00196f
C3537 a_14946_4905# a_16871_4938# 0.00632f
C3538 w_4440_14739# a_4839_12857# 0.00408f
C3539 ua[0] sky130_fd_sc_hd__mux4_1_0.VPB 0.02132f
C3540 a_8755_1779# w_7324_1694# 0.01935f
C3541 a_5765_5409# VGND 0.00306f
C3542 a_24318_14385# a_24774_14701# 0.01242f
C3543 a_6362_1783# a_5069_1787# 0.08907f
C3544 a_9280_5471# a_7845_5295# 0
C3545 a_4213_5413# VGND 0.20073f
C3546 a_12994_4589# VDPWR 0.07505f
C3547 a_7476_1753# w_7324_1694# 0.05213f
C3548 a_13243_5829# sky130_fd_sc_hd__mux4_1_0.A3 0
C3549 a_4763_14525# a_4847_14525# 0.00206f
C3550 a_4753_16339# a_4625_15373# 0
C3551 a_11427_5833# VDPWR 0
C3552 a_8596_5405# sky130_fd_sc_hd__mux4_1_0.A3 0
C3553 VGND w_22960_16387# 0.01911f
C3554 VDPWR a_7845_5295# 0.34676f
C3555 a_15602_1765# w_14694_1680# 0.01154f
C3556 a_16195_4585# sky130_fd_sc_hd__mux4_1_0.A2 0
C3557 a_9809_14509# a_9725_14759# 0.07979f
C3558 a_9280_5471# VDPWR 0.07735f
C3559 a_15017_5825# a_14946_4905# 0
C3560 VDPWR a_9799_16073# 1.07863f
C3561 a_9671_5727# a_10422_5837# 0.00696f
C3562 ui_in[0] a_24241_14651# 0.06328f
C3563 a_13774_5829# a_13411_5829# 0.00847f
C3564 a_7899_5039# sky130_fd_sc_hd__mux4_1_0.A3 0
C3565 uio_out[2] uio_out[1] 0.03102f
C3566 a_13105_2135# a_13369_2135# 0
C3567 a_9629_2033# w_9138_1692# 0.10454f
C3568 a_5099_5047# sky130_fd_sc_hd__mux4_1_0.A3 0
C3569 a_5831_2149# a_2187_1765# 0
C3570 sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_sc_hd__mux4_1_0.A0 0.10334f
C3571 w_9180_5386# a_10611_5471# 0.02026f
C3572 a_16195_4585# VGND 0.08121f
C3573 a_17125_4938# VGND 0.16937f
C3574 a_11541_5723# w_11050_5382# 0.10454f
C3575 VDPWR a_6862_13645# 0.09661f
C3576 a_7635_5405# a_7506_5013# 0.00792f
C3577 a_16871_4938# VDPWR 0.07431f
C3578 a_11289_2139# a_11160_1747# 0.00792f
C3579 VDPWR a_1950_5025# 0.30536f
C3580 a_9360_4571# w_9180_5386# 0.00104f
C3581 w_6570_15449# a_6087_14735# 0.06196f
C3582 a_9877_10533# VGND 0.9946f
C3583 a_12631_13987# a_12075_13379# 0.28206f
C3584 a_11291_12911# a_11049_14719# 0
C3585 a_9809_14509# a_9597_13793# 0
C3586 VGND a_9725_14759# 0.02642f
C3587 a_7869_2145# a_6885_1783# 0.04534f
C3588 a_13105_1769# a_12439_1773# 0
C3589 a_5735_1783# VDPWR 0.00115f
C3590 a_3738_1787# VGND 0.08661f
C3591 a_4755_13107# VDPWR 0.31944f
C3592 a_6915_5043# a_7845_5295# 0.21188f
C3593 a_5809_14763# a_4913_13781# 0
C3594 a_4849_11293# w_4432_13071# 0.00299f
C3595 VDPWR a_3768_5047# 0.07396f
C3596 w_11718_13593# a_11243_11891# 0.00315f
C3597 a_2259_2047# a_2313_1791# 0.00386f
C3598 a_9332_5445# a_7845_5295# 0
C3599 w_5484_4958# VDPWR 0.51493f
C3600 a_15017_5825# VDPWR 0
C3601 VGND w_17940_16403# 0.01236f
C3602 a_6629_15387# a_7173_15235# 0.002f
C3603 a_9280_5471# a_9332_5445# 0.1439f
C3604 a_2217_5025# w_3668_4962# 0.00346f
C3605 a_2289_5307# w_1798_4966# 0.10454f
C3606 a_13315_2025# a_14255_1769# 0.13962f
C3607 a_4183_2153# a_2187_1765# 0
C3608 w_9394_13055# a_9589_12125# 0
C3609 a_6915_5043# VDPWR 1.05198f
C3610 a_14255_1769# w_12824_1684# 0.02026f
C3611 a_13732_2135# VDPWR 0.01969f
C3612 VGND a_18128_16189# 0.25249f
C3613 w_20196_16393# a_19510_16177# 0.05645f
C3614 a_9753_4963# a_10116_4963# 0.00847f
C3615 a_10813_13753# a_11291_12911# 0
C3616 a_12809_13987# a_11243_11891# 0.00264f
C3617 a_9332_5445# VDPWR 0.29533f
C3618 a_4837_16089# w_5786_13983# 0.06973f
C3619 a_3229_5051# a_4576_5413# 0.03325f
C3620 a_9467_13091# a_9801_12841# 0.16952f
C3621 a_6089_11935# VDPWR 0
C3622 w_10748_13967# a_11049_14719# 0
C3623 a_9597_13793# VGND 0.24546f
C3624 a_15672_4951# a_14946_4905# 0.18442f
C3625 a_7899_5039# a_9360_4571# 0
C3626 a_6805_15235# a_6087_14735# 0.00366f
C3627 a_9865_15329# a_10983_13753# 0.00818f
C3628 a_4837_16089# a_6003_11935# 0
C3629 a_12509_4593# sky130_fd_sc_hd__mux4_1_0.A2 0
C3630 a_9717_13091# a_9597_13793# 0
C3631 a_5606_1757# a_5831_2149# 0.00559f
C3632 a_9477_11527# w_9404_11491# 0.06993f
C3633 a_15281_5459# a_15113_5459# 0
C3634 VDPWR a_12439_1773# 1.04462f
C3635 a_4837_16089# a_4903_15345# 0.50561f
C3636 a_11351_13753# a_10983_13753# 0
C3637 VDPWR a_2676_1791# 0.20903f
C3638 a_13271_4955# sky130_fd_sc_hd__mux4_1_0.A3 0
C3639 a_16195_4585# a_8785_5039# 0.42059f
C3640 a_17125_4938# a_8785_5039# 0.31816f
C3641 VGND a_14297_5463# 0.67503f
C3642 w_14736_5374# a_13357_5719# 0
C3643 a_10569_1777# a_11553_1773# 0.08312f
C3644 VDPWR a_11986_4959# 0.02086f
C3645 a_7454_5039# w_7354_4954# 0.01793f
C3646 a_4837_16089# VGND 0.68517f
C3647 a_9477_11527# a_9589_12125# 0
C3648 a_11455_4959# VDPWR 0
C3649 a_9725_5837# a_10088_5837# 0.00847f
C3650 a_4910_5047# a_4159_5303# 0.00682f
C3651 a_11150_5467# a_11202_5441# 0.1439f
C3652 a_9547_16323# a_9799_16073# 0
C3653 a_4183_2153# a_4546_2153# 0.00847f
C3654 a_9467_13091# w_9492_12311# 0.0035f
C3655 a_6915_5043# w_5484_4958# 0.02026f
C3656 a_9699_4853# a_9585_4963# 0
C3657 a_11595_5833# w_11050_5382# 0
C3658 a_12509_4593# VGND 0.67184f
C3659 w_10748_13967# a_10813_13753# 0.08205f
C3660 a_15227_5715# sky130_fd_sc_hd__mux4_1_0.A3 0.00796f
C3661 a_9877_10533# a_12631_13987# 0.0762f
C3662 VDPWR a_9547_16323# 0.0251f
C3663 a_9809_14509# w_11718_13593# 0
C3664 a_12250_2139# VDPWR 0
C3665 a_14946_4905# a_13357_5719# 0
C3666 a_13271_4955# a_13046_4563# 0.00559f
C3667 a_2175_5417# VGND 0.0024f
C3668 a_9809_14509# a_11597_15219# 0.17824f
C3669 a_11569_4849# a_12320_4959# 0.00696f
C3670 w_12866_5378# a_12966_5463# 0.01793f
C3671 a_2313_2157# VDPWR 0.00745f
C3672 VDPWR a_6635_15235# 0.33595f
C3673 a_16195_4585# a_14916_4559# 0
C3674 a_23511_14335# ui_in[0] 0.01792f
C3675 a_5809_14763# a_5895_14763# 0.00658f
C3676 clk rst_n 0.03102f
C3677 a_11499_2029# a_10569_1777# 0.21188f
C3678 a_15255_4841# a_15309_4951# 0.03622f
C3679 a_9475_14759# w_9490_15543# 0
C3680 a_15672_4951# VDPWR 0.02182f
C3681 VGND w_9180_5386# 0.56712f
C3682 a_14836_5459# w_14736_5374# 0.01793f
C3683 a_6862_13645# a_6635_15235# 0
C3684 a_9867_12097# a_11243_11891# 0.03573f
C3685 a_13439_4955# a_13802_4955# 0.00847f
C3686 a_23731_14309# a_24152_14385# 0.01881f
C3687 w_14764_4500# a_15227_5715# 0
C3688 a_9587_15357# w_9392_16287# 0
C3689 a_24234_14385# sky130_fd_sc_hd__mux4_1_0.VPB 0.05795f
C3690 w_10674_14933# a_8113_13753# 0
C3691 a_5765_5043# a_6029_5043# 0
C3692 a_14975_2131# VDPWR 0
C3693 a_14846_1739# sky130_fd_sc_hd__mux4_1_0.A2 0.00279f
C3694 a_4755_12857# a_4839_12857# 0.00208f
C3695 a_9419_2143# a_9238_1777# 0
C3696 a_17125_4938# a_17346_5265# 0.00783f
C3697 a_4837_16089# a_5851_13769# 0.08387f
C3698 a_13732_2135# a_12439_1773# 0.03325f
C3699 a_11767_15219# a_11597_15219# 0.00167f
C3700 a_24241_14651# ui_in[1] 0.00168f
C3701 a_10965_11919# a_9867_12097# 0.18618f
C3702 w_14764_4500# sky130_fd_sc_hd__mux4_1_0.A3 0
C3703 a_11359_4593# VDPWR 0.00133f
C3704 a_13046_4563# sky130_fd_sc_hd__mux4_1_0.A3 0
C3705 a_9811_11277# w_10674_14933# 0.08584f
C3706 a_2313_1791# a_2049_1791# 0
C3707 a_14836_5459# a_14946_4905# 0.00175f
C3708 a_9875_13765# a_11089_13753# 0
C3709 VGND w_11718_13593# 0.01919f
C3710 VDPWR a_4915_10549# 0.69549f
C3711 a_9801_12841# a_10983_13753# 0
C3712 a_12924_1769# w_12824_1684# 0.01793f
C3713 a_9467_13091# a_9475_14759# 0
C3714 a_13243_5829# VGND 0.00268f
C3715 a_14325_4589# w_14736_5374# 0.00258f
C3716 VGND a_11597_15219# 0.13063f
C3717 a_14794_1765# sky130_fd_sc_hd__mux4_1_0.A2 0.00159f
C3718 a_24318_14385# a_24234_14385# 0.0296f
C3719 a_13439_4955# a_13175_4955# 0
C3720 a_8596_5405# VGND 0.00249f
C3721 a_14846_1739# VGND 0.40101f
C3722 VDPWR a_13357_5719# 0.3555f
C3723 a_6862_13645# a_4915_10549# 0
C3724 a_12509_4593# w_12894_4504# 0.24999f
C3725 a_5945_2039# sky130_fd_sc_hd__mux4_1_0.A2 0.00224f
C3726 a_14297_5463# a_8785_5039# 0.04835f
C3727 a_9629_2033# sky130_fd_sc_hd__mux4_1_0.A2 0.00296f
C3728 a_7476_1753# w_5454_1698# 0
C3729 a_23677_14335# sky130_fd_sc_hd__mux4_1_0.A3 0
C3730 a_12481_5467# w_11050_5382# 0.02004f
C3731 a_9238_1777# w_7324_1694# 0.00227f
C3732 w_5786_13983# a_6389_13769# 0.01492f
C3733 a_4503_16339# a_6629_15387# 0
C3734 VGND a_12809_13987# 0
C3735 a_9673_15357# a_9809_14509# 0
C3736 a_12135_15219# a_12075_13379# 0.36868f
C3737 w_10748_13967# a_10771_14747# 0
C3738 a_5636_5017# a_6029_5409# 0.02301f
C3739 ua[1] sky130_fd_sc_hd__mux4_1_0.VNB 0.14696f
C3740 ua[2] sky130_fd_sc_hd__mux4_1_0.VNB 0.14696f
C3741 ua[3] sky130_fd_sc_hd__mux4_1_0.VNB 0.14696f
C3742 ua[4] sky130_fd_sc_hd__mux4_1_0.VNB 0.14465f
C3743 ua[5] sky130_fd_sc_hd__mux4_1_0.VNB 0.14471f
C3744 ua[6] sky130_fd_sc_hd__mux4_1_0.VNB 0.14538f
C3745 ua[7] sky130_fd_sc_hd__mux4_1_0.VNB 0.1455f
C3746 ena sky130_fd_sc_hd__mux4_1_0.VNB 0.07038f
C3747 clk sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3748 rst_n sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3749 ui_in[2] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3750 ui_in[3] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3751 ui_in[4] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3752 ui_in[5] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3753 ui_in[6] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3754 ui_in[7] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3755 uio_in[0] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3756 uio_in[1] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3757 uio_in[2] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3758 uio_in[3] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3759 uio_in[4] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3760 uio_in[5] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3761 uio_in[6] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3762 uio_in[7] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3763 uo_out[0] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3764 uo_out[1] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3765 uo_out[2] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3766 uo_out[3] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3767 uo_out[4] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3768 uo_out[5] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3769 uo_out[6] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3770 uo_out[7] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3771 uio_out[0] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3772 uio_out[1] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3773 uio_out[2] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3774 uio_out[3] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3775 uio_out[4] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3776 uio_out[5] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3777 uio_out[6] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3778 uio_out[7] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3779 uio_oe[0] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3780 uio_oe[1] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3781 uio_oe[2] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3782 uio_oe[3] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3783 uio_oe[4] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3784 uio_oe[5] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3785 uio_oe[6] sky130_fd_sc_hd__mux4_1_0.VNB 0.04288f
C3786 uio_oe[7] sky130_fd_sc_hd__mux4_1_0.VNB 0.07038f
C3787 ua[0] sky130_fd_sc_hd__mux4_1_0.VNB 9.60658f
C3788 ui_in[1] sky130_fd_sc_hd__mux4_1_0.VNB 8.61396f
C3789 ui_in[0] sky130_fd_sc_hd__mux4_1_0.VNB 9.30023f
C3790 VDPWR sky130_fd_sc_hd__mux4_1_0.VNB 81.6264f
C3791 VGND sky130_fd_sc_hd__mux4_1_0.VNB 95.02061f
C3792 a_15602_1765# sky130_fd_sc_hd__mux4_1_0.VNB 0.00345f
C3793 a_15239_1765# sky130_fd_sc_hd__mux4_1_0.VNB 0.00484f
C3794 a_13732_1769# sky130_fd_sc_hd__mux4_1_0.VNB 0.00345f
C3795 a_13369_1769# sky130_fd_sc_hd__mux4_1_0.VNB 0.00484f
C3796 a_15602_2131# sky130_fd_sc_hd__mux4_1_0.VNB 0.01578f
C3797 a_15239_2131# sky130_fd_sc_hd__mux4_1_0.VNB 0.01584f
C3798 a_14794_1765# sky130_fd_sc_hd__mux4_1_0.VNB 0.06682f
C3799 a_15185_2021# sky130_fd_sc_hd__mux4_1_0.VNB 0.27343f
C3800 a_14846_1739# sky130_fd_sc_hd__mux4_1_0.VNB 0.13081f
C3801 a_14255_1769# sky130_fd_sc_hd__mux4_1_0.VNB 0.55211f
C3802 a_11916_1773# sky130_fd_sc_hd__mux4_1_0.VNB 0.00345f
C3803 a_11553_1773# sky130_fd_sc_hd__mux4_1_0.VNB 0.00484f
C3804 a_13732_2135# sky130_fd_sc_hd__mux4_1_0.VNB 0.01578f
C3805 a_13369_2135# sky130_fd_sc_hd__mux4_1_0.VNB 0.01584f
C3806 a_12924_1769# sky130_fd_sc_hd__mux4_1_0.VNB 0.06298f
C3807 a_13315_2025# sky130_fd_sc_hd__mux4_1_0.VNB 0.26543f
C3808 a_12976_1743# sky130_fd_sc_hd__mux4_1_0.VNB 0.13025f
C3809 a_12439_1773# sky130_fd_sc_hd__mux4_1_0.VNB 0.52339f
C3810 a_10046_1777# sky130_fd_sc_hd__mux4_1_0.VNB 0.00345f
C3811 a_9683_1777# sky130_fd_sc_hd__mux4_1_0.VNB 0.00484f
C3812 a_11916_2139# sky130_fd_sc_hd__mux4_1_0.VNB 0.01578f
C3813 a_11553_2139# sky130_fd_sc_hd__mux4_1_0.VNB 0.01584f
C3814 a_11108_1773# sky130_fd_sc_hd__mux4_1_0.VNB 0.06682f
C3815 a_11499_2029# sky130_fd_sc_hd__mux4_1_0.VNB 0.26466f
C3816 a_11160_1747# sky130_fd_sc_hd__mux4_1_0.VNB 0.13081f
C3817 a_10569_1777# sky130_fd_sc_hd__mux4_1_0.VNB 0.55211f
C3818 a_8232_1779# sky130_fd_sc_hd__mux4_1_0.VNB 0.00345f
C3819 a_7869_1779# sky130_fd_sc_hd__mux4_1_0.VNB 0.00484f
C3820 a_10046_2143# sky130_fd_sc_hd__mux4_1_0.VNB 0.01578f
C3821 a_9683_2143# sky130_fd_sc_hd__mux4_1_0.VNB 0.01584f
C3822 a_9238_1777# sky130_fd_sc_hd__mux4_1_0.VNB 0.06285f
C3823 a_9629_2033# sky130_fd_sc_hd__mux4_1_0.VNB 0.26543f
C3824 a_9290_1751# sky130_fd_sc_hd__mux4_1_0.VNB 0.13016f
C3825 a_8755_1779# sky130_fd_sc_hd__mux4_1_0.VNB 0.52093f
C3826 a_6362_1783# sky130_fd_sc_hd__mux4_1_0.VNB 0.00345f
C3827 a_5999_1783# sky130_fd_sc_hd__mux4_1_0.VNB 0.00484f
C3828 a_8232_2145# sky130_fd_sc_hd__mux4_1_0.VNB 0.01578f
C3829 a_7869_2145# sky130_fd_sc_hd__mux4_1_0.VNB 0.01584f
C3830 a_7424_1779# sky130_fd_sc_hd__mux4_1_0.VNB 0.06682f
C3831 a_7815_2035# sky130_fd_sc_hd__mux4_1_0.VNB 0.26452f
C3832 a_7476_1753# sky130_fd_sc_hd__mux4_1_0.VNB 0.13081f
C3833 a_6885_1783# sky130_fd_sc_hd__mux4_1_0.VNB 0.55211f
C3834 a_4546_1787# sky130_fd_sc_hd__mux4_1_0.VNB 0.00345f
C3835 a_4183_1787# sky130_fd_sc_hd__mux4_1_0.VNB 0.00484f
C3836 a_6362_2149# sky130_fd_sc_hd__mux4_1_0.VNB 0.01578f
C3837 a_5999_2149# sky130_fd_sc_hd__mux4_1_0.VNB 0.01584f
C3838 a_5554_1783# sky130_fd_sc_hd__mux4_1_0.VNB 0.06298f
C3839 a_5945_2039# sky130_fd_sc_hd__mux4_1_0.VNB 0.26543f
C3840 a_5606_1757# sky130_fd_sc_hd__mux4_1_0.VNB 0.13025f
C3841 a_5069_1787# sky130_fd_sc_hd__mux4_1_0.VNB 0.52277f
C3842 a_2676_1791# sky130_fd_sc_hd__mux4_1_0.VNB 0.00345f
C3843 a_2313_1791# sky130_fd_sc_hd__mux4_1_0.VNB 0.00484f
C3844 a_4546_2153# sky130_fd_sc_hd__mux4_1_0.VNB 0.01578f
C3845 a_4183_2153# sky130_fd_sc_hd__mux4_1_0.VNB 0.01584f
C3846 a_3738_1787# sky130_fd_sc_hd__mux4_1_0.VNB 0.06682f
C3847 a_4129_2043# sky130_fd_sc_hd__mux4_1_0.VNB 0.26466f
C3848 a_3790_1761# sky130_fd_sc_hd__mux4_1_0.VNB 0.13081f
C3849 a_3199_1791# sky130_fd_sc_hd__mux4_1_0.VNB 0.55211f
C3850 a_2676_2157# sky130_fd_sc_hd__mux4_1_0.VNB 0.01578f
C3851 a_2313_2157# sky130_fd_sc_hd__mux4_1_0.VNB 0.01584f
C3852 a_1868_1791# sky130_fd_sc_hd__mux4_1_0.VNB 0.10031f
C3853 a_2259_2047# sky130_fd_sc_hd__mux4_1_0.VNB 0.26543f
C3854 a_1920_1765# sky130_fd_sc_hd__mux4_1_0.VNB 0.1359f
C3855 a_2187_1765# sky130_fd_sc_hd__mux4_1_0.VNB 2.28963f
C3856 a_15672_4585# sky130_fd_sc_hd__mux4_1_0.VNB 0.00345f
C3857 a_15309_4585# sky130_fd_sc_hd__mux4_1_0.VNB 0.00484f
C3858 a_13802_4589# sky130_fd_sc_hd__mux4_1_0.VNB 0.00345f
C3859 a_13439_4589# sky130_fd_sc_hd__mux4_1_0.VNB 0.00484f
C3860 a_15672_4951# sky130_fd_sc_hd__mux4_1_0.VNB 0.01578f
C3861 a_15309_4951# sky130_fd_sc_hd__mux4_1_0.VNB 0.01584f
C3862 a_14864_4585# sky130_fd_sc_hd__mux4_1_0.VNB 0.06682f
C3863 a_15255_4841# sky130_fd_sc_hd__mux4_1_0.VNB 0.26397f
C3864 a_14946_4905# sky130_fd_sc_hd__mux4_1_0.VNB 1.04897f
C3865 a_14916_4559# sky130_fd_sc_hd__mux4_1_0.VNB 0.12906f
C3866 a_14325_4589# sky130_fd_sc_hd__mux4_1_0.VNB 0.51247f
C3867 a_11986_4593# sky130_fd_sc_hd__mux4_1_0.VNB 0.00345f
C3868 a_11623_4593# sky130_fd_sc_hd__mux4_1_0.VNB 0.00484f
C3869 a_13802_4955# sky130_fd_sc_hd__mux4_1_0.VNB 0.01578f
C3870 a_13439_4955# sky130_fd_sc_hd__mux4_1_0.VNB 0.01584f
C3871 a_12994_4589# sky130_fd_sc_hd__mux4_1_0.VNB 0.06298f
C3872 a_13385_4845# sky130_fd_sc_hd__mux4_1_0.VNB 0.26214f
C3873 a_13046_4563# sky130_fd_sc_hd__mux4_1_0.VNB 0.12849f
C3874 a_12509_4593# sky130_fd_sc_hd__mux4_1_0.VNB 0.48861f
C3875 a_10116_4597# sky130_fd_sc_hd__mux4_1_0.VNB 0.00345f
C3876 a_9753_4597# sky130_fd_sc_hd__mux4_1_0.VNB 0.00484f
C3877 a_11986_4959# sky130_fd_sc_hd__mux4_1_0.VNB 0.01578f
C3878 a_11623_4959# sky130_fd_sc_hd__mux4_1_0.VNB 0.01584f
C3879 a_11178_4593# sky130_fd_sc_hd__mux4_1_0.VNB 0.06682f
C3880 a_11569_4849# sky130_fd_sc_hd__mux4_1_0.VNB 0.26136f
C3881 a_11230_4567# sky130_fd_sc_hd__mux4_1_0.VNB 0.12906f
C3882 a_10639_4597# sky130_fd_sc_hd__mux4_1_0.VNB 0.51206f
C3883 a_10116_4963# sky130_fd_sc_hd__mux4_1_0.VNB 0.01578f
C3884 a_9753_4963# sky130_fd_sc_hd__mux4_1_0.VNB 0.01584f
C3885 a_9308_4597# sky130_fd_sc_hd__mux4_1_0.VNB 0.09346f
C3886 a_9699_4853# sky130_fd_sc_hd__mux4_1_0.VNB 0.26214f
C3887 a_9360_4571# sky130_fd_sc_hd__mux4_1_0.VNB 0.13349f
C3888 a_8262_5039# sky130_fd_sc_hd__mux4_1_0.VNB 0.00345f
C3889 a_7899_5039# sky130_fd_sc_hd__mux4_1_0.VNB 0.00484f
C3890 a_17125_4938# sky130_fd_sc_hd__mux4_1_0.VNB 0.13914f
C3891 a_16195_4585# sky130_fd_sc_hd__mux4_1_0.VNB 0.44799f
C3892 a_16871_4938# sky130_fd_sc_hd__mux4_1_0.VNB 0.23758f
C3893 a_15644_5459# sky130_fd_sc_hd__mux4_1_0.VNB 0.00345f
C3894 a_15281_5459# sky130_fd_sc_hd__mux4_1_0.VNB 0.00484f
C3895 a_16167_5459# sky130_fd_sc_hd__mux4_1_0.VNB 0.5186f
C3896 a_13774_5463# sky130_fd_sc_hd__mux4_1_0.VNB 0.00345f
C3897 a_13411_5463# sky130_fd_sc_hd__mux4_1_0.VNB 0.00484f
C3898 a_15644_5825# sky130_fd_sc_hd__mux4_1_0.VNB 0.01578f
C3899 a_15281_5825# sky130_fd_sc_hd__mux4_1_0.VNB 0.01584f
C3900 a_14836_5459# sky130_fd_sc_hd__mux4_1_0.VNB 0.06682f
C3901 a_15227_5715# sky130_fd_sc_hd__mux4_1_0.VNB 0.27134f
C3902 a_14888_5433# sky130_fd_sc_hd__mux4_1_0.VNB 0.12984f
C3903 a_14297_5463# sky130_fd_sc_hd__mux4_1_0.VNB 0.50345f
C3904 a_11958_5467# sky130_fd_sc_hd__mux4_1_0.VNB 0.00345f
C3905 a_11595_5467# sky130_fd_sc_hd__mux4_1_0.VNB 0.00484f
C3906 a_13774_5829# sky130_fd_sc_hd__mux4_1_0.VNB 0.01578f
C3907 a_13411_5829# sky130_fd_sc_hd__mux4_1_0.VNB 0.01584f
C3908 a_12966_5463# sky130_fd_sc_hd__mux4_1_0.VNB 0.06298f
C3909 a_13357_5719# sky130_fd_sc_hd__mux4_1_0.VNB 0.26335f
C3910 a_13018_5437# sky130_fd_sc_hd__mux4_1_0.VNB 0.12928f
C3911 a_12481_5467# sky130_fd_sc_hd__mux4_1_0.VNB 0.48206f
C3912 a_10088_5471# sky130_fd_sc_hd__mux4_1_0.VNB 0.00345f
C3913 a_9725_5471# sky130_fd_sc_hd__mux4_1_0.VNB 0.00484f
C3914 a_11958_5833# sky130_fd_sc_hd__mux4_1_0.VNB 0.01578f
C3915 a_11595_5833# sky130_fd_sc_hd__mux4_1_0.VNB 0.01584f
C3916 a_11150_5467# sky130_fd_sc_hd__mux4_1_0.VNB 0.06682f
C3917 a_11541_5723# sky130_fd_sc_hd__mux4_1_0.VNB 0.26257f
C3918 a_11202_5441# sky130_fd_sc_hd__mux4_1_0.VNB 0.12984f
C3919 a_10611_5471# sky130_fd_sc_hd__mux4_1_0.VNB 0.50409f
C3920 a_8785_5039# sky130_fd_sc_hd__mux4_1_0.VNB 1.40108f
C3921 a_6392_5043# sky130_fd_sc_hd__mux4_1_0.VNB 0.00345f
C3922 a_6029_5043# sky130_fd_sc_hd__mux4_1_0.VNB 0.00484f
C3923 a_8262_5405# sky130_fd_sc_hd__mux4_1_0.VNB 0.01578f
C3924 a_7899_5405# sky130_fd_sc_hd__mux4_1_0.VNB 0.01584f
C3925 a_7454_5039# sky130_fd_sc_hd__mux4_1_0.VNB 0.06682f
C3926 a_7845_5295# sky130_fd_sc_hd__mux4_1_0.VNB 0.27171f
C3927 a_7506_5013# sky130_fd_sc_hd__mux4_1_0.VNB 0.13081f
C3928 a_6915_5043# sky130_fd_sc_hd__mux4_1_0.VNB 0.55211f
C3929 a_4576_5047# sky130_fd_sc_hd__mux4_1_0.VNB 0.00345f
C3930 a_4213_5047# sky130_fd_sc_hd__mux4_1_0.VNB 0.00484f
C3931 a_6392_5409# sky130_fd_sc_hd__mux4_1_0.VNB 0.01578f
C3932 a_6029_5409# sky130_fd_sc_hd__mux4_1_0.VNB 0.01584f
C3933 a_5584_5043# sky130_fd_sc_hd__mux4_1_0.VNB 0.06298f
C3934 a_5975_5299# sky130_fd_sc_hd__mux4_1_0.VNB 0.26543f
C3935 a_5636_5017# sky130_fd_sc_hd__mux4_1_0.VNB 0.13025f
C3936 a_5099_5047# sky130_fd_sc_hd__mux4_1_0.VNB 0.52543f
C3937 a_2706_5051# sky130_fd_sc_hd__mux4_1_0.VNB 0.00345f
C3938 a_2343_5051# sky130_fd_sc_hd__mux4_1_0.VNB 0.00484f
C3939 a_4576_5413# sky130_fd_sc_hd__mux4_1_0.VNB 0.01578f
C3940 a_4213_5413# sky130_fd_sc_hd__mux4_1_0.VNB 0.01584f
C3941 a_3768_5047# sky130_fd_sc_hd__mux4_1_0.VNB 0.06682f
C3942 a_4159_5303# sky130_fd_sc_hd__mux4_1_0.VNB 0.26466f
C3943 a_3820_5021# sky130_fd_sc_hd__mux4_1_0.VNB 0.13081f
C3944 a_3229_5051# sky130_fd_sc_hd__mux4_1_0.VNB 0.55211f
C3945 a_2706_5417# sky130_fd_sc_hd__mux4_1_0.VNB 0.01578f
C3946 a_2343_5417# sky130_fd_sc_hd__mux4_1_0.VNB 0.01584f
C3947 a_1898_5051# sky130_fd_sc_hd__mux4_1_0.VNB 0.10031f
C3948 a_2289_5307# sky130_fd_sc_hd__mux4_1_0.VNB 0.26543f
C3949 a_1950_5025# sky130_fd_sc_hd__mux4_1_0.VNB 0.1359f
C3950 a_10088_5837# sky130_fd_sc_hd__mux4_1_0.VNB 0.01578f
C3951 a_9725_5837# sky130_fd_sc_hd__mux4_1_0.VNB 0.01584f
C3952 a_9280_5471# sky130_fd_sc_hd__mux4_1_0.VNB 0.09442f
C3953 a_9671_5727# sky130_fd_sc_hd__mux4_1_0.VNB 0.26335f
C3954 a_9332_5445# sky130_fd_sc_hd__mux4_1_0.VNB 0.13493f
C3955 a_2217_5025# sky130_fd_sc_hd__mux4_1_0.VNB 2.29089f
C3956 a_9599_10561# sky130_fd_sc_hd__mux4_1_0.VNB 0.1752f
C3957 a_4637_10577# sky130_fd_sc_hd__mux4_1_0.VNB 0.1752f
C3958 a_9727_11527# sky130_fd_sc_hd__mux4_1_0.VNB 0.00137f
C3959 a_9477_11527# sky130_fd_sc_hd__mux4_1_0.VNB 0.24712f
C3960 a_4765_11543# sky130_fd_sc_hd__mux4_1_0.VNB 0.00137f
C3961 a_4515_11543# sky130_fd_sc_hd__mux4_1_0.VNB 0.24712f
C3962 a_10965_11919# sky130_fd_sc_hd__mux4_1_0.VNB 0.1732f
C3963 a_9867_12097# sky130_fd_sc_hd__mux4_1_0.VNB 0.54635f
C3964 a_6003_11935# sky130_fd_sc_hd__mux4_1_0.VNB 0.1732f
C3965 a_9589_12125# sky130_fd_sc_hd__mux4_1_0.VNB 0.17114f
C3966 a_4905_12113# sky130_fd_sc_hd__mux4_1_0.VNB 0.55094f
C3967 a_4627_12141# sky130_fd_sc_hd__mux4_1_0.VNB 0.17114f
C3968 a_9717_13091# sky130_fd_sc_hd__mux4_1_0.VNB 0.00137f
C3969 a_9467_13091# sky130_fd_sc_hd__mux4_1_0.VNB 0.24424f
C3970 a_10937_12911# sky130_fd_sc_hd__mux4_1_0.VNB 0.16539f
C3971 a_4755_13107# sky130_fd_sc_hd__mux4_1_0.VNB 0.00137f
C3972 a_4505_13107# sky130_fd_sc_hd__mux4_1_0.VNB 0.24424f
C3973 a_5975_12927# sky130_fd_sc_hd__mux4_1_0.VNB 0.16539f
C3974 a_11291_12911# sky130_fd_sc_hd__mux4_1_0.VNB 0.46058f
C3975 a_11824_13629# sky130_fd_sc_hd__mux4_1_0.VNB 0.1516f
C3976 a_12075_13379# sky130_fd_sc_hd__mux4_1_0.VNB 0.40216f
C3977 a_11243_11891# sky130_fd_sc_hd__mux4_1_0.VNB 1.12822f
C3978 a_9877_10533# sky130_fd_sc_hd__mux4_1_0.VNB 3.44942f
C3979 a_12631_13987# sky130_fd_sc_hd__mux4_1_0.VNB 0.15779f
C3980 a_11351_13753# sky130_fd_sc_hd__mux4_1_0.VNB 0.31965f
C3981 a_10813_13753# sky130_fd_sc_hd__mux4_1_0.VNB 0.16387f
C3982 a_9875_13765# sky130_fd_sc_hd__mux4_1_0.VNB 0.45251f
C3983 a_6329_12927# sky130_fd_sc_hd__mux4_1_0.VNB 0.46058f
C3984 a_6862_13645# sky130_fd_sc_hd__mux4_1_0.VNB 0.1516f
C3985 a_7113_13395# sky130_fd_sc_hd__mux4_1_0.VNB 0.39872f
C3986 a_6281_11907# sky130_fd_sc_hd__mux4_1_0.VNB 1.1397f
C3987 a_4915_10549# sky130_fd_sc_hd__mux4_1_0.VNB 3.27518f
C3988 a_9597_13793# sky130_fd_sc_hd__mux4_1_0.VNB 0.16601f
C3989 a_7669_14003# sky130_fd_sc_hd__mux4_1_0.VNB 0.1564f
C3990 a_6389_13769# sky130_fd_sc_hd__mux4_1_0.VNB 0.31965f
C3991 a_5851_13769# sky130_fd_sc_hd__mux4_1_0.VNB 0.16387f
C3992 a_4913_13781# sky130_fd_sc_hd__mux4_1_0.VNB 0.45689f
C3993 a_4635_13809# sky130_fd_sc_hd__mux4_1_0.VNB 0.17003f
C3994 a_24318_14385# sky130_fd_sc_hd__mux4_1_0.VNB 0.02499f
C3995 a_24152_14385# sky130_fd_sc_hd__mux4_1_0.VNB 0.02039f
C3996 a_23511_14335# sky130_fd_sc_hd__mux4_1_0.VNB 0.04207f
C3997 a_24962_14701# sky130_fd_sc_hd__mux4_1_0.VNB 0.16413f
C3998 a_24774_14701# sky130_fd_sc_hd__mux4_1_0.VNB 0.2179f
C3999 a_24234_14385# sky130_fd_sc_hd__mux4_1_0.VNB 0.03874f
C4000 a_24241_14651# sky130_fd_sc_hd__mux4_1_0.VNB 0.00666f
C4001 sky130_fd_sc_hd__mux4_1_0.A2 sky130_fd_sc_hd__mux4_1_0.VNB 11.8725f
C4002 sky130_fd_sc_hd__mux4_1_0.A3 sky130_fd_sc_hd__mux4_1_0.VNB 10.095f
C4003 a_23731_14309# sky130_fd_sc_hd__mux4_1_0.VNB 0.33779f
C4004 a_23677_14701# sky130_fd_sc_hd__mux4_1_0.VNB 0.00373f
C4005 a_23511_14701# sky130_fd_sc_hd__mux4_1_0.VNB 0.02865f
C4006 a_9725_14759# sky130_fd_sc_hd__mux4_1_0.VNB 0.00137f
C4007 a_9475_14759# sky130_fd_sc_hd__mux4_1_0.VNB 0.24496f
C4008 a_9801_12841# sky130_fd_sc_hd__mux4_1_0.VNB 1.33033f
C4009 a_9811_11277# sky130_fd_sc_hd__mux4_1_0.VNB 2.17869f
C4010 a_10771_14747# sky130_fd_sc_hd__mux4_1_0.VNB 0.1671f
C4011 a_4763_14775# sky130_fd_sc_hd__mux4_1_0.VNB 0.00137f
C4012 a_4513_14775# sky130_fd_sc_hd__mux4_1_0.VNB 0.24496f
C4013 a_4839_12857# sky130_fd_sc_hd__mux4_1_0.VNB 1.33478f
C4014 a_4849_11293# sky130_fd_sc_hd__mux4_1_0.VNB 2.17869f
C4015 a_5809_14763# sky130_fd_sc_hd__mux4_1_0.VNB 0.1671f
C4016 a_12135_15219# sky130_fd_sc_hd__mux4_1_0.VNB 0.75127f
C4017 a_11597_15219# sky130_fd_sc_hd__mux4_1_0.VNB 0.17279f
C4018 a_11049_14719# sky130_fd_sc_hd__mux4_1_0.VNB 0.33714f
C4019 a_9809_14509# sky130_fd_sc_hd__mux4_1_0.VNB 0.62284f
C4020 a_8113_13753# sky130_fd_sc_hd__mux4_1_0.VNB 3.07869f
C4021 a_9865_15329# sky130_fd_sc_hd__mux4_1_0.VNB 0.69482f
C4022 a_7173_15235# sky130_fd_sc_hd__mux4_1_0.VNB 0.79677f
C4023 a_6635_15235# sky130_fd_sc_hd__mux4_1_0.VNB 0.17279f
C4024 a_6087_14735# sky130_fd_sc_hd__mux4_1_0.VNB 0.33714f
C4025 a_4847_14525# sky130_fd_sc_hd__mux4_1_0.VNB 0.63122f
C4026 a_9587_15357# sky130_fd_sc_hd__mux4_1_0.VNB 0.17275f
C4027 a_4903_15345# sky130_fd_sc_hd__mux4_1_0.VNB 0.69937f
C4028 a_4625_15373# sky130_fd_sc_hd__mux4_1_0.VNB 0.17275f
C4029 a_22274_16171# sky130_fd_sc_hd__mux4_1_0.VNB 0.45419f
C4030 a_21506_16181# sky130_fd_sc_hd__mux4_1_0.VNB 0.40241f
C4031 a_20384_16179# sky130_fd_sc_hd__mux4_1_0.VNB 0.53611f
C4032 a_19510_16177# sky130_fd_sc_hd__mux4_1_0.VNB 0.45443f
C4033 a_18742_16187# sky130_fd_sc_hd__mux4_1_0.VNB 0.40031f
C4034 a_18128_16189# sky130_fd_sc_hd__mux4_1_0.VNB 0.33935f
C4035 a_17254_16187# sky130_fd_sc_hd__mux4_1_0.VNB 0.45045f
C4036 a_16486_16197# sky130_fd_sc_hd__mux4_1_0.VNB 0.40469f
C4037 a_9799_16073# sky130_fd_sc_hd__mux4_1_0.VNB 1.62449f
C4038 a_9715_16323# sky130_fd_sc_hd__mux4_1_0.VNB 0.00137f
C4039 a_9465_16323# sky130_fd_sc_hd__mux4_1_0.VNB 0.24845f
C4040 a_4837_16089# sky130_fd_sc_hd__mux4_1_0.VNB 1.72323f
C4041 a_4753_16339# sky130_fd_sc_hd__mux4_1_0.VNB 0.00137f
C4042 a_4503_16339# sky130_fd_sc_hd__mux4_1_0.VNB 0.24845f
C4043 sky130_fd_sc_hd__mux4_1_0.A0 sky130_fd_sc_hd__mux4_1_0.VNB 3.82953f
C4044 a_6629_15387# sky130_fd_sc_hd__mux4_1_0.VNB 2.47775f
C4045 sky130_fd_sc_hd__mux4_1_0.A1 sky130_fd_sc_hd__mux4_1_0.VNB 8.29901f
C4046 w_14694_1680# sky130_fd_sc_hd__mux4_1_0.VNB 1.49072f
C4047 w_12824_1684# sky130_fd_sc_hd__mux4_1_0.VNB 1.49072f
C4048 w_11008_1688# sky130_fd_sc_hd__mux4_1_0.VNB 1.49072f
C4049 w_9138_1692# sky130_fd_sc_hd__mux4_1_0.VNB 1.49072f
C4050 w_7324_1694# sky130_fd_sc_hd__mux4_1_0.VNB 1.49072f
C4051 w_5454_1698# sky130_fd_sc_hd__mux4_1_0.VNB 1.49072f
C4052 w_3638_1702# sky130_fd_sc_hd__mux4_1_0.VNB 1.49072f
C4053 w_1768_1706# sky130_fd_sc_hd__mux4_1_0.VNB 1.49072f
C4054 w_6044_2758# sky130_fd_sc_hd__mux4_1_0.VNB 0.33898f
C4055 w_16764_4814# sky130_fd_sc_hd__mux4_1_0.VNB 0.87055f
C4056 w_14764_4500# sky130_fd_sc_hd__mux4_1_0.VNB 1.49072f
C4057 w_12894_4504# sky130_fd_sc_hd__mux4_1_0.VNB 1.49072f
C4058 w_11078_4508# sky130_fd_sc_hd__mux4_1_0.VNB 1.49072f
C4059 w_9208_4512# sky130_fd_sc_hd__mux4_1_0.VNB 1.49072f
C4060 w_7354_4954# sky130_fd_sc_hd__mux4_1_0.VNB 1.49072f
C4061 w_5484_4958# sky130_fd_sc_hd__mux4_1_0.VNB 1.49072f
C4062 w_3668_4962# sky130_fd_sc_hd__mux4_1_0.VNB 1.49072f
C4063 w_1798_4966# sky130_fd_sc_hd__mux4_1_0.VNB 1.49072f
C4064 w_14736_5374# sky130_fd_sc_hd__mux4_1_0.VNB 1.49072f
C4065 w_12866_5378# sky130_fd_sc_hd__mux4_1_0.VNB 1.49072f
C4066 w_11050_5382# sky130_fd_sc_hd__mux4_1_0.VNB 1.49072f
C4067 w_9180_5386# sky130_fd_sc_hd__mux4_1_0.VNB 1.49072f
C4068 w_6074_6018# sky130_fd_sc_hd__mux4_1_0.VNB 0.33898f
C4069 w_9502_10747# sky130_fd_sc_hd__mux4_1_0.VNB 0.51617f
C4070 w_4540_10763# sky130_fd_sc_hd__mux4_1_0.VNB 0.51617f
C4071 w_9404_11491# sky130_fd_sc_hd__mux4_1_0.VNB 0.69336f
C4072 w_4442_11507# sky130_fd_sc_hd__mux4_1_0.VNB 0.69336f
C4073 w_10868_12105# sky130_fd_sc_hd__mux4_1_0.VNB 0.51617f
C4074 w_9492_12311# sky130_fd_sc_hd__mux4_1_0.VNB 0.51617f
C4075 w_5906_12121# sky130_fd_sc_hd__mux4_1_0.VNB 0.51617f
C4076 w_4530_12327# sky130_fd_sc_hd__mux4_1_0.VNB 0.51617f
C4077 w_10872_13125# sky130_fd_sc_hd__mux4_1_0.VNB 0.51617f
C4078 w_9394_13055# sky130_fd_sc_hd__mux4_1_0.VNB 0.69336f
C4079 w_5910_13141# sky130_fd_sc_hd__mux4_1_0.VNB 0.51617f
C4080 w_4432_13071# sky130_fd_sc_hd__mux4_1_0.VNB 0.69336f
C4081 w_11718_13593# sky130_fd_sc_hd__mux4_1_0.VNB 0.51617f
C4082 w_6756_13609# sky130_fd_sc_hd__mux4_1_0.VNB 0.51617f
C4083 w_12566_13951# sky130_fd_sc_hd__mux4_1_0.VNB 0.60476f
C4084 w_10748_13967# sky130_fd_sc_hd__mux4_1_0.VNB 0.69336f
C4085 w_9500_13979# sky130_fd_sc_hd__mux4_1_0.VNB 0.51617f
C4086 w_7604_13967# sky130_fd_sc_hd__mux4_1_0.VNB 0.60476f
C4087 w_5786_13983# sky130_fd_sc_hd__mux4_1_0.VNB 0.69336f
C4088 w_4538_13995# sky130_fd_sc_hd__mux4_1_0.VNB 0.51617f
C4089 sky130_fd_sc_hd__mux4_1_0.VPB sky130_fd_sc_hd__mux4_1_0.VNB 1.9337f
C4090 w_10674_14933# sky130_fd_sc_hd__mux4_1_0.VNB 0.51617f
C4091 w_9402_14723# sky130_fd_sc_hd__mux4_1_0.VNB 0.69336f
C4092 w_5712_14949# sky130_fd_sc_hd__mux4_1_0.VNB 0.51617f
C4093 w_4440_14739# sky130_fd_sc_hd__mux4_1_0.VNB 0.69336f
C4094 w_11532_15433# sky130_fd_sc_hd__mux4_1_0.VNB 0.69336f
C4095 w_9490_15543# sky130_fd_sc_hd__mux4_1_0.VNB 0.51617f
C4096 w_6570_15449# sky130_fd_sc_hd__mux4_1_0.VNB 0.69336f
C4097 w_4528_15559# sky130_fd_sc_hd__mux4_1_0.VNB 0.51617f
C4098 w_22960_16387# sky130_fd_sc_hd__mux4_1_0.VNB 0.33898f
C4099 w_22086_16385# sky130_fd_sc_hd__mux4_1_0.VNB 0.33898f
C4100 w_21318_16395# sky130_fd_sc_hd__mux4_1_0.VNB 0.33898f
C4101 w_20196_16393# sky130_fd_sc_hd__mux4_1_0.VNB 0.33898f
C4102 w_19322_16391# sky130_fd_sc_hd__mux4_1_0.VNB 0.33898f
C4103 w_18554_16401# sky130_fd_sc_hd__mux4_1_0.VNB 0.33898f
C4104 w_17940_16403# sky130_fd_sc_hd__mux4_1_0.VNB 0.33898f
C4105 w_17066_16401# sky130_fd_sc_hd__mux4_1_0.VNB 0.33898f
C4106 w_16298_16411# sky130_fd_sc_hd__mux4_1_0.VNB 0.33898f
C4107 w_9392_16287# sky130_fd_sc_hd__mux4_1_0.VNB 0.69336f
C4108 w_4430_16303# sky130_fd_sc_hd__mux4_1_0.VNB 0.69336f
C4109 w_9392_17212# sky130_fd_sc_hd__mux4_1_0.VNB 0.33898f
.ends

