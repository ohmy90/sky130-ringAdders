VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_ohmy90_adders
  CLASS BLOCK ;
  FOREIGN tt_um_ohmy90_adders ;
  ORIGIN -0.990 0.000 ;
  SIZE 151.720 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.378000 ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.252000 ;
    ANTENNADIFFAREA 0.502250 ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 48.215 88.885 48.385 89.055 ;
        RECT 48.215 88.865 48.320 88.885 ;
        RECT 47.390 87.955 48.320 88.865 ;
      LAYER nwell ;
        RECT 46.960 86.060 48.720 87.665 ;
        RECT 22.150 81.515 25.750 83.120 ;
        RECT 46.960 81.435 50.560 83.040 ;
        RECT 81.490 82.055 83.250 83.660 ;
        RECT 85.330 82.005 87.090 83.610 ;
        RECT 89.700 82.015 91.460 83.620 ;
        RECT 92.770 82.005 94.530 83.610 ;
        RECT 96.610 81.955 98.370 83.560 ;
        RECT 100.980 81.965 102.740 83.570 ;
        RECT 106.590 81.975 108.350 83.580 ;
        RECT 110.430 81.925 112.190 83.530 ;
        RECT 114.800 81.935 116.560 83.540 ;
      LAYER pwell ;
        RECT 22.385 80.315 25.555 81.225 ;
        RECT 22.485 80.125 22.655 80.315 ;
        RECT 47.195 80.235 50.365 81.145 ;
        RECT 81.890 80.855 82.820 81.765 ;
        RECT 81.890 80.835 81.995 80.855 ;
        RECT 81.825 80.665 81.995 80.835 ;
        RECT 85.730 80.805 86.660 81.715 ;
        RECT 90.100 80.815 91.030 81.725 ;
        RECT 85.730 80.785 85.835 80.805 ;
        RECT 90.100 80.795 90.205 80.815 ;
        RECT 85.665 80.615 85.835 80.785 ;
        RECT 90.035 80.625 90.205 80.795 ;
        RECT 93.170 80.805 94.100 81.715 ;
        RECT 93.170 80.785 93.275 80.805 ;
        RECT 93.105 80.615 93.275 80.785 ;
        RECT 97.010 80.755 97.940 81.665 ;
        RECT 101.380 80.765 102.310 81.675 ;
        RECT 106.990 80.775 107.920 81.685 ;
        RECT 97.010 80.735 97.115 80.755 ;
        RECT 101.380 80.745 101.485 80.765 ;
        RECT 106.990 80.755 107.095 80.775 ;
        RECT 96.945 80.565 97.115 80.735 ;
        RECT 101.315 80.575 101.485 80.745 ;
        RECT 106.925 80.585 107.095 80.755 ;
        RECT 110.830 80.725 111.760 81.635 ;
        RECT 115.200 80.735 116.130 81.645 ;
        RECT 110.830 80.705 110.935 80.725 ;
        RECT 115.200 80.715 115.305 80.735 ;
        RECT 110.765 80.535 110.935 80.705 ;
        RECT 115.135 80.545 115.305 80.715 ;
        RECT 47.295 80.045 47.465 80.235 ;
      LAYER nwell ;
        RECT 22.640 77.795 25.320 79.400 ;
      LAYER pwell ;
        RECT 23.975 77.415 24.925 77.505 ;
        RECT 22.995 76.595 24.925 77.415 ;
      LAYER nwell ;
        RECT 32.850 77.245 36.450 78.850 ;
        RECT 47.450 77.715 50.130 79.320 ;
      LAYER pwell ;
        RECT 48.785 77.335 49.735 77.425 ;
        RECT 35.120 76.725 36.255 76.955 ;
        RECT 22.995 76.575 23.145 76.595 ;
        RECT 22.975 76.405 23.145 76.575 ;
      LAYER nwell ;
        RECT 22.200 73.695 25.800 75.300 ;
        RECT 28.560 74.745 31.240 76.350 ;
      LAYER pwell ;
        RECT 33.045 76.045 36.255 76.725 ;
        RECT 47.805 76.515 49.735 77.335 ;
      LAYER nwell ;
        RECT 57.660 77.165 61.260 78.770 ;
      LAYER pwell ;
        RECT 59.930 76.645 61.065 76.875 ;
        RECT 47.805 76.495 47.955 76.515 ;
        RECT 47.785 76.325 47.955 76.495 ;
        RECT 33.185 75.855 33.355 76.045 ;
        RECT 29.895 74.365 30.845 74.455 ;
        RECT 28.915 73.545 30.845 74.365 ;
      LAYER nwell ;
        RECT 47.010 73.615 50.610 75.220 ;
        RECT 53.370 74.665 56.050 76.270 ;
      LAYER pwell ;
        RECT 57.855 75.965 61.065 76.645 ;
        RECT 57.995 75.775 58.165 75.965 ;
        RECT 54.705 74.285 55.655 74.375 ;
        RECT 28.915 73.525 29.065 73.545 ;
        RECT 22.435 72.495 25.605 73.405 ;
        RECT 28.895 73.355 29.065 73.525 ;
        RECT 53.725 73.465 55.655 74.285 ;
        RECT 53.725 73.445 53.875 73.465 ;
        RECT 22.535 72.305 22.705 72.495 ;
        RECT 47.245 72.415 50.415 73.325 ;
        RECT 53.705 73.275 53.875 73.445 ;
      LAYER nwell ;
        RECT 117.230 72.745 127.270 74.350 ;
      LAYER pwell ;
        RECT 120.630 72.440 121.980 72.475 ;
        RECT 47.345 72.225 47.515 72.415 ;
        RECT 119.690 72.395 121.980 72.440 ;
        RECT 118.750 72.225 121.980 72.395 ;
        RECT 125.055 72.455 125.975 72.475 ;
        RECT 125.055 72.225 127.075 72.455 ;
        RECT 117.425 71.795 127.075 72.225 ;
        RECT 117.425 71.760 120.620 71.795 ;
        RECT 117.425 71.715 119.680 71.760 ;
      LAYER nwell ;
        RECT 22.690 69.975 25.370 71.580 ;
      LAYER pwell ;
        RECT 117.425 71.545 119.185 71.715 ;
        RECT 121.980 71.545 127.075 71.795 ;
      LAYER nwell ;
        RECT 28.930 69.915 32.530 71.520 ;
        RECT 38.020 69.835 41.160 71.440 ;
        RECT 47.500 69.895 50.180 71.500 ;
        RECT 53.740 69.835 57.340 71.440 ;
        RECT 62.830 69.755 65.970 71.360 ;
      LAYER pwell ;
        RECT 117.565 71.355 117.735 71.545 ;
        RECT 24.025 69.595 24.975 69.685 ;
        RECT 23.045 68.775 24.975 69.595 ;
        RECT 31.200 69.395 32.335 69.625 ;
        RECT 23.045 68.755 23.195 68.775 ;
        RECT 23.025 68.585 23.195 68.755 ;
        RECT 29.125 68.715 32.335 69.395 ;
        RECT 29.265 68.525 29.435 68.715 ;
      LAYER nwell ;
        RECT 33.780 68.045 36.460 69.650 ;
      LAYER pwell ;
        RECT 40.020 69.345 40.965 69.545 ;
        RECT 48.835 69.515 49.785 69.605 ;
        RECT 38.215 68.665 40.965 69.345 ;
        RECT 47.855 68.695 49.785 69.515 ;
        RECT 56.010 69.315 57.145 69.545 ;
        RECT 47.855 68.675 48.005 68.695 ;
        RECT 38.360 68.445 38.530 68.665 ;
        RECT 40.020 68.635 40.965 68.665 ;
        RECT 47.835 68.505 48.005 68.675 ;
        RECT 53.935 68.635 57.145 69.315 ;
        RECT 54.075 68.445 54.245 68.635 ;
      LAYER nwell ;
        RECT 58.590 67.965 61.270 69.570 ;
      LAYER pwell ;
        RECT 64.830 69.265 65.775 69.465 ;
        RECT 63.025 68.585 65.775 69.265 ;
        RECT 63.170 68.365 63.340 68.585 ;
        RECT 64.830 68.555 65.775 68.585 ;
        RECT 35.025 67.525 35.955 67.755 ;
      LAYER nwell ;
        RECT 22.160 65.355 25.760 66.960 ;
        RECT 29.550 65.705 32.230 67.310 ;
      LAYER pwell ;
        RECT 34.120 66.845 35.955 67.525 ;
        RECT 59.835 67.445 60.765 67.675 ;
        RECT 34.120 66.825 34.285 66.845 ;
        RECT 34.115 66.655 34.285 66.825 ;
        RECT 31.115 65.185 32.035 65.415 ;
      LAYER nwell ;
        RECT 46.970 65.275 50.570 66.880 ;
        RECT 54.360 65.625 57.040 67.230 ;
      LAYER pwell ;
        RECT 58.930 66.765 60.765 67.445 ;
        RECT 58.930 66.745 59.095 66.765 ;
        RECT 58.925 66.575 59.095 66.745 ;
        RECT 22.395 64.155 25.565 65.065 ;
        RECT 29.745 64.505 32.035 65.185 ;
        RECT 55.925 65.105 56.845 65.335 ;
        RECT 29.885 64.315 30.055 64.505 ;
        RECT 22.495 63.965 22.665 64.155 ;
        RECT 47.205 64.075 50.375 64.985 ;
        RECT 54.555 64.425 56.845 65.105 ;
        RECT 54.695 64.235 54.865 64.425 ;
        RECT 47.305 63.885 47.475 64.075 ;
      LAYER nwell ;
        RECT 22.650 61.635 25.330 63.240 ;
      LAYER pwell ;
        RECT 23.985 61.255 24.935 61.345 ;
        RECT 23.005 60.435 24.935 61.255 ;
      LAYER nwell ;
        RECT 29.530 60.605 32.210 62.210 ;
        RECT 47.460 61.555 50.140 63.160 ;
      LAYER pwell ;
        RECT 48.795 61.175 49.745 61.265 ;
        RECT 23.005 60.415 23.155 60.435 ;
        RECT 22.985 60.245 23.155 60.415 ;
        RECT 47.815 60.355 49.745 61.175 ;
      LAYER nwell ;
        RECT 54.340 60.525 57.020 62.130 ;
      LAYER pwell ;
        RECT 47.815 60.335 47.965 60.355 ;
        RECT 30.865 60.225 31.815 60.315 ;
        RECT 29.885 59.405 31.815 60.225 ;
        RECT 47.795 60.165 47.965 60.335 ;
        RECT 55.675 60.145 56.625 60.235 ;
        RECT 29.885 59.385 30.035 59.405 ;
        RECT 29.865 59.215 30.035 59.385 ;
        RECT 54.695 59.325 56.625 60.145 ;
        RECT 54.695 59.305 54.845 59.325 ;
      LAYER nwell ;
        RECT 22.210 57.535 25.810 59.140 ;
      LAYER pwell ;
        RECT 54.675 59.135 54.845 59.305 ;
      LAYER nwell ;
        RECT 47.020 57.455 50.620 59.060 ;
      LAYER pwell ;
        RECT 22.445 56.335 25.615 57.245 ;
        RECT 22.545 56.145 22.715 56.335 ;
        RECT 47.255 56.255 50.425 57.165 ;
        RECT 47.355 56.065 47.525 56.255 ;
      LAYER nwell ;
        RECT 22.700 53.815 25.380 55.420 ;
        RECT 47.510 53.735 50.190 55.340 ;
      LAYER pwell ;
        RECT 24.035 53.435 24.985 53.525 ;
        RECT 23.055 52.615 24.985 53.435 ;
        RECT 48.845 53.355 49.795 53.445 ;
        RECT 23.055 52.595 23.205 52.615 ;
        RECT 23.035 52.425 23.205 52.595 ;
        RECT 47.865 52.535 49.795 53.355 ;
        RECT 47.865 52.515 48.015 52.535 ;
        RECT 47.845 52.345 48.015 52.515 ;
        RECT 31.625 32.915 31.795 33.085 ;
        RECT 31.625 32.895 31.730 32.915 ;
        RECT 30.800 31.985 31.730 32.895 ;
      LAYER nwell ;
        RECT 30.370 30.090 32.130 31.695 ;
      LAYER pwell ;
        RECT 53.130 29.735 53.300 29.925 ;
        RECT 46.270 29.055 53.445 29.735 ;
        RECT 62.480 29.715 62.650 29.905 ;
        RECT 46.270 28.825 47.200 29.055 ;
        RECT 52.515 28.825 53.445 29.055 ;
        RECT 55.620 29.035 62.795 29.715 ;
        RECT 71.560 29.695 71.730 29.885 ;
        RECT 55.620 28.805 56.550 29.035 ;
        RECT 61.865 28.805 62.795 29.035 ;
        RECT 64.700 29.015 71.875 29.695 ;
        RECT 80.910 29.675 81.080 29.865 ;
        RECT 64.700 28.785 65.630 29.015 ;
        RECT 70.945 28.785 71.875 29.015 ;
        RECT 74.050 28.995 81.225 29.675 ;
        RECT 74.050 28.765 74.980 28.995 ;
        RECT 80.295 28.765 81.225 28.995 ;
        RECT 16.220 27.635 16.390 27.825 ;
        RECT 9.360 26.955 16.535 27.635 ;
        RECT 25.570 27.615 25.740 27.805 ;
        RECT 9.360 26.725 10.290 26.955 ;
        RECT 15.605 26.725 16.535 26.955 ;
        RECT 18.710 26.935 25.885 27.615 ;
        RECT 34.650 27.595 34.820 27.785 ;
        RECT 18.710 26.705 19.640 26.935 ;
        RECT 24.955 26.705 25.885 26.935 ;
        RECT 27.790 26.915 34.965 27.595 ;
        RECT 44.000 27.575 44.170 27.765 ;
        RECT 27.790 26.685 28.720 26.915 ;
        RECT 34.035 26.685 34.965 26.915 ;
        RECT 37.140 26.895 44.315 27.575 ;
      LAYER nwell ;
        RECT 45.900 26.930 53.640 28.535 ;
        RECT 55.250 26.910 62.990 28.515 ;
      LAYER pwell ;
        RECT 37.140 26.665 38.070 26.895 ;
        RECT 43.385 26.665 44.315 26.895 ;
      LAYER nwell ;
        RECT 64.330 26.890 72.070 28.495 ;
        RECT 73.680 26.870 81.420 28.475 ;
      LAYER pwell ;
        RECT 87.560 26.875 87.730 27.065 ;
      LAYER nwell ;
        RECT 8.990 24.830 16.730 26.435 ;
        RECT 18.340 24.810 26.080 26.415 ;
        RECT 27.420 24.790 35.160 26.395 ;
        RECT 36.770 24.770 44.510 26.375 ;
      LAYER pwell ;
        RECT 84.245 26.195 88.145 26.875 ;
        RECT 87.215 25.965 88.145 26.195 ;
        RECT 53.270 25.365 53.440 25.555 ;
        RECT 46.410 24.685 53.585 25.365 ;
        RECT 62.620 25.345 62.790 25.535 ;
        RECT 46.410 24.455 47.340 24.685 ;
        RECT 52.655 24.455 53.585 24.685 ;
        RECT 55.760 24.665 62.935 25.345 ;
        RECT 71.700 25.325 71.870 25.515 ;
        RECT 55.760 24.435 56.690 24.665 ;
        RECT 62.005 24.435 62.935 24.665 ;
        RECT 64.840 24.645 72.015 25.325 ;
        RECT 81.050 25.305 81.220 25.495 ;
        RECT 64.840 24.415 65.770 24.645 ;
        RECT 71.085 24.415 72.015 24.645 ;
        RECT 74.190 24.625 81.365 25.305 ;
        RECT 74.190 24.395 75.120 24.625 ;
        RECT 80.435 24.395 81.365 24.625 ;
      LAYER nwell ;
        RECT 46.040 22.560 53.780 24.165 ;
        RECT 55.390 22.540 63.130 24.145 ;
        RECT 64.470 22.520 72.210 24.125 ;
        RECT 73.820 22.500 81.560 24.105 ;
        RECT 83.820 24.070 88.340 25.675 ;
      LAYER pwell ;
        RECT 31.475 16.615 31.645 16.785 ;
        RECT 31.475 16.595 31.580 16.615 ;
        RECT 30.650 15.685 31.580 16.595 ;
      LAYER nwell ;
        RECT 30.220 13.790 31.980 15.395 ;
      LAYER pwell ;
        RECT 16.070 11.335 16.240 11.525 ;
        RECT 9.210 10.655 16.385 11.335 ;
        RECT 25.420 11.315 25.590 11.505 ;
        RECT 9.210 10.425 10.140 10.655 ;
        RECT 15.455 10.425 16.385 10.655 ;
        RECT 18.560 10.635 25.735 11.315 ;
        RECT 34.500 11.295 34.670 11.485 ;
        RECT 18.560 10.405 19.490 10.635 ;
        RECT 24.805 10.405 25.735 10.635 ;
        RECT 27.640 10.615 34.815 11.295 ;
        RECT 43.850 11.275 44.020 11.465 ;
        RECT 27.640 10.385 28.570 10.615 ;
        RECT 33.885 10.385 34.815 10.615 ;
        RECT 36.990 10.595 44.165 11.275 ;
        RECT 52.920 11.265 53.090 11.455 ;
        RECT 36.990 10.365 37.920 10.595 ;
        RECT 43.235 10.365 44.165 10.595 ;
        RECT 46.060 10.585 53.235 11.265 ;
        RECT 62.270 11.245 62.440 11.435 ;
        RECT 46.060 10.355 46.990 10.585 ;
        RECT 52.305 10.355 53.235 10.585 ;
        RECT 55.410 10.565 62.585 11.245 ;
        RECT 71.350 11.225 71.520 11.415 ;
        RECT 55.410 10.335 56.340 10.565 ;
        RECT 61.655 10.335 62.585 10.565 ;
        RECT 64.490 10.545 71.665 11.225 ;
        RECT 80.700 11.205 80.870 11.395 ;
        RECT 64.490 10.315 65.420 10.545 ;
        RECT 70.735 10.315 71.665 10.545 ;
        RECT 73.840 10.525 81.015 11.205 ;
        RECT 73.840 10.295 74.770 10.525 ;
        RECT 80.085 10.295 81.015 10.525 ;
      LAYER nwell ;
        RECT 8.840 8.530 16.580 10.135 ;
        RECT 18.190 8.510 25.930 10.115 ;
        RECT 27.270 8.490 35.010 10.095 ;
        RECT 36.620 8.470 44.360 10.075 ;
        RECT 45.690 8.460 53.430 10.065 ;
        RECT 55.040 8.440 62.780 10.045 ;
        RECT 64.120 8.420 71.860 10.025 ;
        RECT 73.470 8.400 81.210 10.005 ;
      LAYER li1 ;
        RECT 47.150 88.885 48.530 89.055 ;
        RECT 47.480 88.085 47.810 88.715 ;
        RECT 47.480 87.485 47.710 88.085 ;
        RECT 47.980 88.065 48.210 88.885 ;
        RECT 47.880 87.655 48.210 87.895 ;
        RECT 47.480 86.505 47.810 87.485 ;
        RECT 47.980 86.335 48.190 87.475 ;
        RECT 47.150 86.165 48.530 86.335 ;
        RECT 81.680 83.385 83.060 83.555 ;
        RECT 22.340 82.845 25.560 83.015 ;
        RECT 22.425 81.995 22.805 82.675 ;
        RECT 23.395 81.995 23.565 82.845 ;
        RECT 23.735 82.165 24.065 82.675 ;
        RECT 24.235 82.335 24.405 82.845 ;
        RECT 47.150 82.765 50.370 82.935 ;
        RECT 24.575 82.165 24.975 82.675 ;
        RECT 23.735 81.995 24.975 82.165 ;
        RECT 22.425 81.035 22.595 81.995 ;
        RECT 22.765 81.655 24.070 81.825 ;
        RECT 25.155 81.745 25.475 82.675 ;
        RECT 22.765 81.205 23.010 81.655 ;
        RECT 23.180 81.285 23.730 81.485 ;
        RECT 23.900 81.455 24.070 81.655 ;
        RECT 24.845 81.575 25.475 81.745 ;
        RECT 47.235 81.915 47.615 82.595 ;
        RECT 48.205 81.915 48.375 82.765 ;
        RECT 48.545 82.085 48.875 82.595 ;
        RECT 49.045 82.255 49.215 82.765 ;
        RECT 49.385 82.085 49.785 82.595 ;
        RECT 48.545 81.915 49.785 82.085 ;
        RECT 23.900 81.285 24.275 81.455 ;
        RECT 24.445 81.035 24.675 81.535 ;
        RECT 22.425 80.865 24.675 81.035 ;
        RECT 22.475 80.295 22.805 80.685 ;
        RECT 22.975 80.545 23.145 80.865 ;
        RECT 24.845 80.695 25.015 81.575 ;
        RECT 23.315 80.295 23.645 80.685 ;
        RECT 24.060 80.525 25.015 80.695 ;
        RECT 25.185 80.295 25.475 81.130 ;
        RECT 47.235 80.955 47.405 81.915 ;
        RECT 47.575 81.575 48.880 81.745 ;
        RECT 49.965 81.665 50.285 82.595 ;
        RECT 82.020 82.245 82.230 83.385 ;
        RECT 85.520 83.335 86.900 83.505 ;
        RECT 89.890 83.345 91.270 83.515 ;
        RECT 82.400 82.235 82.730 83.215 ;
        RECT 82.000 81.825 82.330 82.065 ;
        RECT 47.575 81.125 47.820 81.575 ;
        RECT 47.990 81.205 48.540 81.405 ;
        RECT 48.710 81.375 48.880 81.575 ;
        RECT 49.655 81.495 50.285 81.665 ;
        RECT 48.710 81.205 49.085 81.375 ;
        RECT 49.255 80.955 49.485 81.455 ;
        RECT 47.235 80.785 49.485 80.955 ;
        RECT 22.340 80.125 25.560 80.295 ;
        RECT 47.285 80.215 47.615 80.605 ;
        RECT 47.785 80.465 47.955 80.785 ;
        RECT 49.655 80.615 49.825 81.495 ;
        RECT 48.125 80.215 48.455 80.605 ;
        RECT 48.870 80.445 49.825 80.615 ;
        RECT 49.995 80.215 50.285 81.050 ;
        RECT 82.000 80.835 82.230 81.655 ;
        RECT 82.500 81.635 82.730 82.235 ;
        RECT 85.860 82.195 86.070 83.335 ;
        RECT 86.240 82.185 86.570 83.165 ;
        RECT 90.230 82.205 90.440 83.345 ;
        RECT 92.960 83.335 94.340 83.505 ;
        RECT 90.610 82.195 90.940 83.175 ;
        RECT 93.300 82.195 93.510 83.335 ;
        RECT 96.800 83.285 98.180 83.455 ;
        RECT 101.170 83.295 102.550 83.465 ;
        RECT 106.780 83.305 108.160 83.475 ;
        RECT 85.840 81.775 86.170 82.015 ;
        RECT 82.400 81.005 82.730 81.635 ;
        RECT 81.680 80.665 83.060 80.835 ;
        RECT 85.840 80.785 86.070 81.605 ;
        RECT 86.340 81.585 86.570 82.185 ;
        RECT 90.210 81.785 90.540 82.025 ;
        RECT 86.240 80.955 86.570 81.585 ;
        RECT 90.210 80.795 90.440 81.615 ;
        RECT 90.710 81.595 90.940 82.195 ;
        RECT 93.680 82.185 94.010 83.165 ;
        RECT 93.280 81.775 93.610 82.015 ;
        RECT 90.610 80.965 90.940 81.595 ;
        RECT 85.520 80.615 86.900 80.785 ;
        RECT 89.890 80.625 91.270 80.795 ;
        RECT 93.280 80.785 93.510 81.605 ;
        RECT 93.780 81.585 94.010 82.185 ;
        RECT 97.140 82.145 97.350 83.285 ;
        RECT 97.520 82.135 97.850 83.115 ;
        RECT 101.510 82.155 101.720 83.295 ;
        RECT 101.890 82.145 102.220 83.125 ;
        RECT 107.120 82.165 107.330 83.305 ;
        RECT 110.620 83.255 112.000 83.425 ;
        RECT 114.990 83.265 116.370 83.435 ;
        RECT 107.500 82.155 107.830 83.135 ;
        RECT 97.120 81.725 97.450 81.965 ;
        RECT 93.680 80.955 94.010 81.585 ;
        RECT 92.960 80.615 94.340 80.785 ;
        RECT 97.120 80.735 97.350 81.555 ;
        RECT 97.620 81.535 97.850 82.135 ;
        RECT 101.490 81.735 101.820 81.975 ;
        RECT 97.520 80.905 97.850 81.535 ;
        RECT 101.490 80.745 101.720 81.565 ;
        RECT 101.990 81.545 102.220 82.145 ;
        RECT 107.100 81.745 107.430 81.985 ;
        RECT 101.890 80.915 102.220 81.545 ;
        RECT 107.100 80.755 107.330 81.575 ;
        RECT 107.600 81.555 107.830 82.155 ;
        RECT 110.960 82.115 111.170 83.255 ;
        RECT 111.340 82.105 111.670 83.085 ;
        RECT 115.330 82.125 115.540 83.265 ;
        RECT 115.710 82.115 116.040 83.095 ;
        RECT 110.940 81.695 111.270 81.935 ;
        RECT 107.500 80.925 107.830 81.555 ;
        RECT 96.800 80.565 98.180 80.735 ;
        RECT 101.170 80.575 102.550 80.745 ;
        RECT 106.780 80.585 108.160 80.755 ;
        RECT 110.940 80.705 111.170 81.525 ;
        RECT 111.440 81.505 111.670 82.105 ;
        RECT 115.310 81.705 115.640 81.945 ;
        RECT 111.340 80.875 111.670 81.505 ;
        RECT 115.310 80.715 115.540 81.535 ;
        RECT 115.810 81.515 116.040 82.115 ;
        RECT 115.710 80.885 116.040 81.515 ;
        RECT 110.620 80.535 112.000 80.705 ;
        RECT 114.990 80.545 116.370 80.715 ;
        RECT 47.150 80.045 50.370 80.215 ;
        RECT 22.830 79.125 25.130 79.295 ;
        RECT 23.115 78.455 23.395 79.125 ;
        RECT 23.565 78.235 23.865 78.785 ;
        RECT 24.065 78.405 24.395 79.125 ;
        RECT 47.640 79.045 49.940 79.215 ;
        RECT 24.585 78.405 25.045 78.955 ;
        RECT 33.040 78.575 36.260 78.745 ;
        RECT 22.930 77.815 23.195 78.175 ;
        RECT 23.565 78.065 24.505 78.235 ;
        RECT 24.335 77.815 24.505 78.065 ;
        RECT 22.930 77.565 23.605 77.815 ;
        RECT 23.825 77.565 24.165 77.815 ;
        RECT 24.335 77.485 24.625 77.815 ;
        RECT 24.335 77.395 24.505 77.485 ;
        RECT 23.115 77.205 24.505 77.395 ;
        RECT 23.115 76.845 23.445 77.205 ;
        RECT 24.795 77.035 25.045 78.405 ;
        RECT 33.130 78.195 33.465 78.575 ;
        RECT 24.065 76.575 24.315 77.035 ;
        RECT 24.485 76.745 25.045 77.035 ;
        RECT 33.125 76.705 33.365 78.015 ;
        RECT 33.635 77.605 33.885 78.405 ;
        RECT 34.105 77.855 34.435 78.575 ;
        RECT 34.620 77.605 34.870 78.405 ;
        RECT 35.335 77.775 35.665 78.575 ;
        RECT 35.835 78.145 36.175 78.405 ;
        RECT 47.925 78.375 48.205 79.045 ;
        RECT 33.535 77.435 35.725 77.605 ;
        RECT 22.830 76.405 25.130 76.575 ;
        RECT 33.535 76.525 33.705 77.435 ;
        RECT 35.410 77.265 35.725 77.435 ;
        RECT 28.750 76.075 31.050 76.245 ;
        RECT 33.210 76.195 33.705 76.525 ;
        RECT 33.925 76.300 34.275 77.265 ;
        RECT 34.455 76.295 34.755 77.265 ;
        RECT 34.935 76.295 35.215 77.265 ;
        RECT 35.410 77.015 35.740 77.265 ;
        RECT 29.035 75.405 29.315 76.075 ;
        RECT 22.390 75.025 25.610 75.195 ;
        RECT 29.485 75.185 29.785 75.735 ;
        RECT 29.985 75.355 30.315 76.075 ;
        RECT 35.395 76.025 35.665 76.825 ;
        RECT 35.915 76.745 36.175 78.145 ;
        RECT 48.375 78.155 48.675 78.705 ;
        RECT 48.875 78.325 49.205 79.045 ;
        RECT 49.395 78.325 49.855 78.875 ;
        RECT 57.850 78.495 61.070 78.665 ;
        RECT 47.740 77.735 48.005 78.095 ;
        RECT 48.375 77.985 49.315 78.155 ;
        RECT 49.145 77.735 49.315 77.985 ;
        RECT 47.740 77.485 48.415 77.735 ;
        RECT 48.635 77.485 48.975 77.735 ;
        RECT 49.145 77.405 49.435 77.735 ;
        RECT 49.145 77.315 49.315 77.405 ;
        RECT 47.925 77.125 49.315 77.315 ;
        RECT 47.925 76.765 48.255 77.125 ;
        RECT 49.605 76.955 49.855 78.325 ;
        RECT 57.940 78.115 58.275 78.495 ;
        RECT 35.835 76.235 36.175 76.745 ;
        RECT 48.875 76.495 49.125 76.955 ;
        RECT 49.295 76.665 49.855 76.955 ;
        RECT 57.935 76.625 58.175 77.935 ;
        RECT 58.445 77.525 58.695 78.325 ;
        RECT 58.915 77.775 59.245 78.495 ;
        RECT 59.430 77.525 59.680 78.325 ;
        RECT 60.145 77.695 60.475 78.495 ;
        RECT 60.645 78.065 60.985 78.325 ;
        RECT 58.345 77.355 60.535 77.525 ;
        RECT 47.640 76.325 49.940 76.495 ;
        RECT 58.345 76.445 58.515 77.355 ;
        RECT 60.220 77.185 60.535 77.355 ;
        RECT 30.505 75.355 30.965 75.905 ;
        RECT 33.040 75.855 36.260 76.025 ;
        RECT 53.560 75.995 55.860 76.165 ;
        RECT 58.020 76.115 58.515 76.445 ;
        RECT 58.735 76.220 59.085 77.185 ;
        RECT 59.265 76.215 59.565 77.185 ;
        RECT 59.745 76.215 60.025 77.185 ;
        RECT 60.220 76.935 60.550 77.185 ;
        RECT 22.475 74.175 22.855 74.855 ;
        RECT 23.445 74.175 23.615 75.025 ;
        RECT 23.785 74.345 24.115 74.855 ;
        RECT 24.285 74.515 24.455 75.025 ;
        RECT 24.625 74.345 25.025 74.855 ;
        RECT 23.785 74.175 25.025 74.345 ;
        RECT 22.475 73.215 22.645 74.175 ;
        RECT 22.815 73.835 24.120 74.005 ;
        RECT 25.205 73.925 25.525 74.855 ;
        RECT 28.850 74.765 29.115 75.125 ;
        RECT 29.485 75.015 30.425 75.185 ;
        RECT 30.255 74.765 30.425 75.015 ;
        RECT 28.850 74.515 29.525 74.765 ;
        RECT 29.745 74.515 30.085 74.765 ;
        RECT 30.255 74.435 30.545 74.765 ;
        RECT 30.255 74.345 30.425 74.435 ;
        RECT 22.815 73.385 23.060 73.835 ;
        RECT 23.230 73.465 23.780 73.665 ;
        RECT 23.950 73.635 24.120 73.835 ;
        RECT 24.895 73.755 25.525 73.925 ;
        RECT 29.035 74.155 30.425 74.345 ;
        RECT 29.035 73.795 29.365 74.155 ;
        RECT 30.715 73.985 30.965 75.355 ;
        RECT 53.845 75.325 54.125 75.995 ;
        RECT 47.200 74.945 50.420 75.115 ;
        RECT 54.295 75.105 54.595 75.655 ;
        RECT 54.795 75.275 55.125 75.995 ;
        RECT 60.205 75.945 60.475 76.745 ;
        RECT 60.725 76.665 60.985 78.065 ;
        RECT 60.645 76.155 60.985 76.665 ;
        RECT 55.315 75.275 55.775 75.825 ;
        RECT 57.850 75.775 61.070 75.945 ;
        RECT 23.950 73.465 24.325 73.635 ;
        RECT 24.495 73.215 24.725 73.715 ;
        RECT 22.475 73.045 24.725 73.215 ;
        RECT 22.525 72.475 22.855 72.865 ;
        RECT 23.025 72.725 23.195 73.045 ;
        RECT 24.895 72.875 25.065 73.755 ;
        RECT 29.985 73.525 30.235 73.985 ;
        RECT 30.405 73.695 30.965 73.985 ;
        RECT 47.285 74.095 47.665 74.775 ;
        RECT 48.255 74.095 48.425 74.945 ;
        RECT 48.595 74.265 48.925 74.775 ;
        RECT 49.095 74.435 49.265 74.945 ;
        RECT 49.435 74.265 49.835 74.775 ;
        RECT 48.595 74.095 49.835 74.265 ;
        RECT 28.750 73.355 31.050 73.525 ;
        RECT 23.365 72.475 23.695 72.865 ;
        RECT 24.110 72.705 25.065 72.875 ;
        RECT 25.235 72.475 25.525 73.310 ;
        RECT 47.285 73.135 47.455 74.095 ;
        RECT 47.625 73.755 48.930 73.925 ;
        RECT 50.015 73.845 50.335 74.775 ;
        RECT 53.660 74.685 53.925 75.045 ;
        RECT 54.295 74.935 55.235 75.105 ;
        RECT 55.065 74.685 55.235 74.935 ;
        RECT 53.660 74.435 54.335 74.685 ;
        RECT 54.555 74.435 54.895 74.685 ;
        RECT 55.065 74.355 55.355 74.685 ;
        RECT 55.065 74.265 55.235 74.355 ;
        RECT 47.625 73.305 47.870 73.755 ;
        RECT 48.040 73.385 48.590 73.585 ;
        RECT 48.760 73.555 48.930 73.755 ;
        RECT 49.705 73.675 50.335 73.845 ;
        RECT 53.845 74.075 55.235 74.265 ;
        RECT 53.845 73.715 54.175 74.075 ;
        RECT 55.525 73.905 55.775 75.275 ;
        RECT 117.420 74.075 127.080 74.245 ;
        RECT 48.760 73.385 49.135 73.555 ;
        RECT 49.305 73.135 49.535 73.635 ;
        RECT 47.285 72.965 49.535 73.135 ;
        RECT 22.390 72.305 25.610 72.475 ;
        RECT 47.335 72.395 47.665 72.785 ;
        RECT 47.835 72.645 48.005 72.965 ;
        RECT 49.705 72.795 49.875 73.675 ;
        RECT 54.795 73.445 55.045 73.905 ;
        RECT 55.215 73.615 55.775 73.905 ;
        RECT 53.560 73.275 55.860 73.445 ;
        RECT 117.595 73.405 117.765 73.905 ;
        RECT 117.935 73.695 118.265 74.075 ;
        RECT 118.435 73.735 119.965 73.905 ;
        RECT 118.435 73.575 118.605 73.735 ;
        RECT 118.955 73.405 119.125 73.565 ;
        RECT 117.595 73.235 119.125 73.405 ;
        RECT 119.295 73.395 119.625 73.565 ;
        RECT 48.175 72.395 48.505 72.785 ;
        RECT 48.920 72.625 49.875 72.795 ;
        RECT 50.045 72.395 50.335 73.230 ;
        RECT 119.295 73.065 119.465 73.395 ;
        RECT 119.795 73.235 119.965 73.735 ;
        RECT 120.135 73.065 120.485 73.905 ;
        RECT 120.655 73.695 120.985 74.075 ;
        RECT 121.245 73.735 122.255 73.905 ;
        RECT 117.570 72.435 117.915 73.055 ;
        RECT 118.225 72.435 118.660 73.055 ;
        RECT 118.830 72.895 119.465 73.065 ;
        RECT 47.200 72.225 50.420 72.395 ;
        RECT 118.830 72.375 119.000 72.895 ;
        RECT 119.680 72.835 120.485 73.065 ;
        RECT 119.680 72.725 120.040 72.835 ;
        RECT 119.500 72.545 120.040 72.725 ;
        RECT 117.595 72.075 118.605 72.245 ;
        RECT 117.595 71.700 117.765 72.075 ;
        RECT 117.935 71.525 118.265 71.905 ;
        RECT 118.435 71.865 118.605 72.075 ;
        RECT 118.830 72.205 119.120 72.375 ;
        RECT 118.830 72.035 119.170 72.205 ;
        RECT 119.340 71.865 119.510 72.200 ;
        RECT 119.680 71.870 120.040 72.545 ;
        RECT 120.685 72.435 120.985 73.435 ;
        RECT 121.245 73.225 121.415 73.735 ;
        RECT 121.585 73.055 121.915 73.565 ;
        RECT 122.085 73.525 122.255 73.735 ;
        RECT 122.480 73.695 122.810 74.075 ;
        RECT 122.980 73.525 123.150 73.905 ;
        RECT 123.400 73.695 123.750 74.075 ;
        RECT 123.920 73.575 124.105 73.905 ;
        RECT 122.085 73.355 123.150 73.525 ;
        RECT 121.155 72.885 121.915 73.055 ;
        RECT 121.155 72.360 121.325 72.885 ;
        RECT 121.710 72.705 121.880 72.715 ;
        RECT 121.495 72.545 121.880 72.705 ;
        RECT 121.495 72.535 121.825 72.545 ;
        RECT 122.220 72.495 122.465 73.115 ;
        RECT 122.670 72.495 123.000 73.115 ;
        RECT 123.475 72.435 123.765 73.115 ;
        RECT 123.935 72.715 124.105 73.575 ;
        RECT 124.400 73.575 124.610 73.905 ;
        RECT 124.780 73.735 126.065 73.905 ;
        RECT 124.780 73.695 125.110 73.735 ;
        RECT 123.935 72.545 124.225 72.715 ;
        RECT 121.155 72.285 121.470 72.360 ;
        RECT 118.435 71.695 119.510 71.865 ;
        RECT 120.220 71.525 120.510 72.245 ;
        RECT 120.800 71.865 120.970 72.235 ;
        RECT 121.140 72.035 121.470 72.285 ;
        RECT 121.640 72.325 121.810 72.365 ;
        RECT 121.640 72.155 123.160 72.325 ;
        RECT 121.640 72.035 121.810 72.155 ;
        RECT 122.045 71.865 122.400 71.905 ;
        RECT 120.800 71.695 122.400 71.865 ;
        RECT 122.570 71.525 122.740 71.985 ;
        RECT 122.915 71.735 123.160 72.155 ;
        RECT 123.935 72.095 124.105 72.545 ;
        RECT 124.400 72.375 124.570 73.575 ;
        RECT 125.265 73.425 125.595 73.565 ;
        RECT 124.810 73.195 125.595 73.425 ;
        RECT 125.895 73.275 126.065 73.735 ;
        RECT 126.235 73.695 126.565 74.075 ;
        RECT 124.400 72.205 124.640 72.375 ;
        RECT 123.430 71.525 123.760 71.905 ;
        RECT 123.930 71.765 124.105 72.095 ;
        RECT 124.810 72.025 124.980 73.195 ;
        RECT 125.895 73.105 126.545 73.275 ;
        RECT 125.610 72.545 126.065 72.715 ;
        RECT 125.390 72.365 125.800 72.375 ;
        RECT 125.390 72.205 125.805 72.365 ;
        RECT 126.375 72.325 126.545 73.105 ;
        RECT 125.630 72.035 125.805 72.205 ;
        RECT 125.975 72.155 126.545 72.325 ;
        RECT 126.735 72.990 126.995 73.905 ;
        RECT 126.735 72.810 127.000 72.990 ;
        RECT 124.450 71.855 124.980 72.025 ;
        RECT 125.150 71.865 125.320 72.025 ;
        RECT 125.975 71.865 126.145 72.155 ;
        RECT 124.450 71.695 124.620 71.855 ;
        RECT 125.150 71.695 126.145 71.865 ;
        RECT 126.315 71.525 126.485 71.985 ;
        RECT 126.735 71.695 126.995 72.810 ;
        RECT 22.880 71.305 25.180 71.475 ;
        RECT 23.165 70.635 23.445 71.305 ;
        RECT 23.615 70.415 23.915 70.965 ;
        RECT 24.115 70.585 24.445 71.305 ;
        RECT 29.120 71.245 32.340 71.415 ;
        RECT 24.635 70.585 25.095 71.135 ;
        RECT 29.210 70.865 29.545 71.245 ;
        RECT 22.980 69.995 23.245 70.355 ;
        RECT 23.615 70.245 24.555 70.415 ;
        RECT 24.385 69.995 24.555 70.245 ;
        RECT 22.980 69.745 23.655 69.995 ;
        RECT 23.875 69.745 24.215 69.995 ;
        RECT 24.385 69.665 24.675 69.995 ;
        RECT 24.385 69.575 24.555 69.665 ;
        RECT 23.165 69.385 24.555 69.575 ;
        RECT 23.165 69.025 23.495 69.385 ;
        RECT 24.845 69.215 25.095 70.585 ;
        RECT 29.205 69.375 29.445 70.685 ;
        RECT 29.715 70.275 29.965 71.075 ;
        RECT 30.185 70.525 30.515 71.245 ;
        RECT 30.700 70.275 30.950 71.075 ;
        RECT 31.415 70.445 31.745 71.245 ;
        RECT 38.210 71.165 40.970 71.335 ;
        RECT 47.690 71.225 49.990 71.395 ;
        RECT 117.420 71.355 127.080 71.525 ;
        RECT 31.915 70.815 32.255 71.075 ;
        RECT 29.615 70.105 31.805 70.275 ;
        RECT 24.115 68.755 24.365 69.215 ;
        RECT 24.535 68.925 25.095 69.215 ;
        RECT 29.615 69.195 29.785 70.105 ;
        RECT 31.490 69.935 31.805 70.105 ;
        RECT 29.290 68.865 29.785 69.195 ;
        RECT 30.005 68.970 30.355 69.935 ;
        RECT 30.535 68.965 30.835 69.935 ;
        RECT 31.015 68.965 31.295 69.935 ;
        RECT 31.490 69.685 31.820 69.935 ;
        RECT 22.880 68.585 25.180 68.755 ;
        RECT 31.475 68.695 31.745 69.495 ;
        RECT 31.995 69.415 32.255 70.815 ;
        RECT 38.300 70.655 39.955 70.945 ;
        RECT 38.300 70.315 39.890 70.485 ;
        RECT 40.125 70.365 40.405 71.165 ;
        RECT 38.300 70.025 38.620 70.315 ;
        RECT 39.720 70.195 39.890 70.315 ;
        RECT 31.915 68.905 32.255 69.415 ;
        RECT 33.970 69.375 36.270 69.545 ;
        RECT 29.120 68.525 32.340 68.695 ;
        RECT 34.240 68.405 34.630 68.580 ;
        RECT 35.115 68.575 35.445 69.375 ;
        RECT 38.300 69.285 38.650 69.855 ;
        RECT 38.820 69.525 39.530 70.145 ;
        RECT 39.720 70.025 40.445 70.195 ;
        RECT 40.615 70.025 40.885 70.995 ;
        RECT 47.975 70.555 48.255 71.225 ;
        RECT 48.425 70.335 48.725 70.885 ;
        RECT 48.925 70.505 49.255 71.225 ;
        RECT 53.930 71.165 57.150 71.335 ;
        RECT 49.445 70.505 49.905 71.055 ;
        RECT 54.020 70.785 54.355 71.165 ;
        RECT 40.275 69.855 40.445 70.025 ;
        RECT 39.700 69.525 40.105 69.855 ;
        RECT 40.275 69.525 40.545 69.855 ;
        RECT 40.275 69.355 40.445 69.525 ;
        RECT 35.615 68.585 36.150 69.205 ;
        RECT 38.835 69.185 40.445 69.355 ;
        RECT 40.715 69.290 40.885 70.025 ;
        RECT 47.790 69.915 48.055 70.275 ;
        RECT 48.425 70.165 49.365 70.335 ;
        RECT 49.195 69.915 49.365 70.165 ;
        RECT 47.790 69.665 48.465 69.915 ;
        RECT 48.685 69.665 49.025 69.915 ;
        RECT 49.195 69.585 49.485 69.915 ;
        RECT 49.195 69.495 49.365 69.585 ;
        RECT 38.305 68.615 38.635 69.115 ;
        RECT 38.835 68.835 39.005 69.185 ;
        RECT 39.205 68.615 39.535 69.015 ;
        RECT 39.705 68.835 39.875 69.185 ;
        RECT 40.045 68.615 40.425 69.015 ;
        RECT 40.615 68.945 40.885 69.290 ;
        RECT 47.975 69.305 49.365 69.495 ;
        RECT 47.975 68.945 48.305 69.305 ;
        RECT 49.655 69.135 49.905 70.505 ;
        RECT 54.015 69.295 54.255 70.605 ;
        RECT 54.525 70.195 54.775 70.995 ;
        RECT 54.995 70.445 55.325 71.165 ;
        RECT 55.510 70.195 55.760 70.995 ;
        RECT 56.225 70.365 56.555 71.165 ;
        RECT 63.020 71.085 65.780 71.255 ;
        RECT 56.725 70.735 57.065 70.995 ;
        RECT 54.425 70.025 56.615 70.195 ;
        RECT 48.925 68.675 49.175 69.135 ;
        RECT 49.345 68.845 49.905 69.135 ;
        RECT 54.425 69.115 54.595 70.025 ;
        RECT 56.300 69.855 56.615 70.025 ;
        RECT 54.100 68.785 54.595 69.115 ;
        RECT 54.815 68.890 55.165 69.855 ;
        RECT 55.345 68.885 55.645 69.855 ;
        RECT 55.825 68.885 56.105 69.855 ;
        RECT 56.300 69.605 56.630 69.855 ;
        RECT 34.240 68.235 35.665 68.405 ;
        RECT 34.115 67.505 34.470 68.065 ;
        RECT 34.640 67.335 34.810 68.235 ;
        RECT 34.980 67.505 35.245 68.065 ;
        RECT 35.495 67.735 35.665 68.235 ;
        RECT 35.835 67.565 36.150 68.585 ;
        RECT 38.210 68.445 40.970 68.615 ;
        RECT 47.690 68.505 49.990 68.675 ;
        RECT 56.285 68.615 56.555 69.415 ;
        RECT 56.805 69.335 57.065 70.735 ;
        RECT 63.110 70.575 64.765 70.865 ;
        RECT 63.110 70.235 64.700 70.405 ;
        RECT 64.935 70.285 65.215 71.085 ;
        RECT 63.110 69.945 63.430 70.235 ;
        RECT 64.530 70.115 64.700 70.235 ;
        RECT 56.725 68.825 57.065 69.335 ;
        RECT 58.780 69.295 61.080 69.465 ;
        RECT 53.930 68.445 57.150 68.615 ;
        RECT 59.050 68.325 59.440 68.500 ;
        RECT 59.925 68.495 60.255 69.295 ;
        RECT 63.110 69.205 63.460 69.775 ;
        RECT 63.630 69.445 64.340 70.065 ;
        RECT 64.530 69.945 65.255 70.115 ;
        RECT 65.425 69.945 65.695 70.915 ;
        RECT 65.085 69.775 65.255 69.945 ;
        RECT 64.510 69.445 64.915 69.775 ;
        RECT 65.085 69.445 65.355 69.775 ;
        RECT 65.085 69.275 65.255 69.445 ;
        RECT 60.425 68.505 60.960 69.125 ;
        RECT 63.645 69.105 65.255 69.275 ;
        RECT 65.525 69.210 65.695 69.945 ;
        RECT 63.115 68.535 63.445 69.035 ;
        RECT 63.645 68.755 63.815 69.105 ;
        RECT 64.015 68.535 64.345 68.935 ;
        RECT 64.515 68.755 64.685 69.105 ;
        RECT 64.855 68.535 65.235 68.935 ;
        RECT 65.425 68.865 65.695 69.210 ;
        RECT 59.050 68.155 60.475 68.325 ;
        RECT 29.740 67.035 32.040 67.205 ;
        RECT 22.350 66.685 25.570 66.855 ;
        RECT 22.435 65.835 22.815 66.515 ;
        RECT 23.405 65.835 23.575 66.685 ;
        RECT 23.745 66.005 24.075 66.515 ;
        RECT 24.245 66.175 24.415 66.685 ;
        RECT 24.585 66.005 24.985 66.515 ;
        RECT 23.745 65.835 24.985 66.005 ;
        RECT 22.435 64.875 22.605 65.835 ;
        RECT 22.775 65.495 24.080 65.665 ;
        RECT 25.165 65.585 25.485 66.515 ;
        RECT 29.825 66.480 30.430 67.035 ;
        RECT 30.605 66.525 31.085 66.865 ;
        RECT 30.730 66.490 30.910 66.525 ;
        RECT 31.255 66.490 31.510 67.035 ;
        RECT 29.825 66.380 30.440 66.480 ;
        RECT 30.255 66.355 30.440 66.380 ;
        RECT 29.825 65.760 30.085 66.210 ;
        RECT 30.255 66.110 30.585 66.355 ;
        RECT 30.755 66.035 31.510 66.285 ;
        RECT 31.680 66.165 31.955 66.865 ;
        RECT 34.220 66.825 34.460 67.335 ;
        RECT 34.640 67.005 34.920 67.335 ;
        RECT 35.150 66.825 35.365 67.335 ;
        RECT 35.535 66.995 36.150 67.565 ;
        RECT 58.925 67.425 59.280 67.985 ;
        RECT 59.450 67.255 59.620 68.155 ;
        RECT 59.790 67.425 60.055 67.985 ;
        RECT 60.305 67.655 60.475 68.155 ;
        RECT 60.645 67.485 60.960 68.505 ;
        RECT 63.020 68.365 65.780 68.535 ;
        RECT 54.550 66.955 56.850 67.125 ;
        RECT 33.970 66.655 36.270 66.825 ;
        RECT 47.160 66.605 50.380 66.775 ;
        RECT 30.740 66.000 31.510 66.035 ;
        RECT 30.725 65.990 31.510 66.000 ;
        RECT 30.720 65.975 31.615 65.990 ;
        RECT 30.700 65.960 31.615 65.975 ;
        RECT 30.680 65.950 31.615 65.960 ;
        RECT 30.655 65.940 31.615 65.950 ;
        RECT 30.585 65.910 31.615 65.940 ;
        RECT 30.565 65.880 31.615 65.910 ;
        RECT 30.545 65.850 31.615 65.880 ;
        RECT 30.515 65.825 31.615 65.850 ;
        RECT 30.480 65.790 31.615 65.825 ;
        RECT 30.450 65.785 31.615 65.790 ;
        RECT 30.450 65.780 30.840 65.785 ;
        RECT 30.450 65.770 30.815 65.780 ;
        RECT 30.450 65.765 30.800 65.770 ;
        RECT 30.450 65.760 30.785 65.765 ;
        RECT 29.825 65.755 30.785 65.760 ;
        RECT 29.825 65.745 30.775 65.755 ;
        RECT 29.825 65.740 30.765 65.745 ;
        RECT 29.825 65.730 30.755 65.740 ;
        RECT 29.825 65.720 30.750 65.730 ;
        RECT 29.825 65.715 30.745 65.720 ;
        RECT 29.825 65.700 30.735 65.715 ;
        RECT 29.825 65.685 30.730 65.700 ;
        RECT 29.825 65.660 30.720 65.685 ;
        RECT 29.825 65.590 30.715 65.660 ;
        RECT 22.775 65.045 23.020 65.495 ;
        RECT 23.190 65.125 23.740 65.325 ;
        RECT 23.910 65.295 24.080 65.495 ;
        RECT 24.855 65.415 25.485 65.585 ;
        RECT 23.910 65.125 24.285 65.295 ;
        RECT 24.455 64.875 24.685 65.375 ;
        RECT 22.435 64.705 24.685 64.875 ;
        RECT 22.485 64.135 22.815 64.525 ;
        RECT 22.985 64.385 23.155 64.705 ;
        RECT 24.855 64.535 25.025 65.415 ;
        RECT 29.825 65.035 30.375 65.420 ;
        RECT 23.325 64.135 23.655 64.525 ;
        RECT 24.070 64.365 25.025 64.535 ;
        RECT 25.195 64.135 25.485 64.970 ;
        RECT 30.545 64.865 30.715 65.590 ;
        RECT 29.825 64.695 30.715 64.865 ;
        RECT 30.885 65.190 31.215 65.615 ;
        RECT 31.385 65.390 31.615 65.785 ;
        RECT 30.885 65.160 31.160 65.190 ;
        RECT 30.885 64.705 31.105 65.160 ;
        RECT 31.785 65.135 31.955 66.165 ;
        RECT 31.275 64.485 31.525 65.025 ;
        RECT 31.695 64.655 31.955 65.135 ;
        RECT 47.245 65.755 47.625 66.435 ;
        RECT 48.215 65.755 48.385 66.605 ;
        RECT 48.555 65.925 48.885 66.435 ;
        RECT 49.055 66.095 49.225 66.605 ;
        RECT 49.395 65.925 49.795 66.435 ;
        RECT 48.555 65.755 49.795 65.925 ;
        RECT 47.245 64.795 47.415 65.755 ;
        RECT 47.585 65.415 48.890 65.585 ;
        RECT 49.975 65.505 50.295 66.435 ;
        RECT 54.635 66.400 55.240 66.955 ;
        RECT 55.415 66.445 55.895 66.785 ;
        RECT 55.540 66.410 55.720 66.445 ;
        RECT 56.065 66.410 56.320 66.955 ;
        RECT 54.635 66.300 55.250 66.400 ;
        RECT 55.065 66.275 55.250 66.300 ;
        RECT 54.635 65.680 54.895 66.130 ;
        RECT 55.065 66.030 55.395 66.275 ;
        RECT 55.565 65.955 56.320 66.205 ;
        RECT 56.490 66.085 56.765 66.785 ;
        RECT 59.030 66.745 59.270 67.255 ;
        RECT 59.450 66.925 59.730 67.255 ;
        RECT 59.960 66.745 60.175 67.255 ;
        RECT 60.345 66.915 60.960 67.485 ;
        RECT 58.780 66.575 61.080 66.745 ;
        RECT 55.550 65.920 56.320 65.955 ;
        RECT 55.535 65.910 56.320 65.920 ;
        RECT 55.530 65.895 56.425 65.910 ;
        RECT 55.510 65.880 56.425 65.895 ;
        RECT 55.490 65.870 56.425 65.880 ;
        RECT 55.465 65.860 56.425 65.870 ;
        RECT 55.395 65.830 56.425 65.860 ;
        RECT 55.375 65.800 56.425 65.830 ;
        RECT 55.355 65.770 56.425 65.800 ;
        RECT 55.325 65.745 56.425 65.770 ;
        RECT 55.290 65.710 56.425 65.745 ;
        RECT 55.260 65.705 56.425 65.710 ;
        RECT 55.260 65.700 55.650 65.705 ;
        RECT 55.260 65.690 55.625 65.700 ;
        RECT 55.260 65.685 55.610 65.690 ;
        RECT 55.260 65.680 55.595 65.685 ;
        RECT 54.635 65.675 55.595 65.680 ;
        RECT 54.635 65.665 55.585 65.675 ;
        RECT 54.635 65.660 55.575 65.665 ;
        RECT 54.635 65.650 55.565 65.660 ;
        RECT 54.635 65.640 55.560 65.650 ;
        RECT 54.635 65.635 55.555 65.640 ;
        RECT 54.635 65.620 55.545 65.635 ;
        RECT 54.635 65.605 55.540 65.620 ;
        RECT 54.635 65.580 55.530 65.605 ;
        RECT 54.635 65.510 55.525 65.580 ;
        RECT 47.585 64.965 47.830 65.415 ;
        RECT 48.000 65.045 48.550 65.245 ;
        RECT 48.720 65.215 48.890 65.415 ;
        RECT 49.665 65.335 50.295 65.505 ;
        RECT 48.720 65.045 49.095 65.215 ;
        RECT 49.265 64.795 49.495 65.295 ;
        RECT 47.245 64.625 49.495 64.795 ;
        RECT 29.740 64.315 32.040 64.485 ;
        RECT 22.350 63.965 25.570 64.135 ;
        RECT 47.295 64.055 47.625 64.445 ;
        RECT 47.795 64.305 47.965 64.625 ;
        RECT 49.665 64.455 49.835 65.335 ;
        RECT 54.635 64.955 55.185 65.340 ;
        RECT 48.135 64.055 48.465 64.445 ;
        RECT 48.880 64.285 49.835 64.455 ;
        RECT 50.005 64.055 50.295 64.890 ;
        RECT 55.355 64.785 55.525 65.510 ;
        RECT 54.635 64.615 55.525 64.785 ;
        RECT 55.695 65.110 56.025 65.535 ;
        RECT 56.195 65.310 56.425 65.705 ;
        RECT 55.695 65.080 55.970 65.110 ;
        RECT 55.695 64.625 55.915 65.080 ;
        RECT 56.595 65.055 56.765 66.085 ;
        RECT 56.085 64.405 56.335 64.945 ;
        RECT 56.505 64.575 56.765 65.055 ;
        RECT 54.550 64.235 56.850 64.405 ;
        RECT 47.160 63.885 50.380 64.055 ;
        RECT 22.840 62.965 25.140 63.135 ;
        RECT 23.125 62.295 23.405 62.965 ;
        RECT 23.575 62.075 23.875 62.625 ;
        RECT 24.075 62.245 24.405 62.965 ;
        RECT 47.650 62.885 49.950 63.055 ;
        RECT 24.595 62.245 25.055 62.795 ;
        RECT 22.940 61.655 23.205 62.015 ;
        RECT 23.575 61.905 24.515 62.075 ;
        RECT 24.345 61.655 24.515 61.905 ;
        RECT 22.940 61.405 23.615 61.655 ;
        RECT 23.835 61.405 24.175 61.655 ;
        RECT 24.345 61.325 24.635 61.655 ;
        RECT 24.345 61.235 24.515 61.325 ;
        RECT 23.125 61.045 24.515 61.235 ;
        RECT 23.125 60.685 23.455 61.045 ;
        RECT 24.805 60.875 25.055 62.245 ;
        RECT 47.935 62.215 48.215 62.885 ;
        RECT 29.720 61.935 32.020 62.105 ;
        RECT 48.385 61.995 48.685 62.545 ;
        RECT 48.885 62.165 49.215 62.885 ;
        RECT 49.405 62.165 49.865 62.715 ;
        RECT 30.005 61.265 30.285 61.935 ;
        RECT 30.455 61.045 30.755 61.595 ;
        RECT 30.955 61.215 31.285 61.935 ;
        RECT 31.475 61.215 31.935 61.765 ;
        RECT 47.750 61.575 48.015 61.935 ;
        RECT 48.385 61.825 49.325 61.995 ;
        RECT 49.155 61.575 49.325 61.825 ;
        RECT 47.750 61.325 48.425 61.575 ;
        RECT 48.645 61.325 48.985 61.575 ;
        RECT 24.075 60.415 24.325 60.875 ;
        RECT 24.495 60.585 25.055 60.875 ;
        RECT 29.820 60.625 30.085 60.985 ;
        RECT 30.455 60.875 31.395 61.045 ;
        RECT 31.225 60.625 31.395 60.875 ;
        RECT 22.840 60.245 25.140 60.415 ;
        RECT 29.820 60.375 30.495 60.625 ;
        RECT 30.715 60.375 31.055 60.625 ;
        RECT 31.225 60.295 31.515 60.625 ;
        RECT 31.225 60.205 31.395 60.295 ;
        RECT 30.005 60.015 31.395 60.205 ;
        RECT 30.005 59.655 30.335 60.015 ;
        RECT 31.685 59.845 31.935 61.215 ;
        RECT 49.155 61.245 49.445 61.575 ;
        RECT 49.155 61.155 49.325 61.245 ;
        RECT 47.935 60.965 49.325 61.155 ;
        RECT 47.935 60.605 48.265 60.965 ;
        RECT 49.615 60.795 49.865 62.165 ;
        RECT 54.530 61.855 56.830 62.025 ;
        RECT 54.815 61.185 55.095 61.855 ;
        RECT 55.265 60.965 55.565 61.515 ;
        RECT 55.765 61.135 56.095 61.855 ;
        RECT 56.285 61.135 56.745 61.685 ;
        RECT 48.885 60.335 49.135 60.795 ;
        RECT 49.305 60.505 49.865 60.795 ;
        RECT 54.630 60.545 54.895 60.905 ;
        RECT 55.265 60.795 56.205 60.965 ;
        RECT 56.035 60.545 56.205 60.795 ;
        RECT 47.650 60.165 49.950 60.335 ;
        RECT 54.630 60.295 55.305 60.545 ;
        RECT 55.525 60.295 55.865 60.545 ;
        RECT 56.035 60.215 56.325 60.545 ;
        RECT 56.035 60.125 56.205 60.215 ;
        RECT 30.955 59.385 31.205 59.845 ;
        RECT 31.375 59.555 31.935 59.845 ;
        RECT 54.815 59.935 56.205 60.125 ;
        RECT 54.815 59.575 55.145 59.935 ;
        RECT 56.495 59.765 56.745 61.135 ;
        RECT 29.720 59.215 32.020 59.385 ;
        RECT 55.765 59.305 56.015 59.765 ;
        RECT 56.185 59.475 56.745 59.765 ;
        RECT 54.530 59.135 56.830 59.305 ;
        RECT 22.400 58.865 25.620 59.035 ;
        RECT 22.485 58.015 22.865 58.695 ;
        RECT 23.455 58.015 23.625 58.865 ;
        RECT 23.795 58.185 24.125 58.695 ;
        RECT 24.295 58.355 24.465 58.865 ;
        RECT 47.210 58.785 50.430 58.955 ;
        RECT 24.635 58.185 25.035 58.695 ;
        RECT 23.795 58.015 25.035 58.185 ;
        RECT 22.485 57.055 22.655 58.015 ;
        RECT 22.825 57.675 24.130 57.845 ;
        RECT 25.215 57.765 25.535 58.695 ;
        RECT 22.825 57.225 23.070 57.675 ;
        RECT 23.240 57.305 23.790 57.505 ;
        RECT 23.960 57.475 24.130 57.675 ;
        RECT 24.905 57.595 25.535 57.765 ;
        RECT 47.295 57.935 47.675 58.615 ;
        RECT 48.265 57.935 48.435 58.785 ;
        RECT 48.605 58.105 48.935 58.615 ;
        RECT 49.105 58.275 49.275 58.785 ;
        RECT 49.445 58.105 49.845 58.615 ;
        RECT 48.605 57.935 49.845 58.105 ;
        RECT 23.960 57.305 24.335 57.475 ;
        RECT 24.505 57.055 24.735 57.555 ;
        RECT 22.485 56.885 24.735 57.055 ;
        RECT 22.535 56.315 22.865 56.705 ;
        RECT 23.035 56.565 23.205 56.885 ;
        RECT 24.905 56.715 25.075 57.595 ;
        RECT 23.375 56.315 23.705 56.705 ;
        RECT 24.120 56.545 25.075 56.715 ;
        RECT 25.245 56.315 25.535 57.150 ;
        RECT 47.295 56.975 47.465 57.935 ;
        RECT 47.635 57.595 48.940 57.765 ;
        RECT 50.025 57.685 50.345 58.615 ;
        RECT 47.635 57.145 47.880 57.595 ;
        RECT 48.050 57.225 48.600 57.425 ;
        RECT 48.770 57.395 48.940 57.595 ;
        RECT 49.715 57.515 50.345 57.685 ;
        RECT 48.770 57.225 49.145 57.395 ;
        RECT 49.315 56.975 49.545 57.475 ;
        RECT 47.295 56.805 49.545 56.975 ;
        RECT 22.400 56.145 25.620 56.315 ;
        RECT 47.345 56.235 47.675 56.625 ;
        RECT 47.845 56.485 48.015 56.805 ;
        RECT 49.715 56.635 49.885 57.515 ;
        RECT 48.185 56.235 48.515 56.625 ;
        RECT 48.930 56.465 49.885 56.635 ;
        RECT 50.055 56.235 50.345 57.070 ;
        RECT 47.210 56.065 50.430 56.235 ;
        RECT 22.890 55.145 25.190 55.315 ;
        RECT 23.175 54.475 23.455 55.145 ;
        RECT 23.625 54.255 23.925 54.805 ;
        RECT 24.125 54.425 24.455 55.145 ;
        RECT 47.700 55.065 50.000 55.235 ;
        RECT 24.645 54.425 25.105 54.975 ;
        RECT 22.990 53.835 23.255 54.195 ;
        RECT 23.625 54.085 24.565 54.255 ;
        RECT 24.395 53.835 24.565 54.085 ;
        RECT 22.990 53.585 23.665 53.835 ;
        RECT 23.885 53.585 24.225 53.835 ;
        RECT 24.395 53.505 24.685 53.835 ;
        RECT 24.395 53.415 24.565 53.505 ;
        RECT 23.175 53.225 24.565 53.415 ;
        RECT 23.175 52.865 23.505 53.225 ;
        RECT 24.855 53.055 25.105 54.425 ;
        RECT 47.985 54.395 48.265 55.065 ;
        RECT 48.435 54.175 48.735 54.725 ;
        RECT 48.935 54.345 49.265 55.065 ;
        RECT 49.455 54.345 49.915 54.895 ;
        RECT 47.800 53.755 48.065 54.115 ;
        RECT 48.435 54.005 49.375 54.175 ;
        RECT 49.205 53.755 49.375 54.005 ;
        RECT 47.800 53.505 48.475 53.755 ;
        RECT 48.695 53.505 49.035 53.755 ;
        RECT 49.205 53.425 49.495 53.755 ;
        RECT 49.205 53.335 49.375 53.425 ;
        RECT 24.125 52.595 24.375 53.055 ;
        RECT 24.545 52.765 25.105 53.055 ;
        RECT 47.985 53.145 49.375 53.335 ;
        RECT 47.985 52.785 48.315 53.145 ;
        RECT 49.665 52.975 49.915 54.345 ;
        RECT 22.890 52.425 25.190 52.595 ;
        RECT 48.935 52.515 49.185 52.975 ;
        RECT 49.355 52.685 49.915 52.975 ;
        RECT 47.700 52.345 50.000 52.515 ;
        RECT 30.560 32.915 31.940 33.085 ;
        RECT 30.890 32.115 31.220 32.745 ;
        RECT 30.890 31.515 31.120 32.115 ;
        RECT 31.390 32.095 31.620 32.915 ;
        RECT 31.290 31.685 31.620 31.925 ;
        RECT 30.890 30.535 31.220 31.515 ;
        RECT 31.390 30.365 31.600 31.505 ;
        RECT 30.560 30.195 31.940 30.365 ;
        RECT 46.090 29.755 53.450 29.925 ;
        RECT 46.210 29.030 46.610 29.585 ;
        RECT 46.855 29.395 47.185 29.755 ;
        RECT 47.355 29.335 48.365 29.585 ;
        RECT 47.355 29.225 47.525 29.335 ;
        RECT 48.195 29.245 48.365 29.335 ;
        RECT 46.785 29.055 47.525 29.225 ;
        RECT 48.700 29.225 48.870 29.585 ;
        RECT 49.040 29.395 49.370 29.755 ;
        RECT 49.540 29.225 49.710 29.585 ;
        RECT 49.880 29.350 50.210 29.755 ;
        RECT 46.210 28.355 46.540 29.030 ;
        RECT 46.785 28.845 46.955 29.055 ;
        RECT 46.710 28.515 46.955 28.845 ;
        RECT 47.990 28.885 48.485 29.075 ;
        RECT 48.700 29.055 49.710 29.225 ;
        RECT 50.480 29.225 50.650 29.585 ;
        RECT 50.820 29.395 51.150 29.755 ;
        RECT 51.320 29.225 51.490 29.585 ;
        RECT 50.480 29.055 51.490 29.225 ;
        RECT 51.740 29.205 52.340 29.585 ;
        RECT 52.605 29.375 52.935 29.755 ;
        RECT 55.440 29.735 62.800 29.905 ;
        RECT 51.740 29.035 52.935 29.205 ;
        RECT 51.740 28.905 51.980 29.035 ;
        RECT 47.125 28.565 47.565 28.805 ;
        RECT 47.990 28.715 48.655 28.885 ;
        RECT 48.825 28.565 49.200 28.885 ;
        RECT 49.495 28.590 50.660 28.875 ;
        RECT 52.765 28.845 52.935 29.035 ;
        RECT 53.105 29.010 53.365 29.585 ;
        RECT 9.180 27.655 16.540 27.825 ;
        RECT 9.300 26.930 9.700 27.485 ;
        RECT 9.945 27.295 10.275 27.655 ;
        RECT 10.445 27.235 11.455 27.485 ;
        RECT 10.445 27.125 10.615 27.235 ;
        RECT 11.285 27.145 11.455 27.235 ;
        RECT 9.875 26.955 10.615 27.125 ;
        RECT 11.790 27.125 11.960 27.485 ;
        RECT 12.130 27.295 12.460 27.655 ;
        RECT 12.630 27.125 12.800 27.485 ;
        RECT 12.970 27.250 13.300 27.655 ;
        RECT 9.300 26.255 9.630 26.930 ;
        RECT 9.875 26.745 10.045 26.955 ;
        RECT 9.800 26.415 10.045 26.745 ;
        RECT 11.080 26.785 11.575 26.975 ;
        RECT 11.790 26.955 12.800 27.125 ;
        RECT 13.570 27.125 13.740 27.485 ;
        RECT 13.910 27.295 14.240 27.655 ;
        RECT 14.410 27.125 14.580 27.485 ;
        RECT 13.570 26.955 14.580 27.125 ;
        RECT 14.830 27.105 15.430 27.485 ;
        RECT 15.695 27.275 16.025 27.655 ;
        RECT 18.530 27.635 25.890 27.805 ;
        RECT 14.830 26.935 16.025 27.105 ;
        RECT 14.830 26.805 15.070 26.935 ;
        RECT 10.215 26.465 10.655 26.705 ;
        RECT 11.080 26.615 11.745 26.785 ;
        RECT 11.915 26.465 12.290 26.785 ;
        RECT 12.585 26.490 13.750 26.775 ;
        RECT 15.855 26.745 16.025 26.935 ;
        RECT 16.195 26.910 16.455 27.485 ;
        RECT 9.300 25.275 9.700 26.255 ;
        RECT 9.875 25.805 10.045 26.415 ;
        RECT 10.485 25.975 10.905 26.295 ;
        RECT 12.585 26.225 12.755 26.490 ;
        RECT 11.135 26.055 12.755 26.225 ;
        RECT 9.875 25.635 10.540 25.805 ;
        RECT 11.135 25.785 11.385 26.055 ;
        RECT 12.980 25.975 13.340 26.305 ;
        RECT 13.580 26.145 13.750 26.490 ;
        RECT 13.920 26.380 14.310 26.710 ;
        RECT 14.500 26.465 14.870 26.635 ;
        RECT 15.300 26.465 15.630 26.745 ;
        RECT 14.500 26.145 14.670 26.465 ;
        RECT 15.460 26.415 15.630 26.465 ;
        RECT 15.855 26.415 16.110 26.745 ;
        RECT 13.580 25.975 14.670 26.145 ;
        RECT 14.840 25.860 15.240 26.295 ;
        RECT 15.855 26.115 16.025 26.415 ;
        RECT 16.280 26.255 16.455 26.910 ;
        RECT 10.370 25.615 10.540 25.635 ;
        RECT 11.790 25.635 12.800 25.805 ;
        RECT 9.870 25.105 10.200 25.465 ;
        RECT 10.370 25.275 11.455 25.615 ;
        RECT 11.790 25.275 11.960 25.635 ;
        RECT 12.130 25.105 12.460 25.465 ;
        RECT 12.630 25.275 12.800 25.635 ;
        RECT 13.505 25.635 14.580 25.805 ;
        RECT 15.435 25.795 16.025 26.115 ;
        RECT 15.435 25.675 15.605 25.795 ;
        RECT 12.970 25.105 13.300 25.485 ;
        RECT 13.505 25.275 13.740 25.635 ;
        RECT 13.910 25.105 14.240 25.465 ;
        RECT 14.410 25.275 14.580 25.635 ;
        RECT 14.830 25.275 15.605 25.675 ;
        RECT 15.775 25.105 16.025 25.590 ;
        RECT 16.195 25.275 16.455 26.255 ;
        RECT 18.650 26.910 19.050 27.465 ;
        RECT 19.295 27.275 19.625 27.635 ;
        RECT 19.795 27.215 20.805 27.465 ;
        RECT 19.795 27.105 19.965 27.215 ;
        RECT 20.635 27.125 20.805 27.215 ;
        RECT 19.225 26.935 19.965 27.105 ;
        RECT 21.140 27.105 21.310 27.465 ;
        RECT 21.480 27.275 21.810 27.635 ;
        RECT 21.980 27.105 22.150 27.465 ;
        RECT 22.320 27.230 22.650 27.635 ;
        RECT 18.650 26.235 18.980 26.910 ;
        RECT 19.225 26.725 19.395 26.935 ;
        RECT 19.150 26.395 19.395 26.725 ;
        RECT 20.430 26.765 20.925 26.955 ;
        RECT 21.140 26.935 22.150 27.105 ;
        RECT 22.920 27.105 23.090 27.465 ;
        RECT 23.260 27.275 23.590 27.635 ;
        RECT 23.760 27.105 23.930 27.465 ;
        RECT 22.920 26.935 23.930 27.105 ;
        RECT 24.180 27.085 24.780 27.465 ;
        RECT 25.045 27.255 25.375 27.635 ;
        RECT 27.610 27.615 34.970 27.785 ;
        RECT 24.180 26.915 25.375 27.085 ;
        RECT 24.180 26.785 24.420 26.915 ;
        RECT 19.565 26.445 20.005 26.685 ;
        RECT 20.430 26.595 21.095 26.765 ;
        RECT 21.265 26.445 21.640 26.765 ;
        RECT 21.935 26.470 23.100 26.755 ;
        RECT 25.205 26.725 25.375 26.915 ;
        RECT 25.545 26.890 25.805 27.465 ;
        RECT 18.650 25.255 19.050 26.235 ;
        RECT 19.225 25.785 19.395 26.395 ;
        RECT 19.835 25.955 20.255 26.275 ;
        RECT 21.935 26.205 22.105 26.470 ;
        RECT 20.485 26.035 22.105 26.205 ;
        RECT 19.225 25.615 19.890 25.785 ;
        RECT 20.485 25.765 20.735 26.035 ;
        RECT 22.330 25.955 22.690 26.285 ;
        RECT 22.930 26.125 23.100 26.470 ;
        RECT 23.270 26.360 23.660 26.690 ;
        RECT 23.850 26.445 24.220 26.615 ;
        RECT 24.650 26.445 24.980 26.725 ;
        RECT 23.850 26.125 24.020 26.445 ;
        RECT 24.810 26.395 24.980 26.445 ;
        RECT 25.205 26.395 25.460 26.725 ;
        RECT 22.930 25.955 24.020 26.125 ;
        RECT 24.190 25.840 24.590 26.275 ;
        RECT 25.205 26.095 25.375 26.395 ;
        RECT 25.630 26.235 25.805 26.890 ;
        RECT 19.720 25.595 19.890 25.615 ;
        RECT 21.140 25.615 22.150 25.785 ;
        RECT 9.180 24.935 16.540 25.105 ;
        RECT 19.220 25.085 19.550 25.445 ;
        RECT 19.720 25.255 20.805 25.595 ;
        RECT 21.140 25.255 21.310 25.615 ;
        RECT 21.480 25.085 21.810 25.445 ;
        RECT 21.980 25.255 22.150 25.615 ;
        RECT 22.855 25.615 23.930 25.785 ;
        RECT 24.785 25.775 25.375 26.095 ;
        RECT 24.785 25.655 24.955 25.775 ;
        RECT 22.320 25.085 22.650 25.465 ;
        RECT 22.855 25.255 23.090 25.615 ;
        RECT 23.260 25.085 23.590 25.445 ;
        RECT 23.760 25.255 23.930 25.615 ;
        RECT 24.180 25.255 24.955 25.655 ;
        RECT 25.125 25.085 25.375 25.570 ;
        RECT 25.545 25.255 25.805 26.235 ;
        RECT 27.730 26.890 28.130 27.445 ;
        RECT 28.375 27.255 28.705 27.615 ;
        RECT 28.875 27.195 29.885 27.445 ;
        RECT 28.875 27.085 29.045 27.195 ;
        RECT 29.715 27.105 29.885 27.195 ;
        RECT 28.305 26.915 29.045 27.085 ;
        RECT 30.220 27.085 30.390 27.445 ;
        RECT 30.560 27.255 30.890 27.615 ;
        RECT 31.060 27.085 31.230 27.445 ;
        RECT 31.400 27.210 31.730 27.615 ;
        RECT 27.730 26.215 28.060 26.890 ;
        RECT 28.305 26.705 28.475 26.915 ;
        RECT 28.230 26.375 28.475 26.705 ;
        RECT 29.510 26.745 30.005 26.935 ;
        RECT 30.220 26.915 31.230 27.085 ;
        RECT 32.000 27.085 32.170 27.445 ;
        RECT 32.340 27.255 32.670 27.615 ;
        RECT 32.840 27.085 33.010 27.445 ;
        RECT 32.000 26.915 33.010 27.085 ;
        RECT 33.260 27.065 33.860 27.445 ;
        RECT 34.125 27.235 34.455 27.615 ;
        RECT 36.960 27.595 44.320 27.765 ;
        RECT 33.260 26.895 34.455 27.065 ;
        RECT 33.260 26.765 33.500 26.895 ;
        RECT 28.645 26.425 29.085 26.665 ;
        RECT 29.510 26.575 30.175 26.745 ;
        RECT 30.345 26.425 30.720 26.745 ;
        RECT 31.015 26.450 32.180 26.735 ;
        RECT 34.285 26.705 34.455 26.895 ;
        RECT 34.625 26.870 34.885 27.445 ;
        RECT 27.730 25.235 28.130 26.215 ;
        RECT 28.305 25.765 28.475 26.375 ;
        RECT 28.915 25.935 29.335 26.255 ;
        RECT 31.015 26.185 31.185 26.450 ;
        RECT 29.565 26.015 31.185 26.185 ;
        RECT 28.305 25.595 28.970 25.765 ;
        RECT 29.565 25.745 29.815 26.015 ;
        RECT 31.410 25.935 31.770 26.265 ;
        RECT 32.010 26.105 32.180 26.450 ;
        RECT 32.350 26.340 32.740 26.670 ;
        RECT 32.930 26.425 33.300 26.595 ;
        RECT 33.730 26.425 34.060 26.705 ;
        RECT 32.930 26.105 33.100 26.425 ;
        RECT 33.890 26.375 34.060 26.425 ;
        RECT 34.285 26.375 34.540 26.705 ;
        RECT 32.010 25.935 33.100 26.105 ;
        RECT 33.270 25.820 33.670 26.255 ;
        RECT 34.285 26.075 34.455 26.375 ;
        RECT 34.710 26.215 34.885 26.870 ;
        RECT 28.800 25.575 28.970 25.595 ;
        RECT 30.220 25.595 31.230 25.765 ;
        RECT 18.530 24.915 25.890 25.085 ;
        RECT 28.300 25.065 28.630 25.425 ;
        RECT 28.800 25.235 29.885 25.575 ;
        RECT 30.220 25.235 30.390 25.595 ;
        RECT 30.560 25.065 30.890 25.425 ;
        RECT 31.060 25.235 31.230 25.595 ;
        RECT 31.935 25.595 33.010 25.765 ;
        RECT 33.865 25.755 34.455 26.075 ;
        RECT 33.865 25.635 34.035 25.755 ;
        RECT 31.400 25.065 31.730 25.445 ;
        RECT 31.935 25.235 32.170 25.595 ;
        RECT 32.340 25.065 32.670 25.425 ;
        RECT 32.840 25.235 33.010 25.595 ;
        RECT 33.260 25.235 34.035 25.635 ;
        RECT 34.205 25.065 34.455 25.550 ;
        RECT 34.625 25.235 34.885 26.215 ;
        RECT 37.080 26.870 37.480 27.425 ;
        RECT 37.725 27.235 38.055 27.595 ;
        RECT 38.225 27.175 39.235 27.425 ;
        RECT 38.225 27.065 38.395 27.175 ;
        RECT 39.065 27.085 39.235 27.175 ;
        RECT 37.655 26.895 38.395 27.065 ;
        RECT 39.570 27.065 39.740 27.425 ;
        RECT 39.910 27.235 40.240 27.595 ;
        RECT 40.410 27.065 40.580 27.425 ;
        RECT 40.750 27.190 41.080 27.595 ;
        RECT 37.080 26.195 37.410 26.870 ;
        RECT 37.655 26.685 37.825 26.895 ;
        RECT 37.580 26.355 37.825 26.685 ;
        RECT 38.860 26.725 39.355 26.915 ;
        RECT 39.570 26.895 40.580 27.065 ;
        RECT 41.350 27.065 41.520 27.425 ;
        RECT 41.690 27.235 42.020 27.595 ;
        RECT 42.190 27.065 42.360 27.425 ;
        RECT 41.350 26.895 42.360 27.065 ;
        RECT 42.610 27.045 43.210 27.425 ;
        RECT 43.475 27.215 43.805 27.595 ;
        RECT 42.610 26.875 43.805 27.045 ;
        RECT 42.610 26.745 42.850 26.875 ;
        RECT 37.995 26.405 38.435 26.645 ;
        RECT 38.860 26.555 39.525 26.725 ;
        RECT 39.695 26.405 40.070 26.725 ;
        RECT 40.365 26.430 41.530 26.715 ;
        RECT 43.635 26.685 43.805 26.875 ;
        RECT 43.975 26.850 44.235 27.425 ;
        RECT 46.210 27.375 46.610 28.355 ;
        RECT 46.785 27.905 46.955 28.515 ;
        RECT 47.395 28.075 47.815 28.395 ;
        RECT 49.495 28.325 49.665 28.590 ;
        RECT 48.045 28.155 49.665 28.325 ;
        RECT 46.785 27.735 47.450 27.905 ;
        RECT 48.045 27.885 48.295 28.155 ;
        RECT 49.890 28.075 50.250 28.405 ;
        RECT 50.490 28.245 50.660 28.590 ;
        RECT 50.830 28.480 51.220 28.810 ;
        RECT 51.410 28.565 51.780 28.735 ;
        RECT 52.210 28.565 52.540 28.845 ;
        RECT 51.410 28.245 51.580 28.565 ;
        RECT 52.370 28.515 52.540 28.565 ;
        RECT 52.765 28.515 53.020 28.845 ;
        RECT 50.490 28.075 51.580 28.245 ;
        RECT 51.750 27.960 52.150 28.395 ;
        RECT 52.765 28.215 52.935 28.515 ;
        RECT 53.190 28.355 53.365 29.010 ;
        RECT 47.280 27.715 47.450 27.735 ;
        RECT 48.700 27.735 49.710 27.905 ;
        RECT 46.780 27.205 47.110 27.565 ;
        RECT 47.280 27.375 48.365 27.715 ;
        RECT 48.700 27.375 48.870 27.735 ;
        RECT 49.040 27.205 49.370 27.565 ;
        RECT 49.540 27.375 49.710 27.735 ;
        RECT 50.415 27.735 51.490 27.905 ;
        RECT 52.345 27.895 52.935 28.215 ;
        RECT 52.345 27.775 52.515 27.895 ;
        RECT 49.880 27.205 50.210 27.585 ;
        RECT 50.415 27.375 50.650 27.735 ;
        RECT 50.820 27.205 51.150 27.565 ;
        RECT 51.320 27.375 51.490 27.735 ;
        RECT 51.740 27.375 52.515 27.775 ;
        RECT 52.685 27.205 52.935 27.690 ;
        RECT 53.105 27.375 53.365 28.355 ;
        RECT 55.560 29.010 55.960 29.565 ;
        RECT 56.205 29.375 56.535 29.735 ;
        RECT 56.705 29.315 57.715 29.565 ;
        RECT 56.705 29.205 56.875 29.315 ;
        RECT 57.545 29.225 57.715 29.315 ;
        RECT 56.135 29.035 56.875 29.205 ;
        RECT 58.050 29.205 58.220 29.565 ;
        RECT 58.390 29.375 58.720 29.735 ;
        RECT 58.890 29.205 59.060 29.565 ;
        RECT 59.230 29.330 59.560 29.735 ;
        RECT 55.560 28.335 55.890 29.010 ;
        RECT 56.135 28.825 56.305 29.035 ;
        RECT 56.060 28.495 56.305 28.825 ;
        RECT 57.340 28.865 57.835 29.055 ;
        RECT 58.050 29.035 59.060 29.205 ;
        RECT 59.830 29.205 60.000 29.565 ;
        RECT 60.170 29.375 60.500 29.735 ;
        RECT 60.670 29.205 60.840 29.565 ;
        RECT 59.830 29.035 60.840 29.205 ;
        RECT 61.090 29.185 61.690 29.565 ;
        RECT 61.955 29.355 62.285 29.735 ;
        RECT 64.520 29.715 71.880 29.885 ;
        RECT 61.090 29.015 62.285 29.185 ;
        RECT 61.090 28.885 61.330 29.015 ;
        RECT 56.475 28.545 56.915 28.785 ;
        RECT 57.340 28.695 58.005 28.865 ;
        RECT 58.175 28.545 58.550 28.865 ;
        RECT 58.845 28.570 60.010 28.855 ;
        RECT 62.115 28.825 62.285 29.015 ;
        RECT 62.455 28.990 62.715 29.565 ;
        RECT 55.560 27.355 55.960 28.335 ;
        RECT 56.135 27.885 56.305 28.495 ;
        RECT 56.745 28.055 57.165 28.375 ;
        RECT 58.845 28.305 59.015 28.570 ;
        RECT 57.395 28.135 59.015 28.305 ;
        RECT 56.135 27.715 56.800 27.885 ;
        RECT 57.395 27.865 57.645 28.135 ;
        RECT 59.240 28.055 59.600 28.385 ;
        RECT 59.840 28.225 60.010 28.570 ;
        RECT 60.180 28.460 60.570 28.790 ;
        RECT 60.760 28.545 61.130 28.715 ;
        RECT 61.560 28.545 61.890 28.825 ;
        RECT 60.760 28.225 60.930 28.545 ;
        RECT 61.720 28.495 61.890 28.545 ;
        RECT 62.115 28.495 62.370 28.825 ;
        RECT 59.840 28.055 60.930 28.225 ;
        RECT 61.100 27.940 61.500 28.375 ;
        RECT 62.115 28.195 62.285 28.495 ;
        RECT 62.540 28.335 62.715 28.990 ;
        RECT 56.630 27.695 56.800 27.715 ;
        RECT 58.050 27.715 59.060 27.885 ;
        RECT 46.090 27.035 53.450 27.205 ;
        RECT 56.130 27.185 56.460 27.545 ;
        RECT 56.630 27.355 57.715 27.695 ;
        RECT 58.050 27.355 58.220 27.715 ;
        RECT 58.390 27.185 58.720 27.545 ;
        RECT 58.890 27.355 59.060 27.715 ;
        RECT 59.765 27.715 60.840 27.885 ;
        RECT 61.695 27.875 62.285 28.195 ;
        RECT 61.695 27.755 61.865 27.875 ;
        RECT 59.230 27.185 59.560 27.565 ;
        RECT 59.765 27.355 60.000 27.715 ;
        RECT 60.170 27.185 60.500 27.545 ;
        RECT 60.670 27.355 60.840 27.715 ;
        RECT 61.090 27.355 61.865 27.755 ;
        RECT 62.035 27.185 62.285 27.670 ;
        RECT 62.455 27.355 62.715 28.335 ;
        RECT 64.640 28.990 65.040 29.545 ;
        RECT 65.285 29.355 65.615 29.715 ;
        RECT 65.785 29.295 66.795 29.545 ;
        RECT 65.785 29.185 65.955 29.295 ;
        RECT 66.625 29.205 66.795 29.295 ;
        RECT 65.215 29.015 65.955 29.185 ;
        RECT 67.130 29.185 67.300 29.545 ;
        RECT 67.470 29.355 67.800 29.715 ;
        RECT 67.970 29.185 68.140 29.545 ;
        RECT 68.310 29.310 68.640 29.715 ;
        RECT 64.640 28.315 64.970 28.990 ;
        RECT 65.215 28.805 65.385 29.015 ;
        RECT 65.140 28.475 65.385 28.805 ;
        RECT 66.420 28.845 66.915 29.035 ;
        RECT 67.130 29.015 68.140 29.185 ;
        RECT 68.910 29.185 69.080 29.545 ;
        RECT 69.250 29.355 69.580 29.715 ;
        RECT 69.750 29.185 69.920 29.545 ;
        RECT 68.910 29.015 69.920 29.185 ;
        RECT 70.170 29.165 70.770 29.545 ;
        RECT 71.035 29.335 71.365 29.715 ;
        RECT 73.870 29.695 81.230 29.865 ;
        RECT 70.170 28.995 71.365 29.165 ;
        RECT 70.170 28.865 70.410 28.995 ;
        RECT 65.555 28.525 65.995 28.765 ;
        RECT 66.420 28.675 67.085 28.845 ;
        RECT 67.255 28.525 67.630 28.845 ;
        RECT 67.925 28.550 69.090 28.835 ;
        RECT 71.195 28.805 71.365 28.995 ;
        RECT 71.535 28.970 71.795 29.545 ;
        RECT 64.640 27.335 65.040 28.315 ;
        RECT 65.215 27.865 65.385 28.475 ;
        RECT 65.825 28.035 66.245 28.355 ;
        RECT 67.925 28.285 68.095 28.550 ;
        RECT 66.475 28.115 68.095 28.285 ;
        RECT 65.215 27.695 65.880 27.865 ;
        RECT 66.475 27.845 66.725 28.115 ;
        RECT 68.320 28.035 68.680 28.365 ;
        RECT 68.920 28.205 69.090 28.550 ;
        RECT 69.260 28.440 69.650 28.770 ;
        RECT 69.840 28.525 70.210 28.695 ;
        RECT 70.640 28.525 70.970 28.805 ;
        RECT 69.840 28.205 70.010 28.525 ;
        RECT 70.800 28.475 70.970 28.525 ;
        RECT 71.195 28.475 71.450 28.805 ;
        RECT 68.920 28.035 70.010 28.205 ;
        RECT 70.180 27.920 70.580 28.355 ;
        RECT 71.195 28.175 71.365 28.475 ;
        RECT 71.620 28.315 71.795 28.970 ;
        RECT 65.710 27.675 65.880 27.695 ;
        RECT 67.130 27.695 68.140 27.865 ;
        RECT 55.440 27.015 62.800 27.185 ;
        RECT 65.210 27.165 65.540 27.525 ;
        RECT 65.710 27.335 66.795 27.675 ;
        RECT 67.130 27.335 67.300 27.695 ;
        RECT 67.470 27.165 67.800 27.525 ;
        RECT 67.970 27.335 68.140 27.695 ;
        RECT 68.845 27.695 69.920 27.865 ;
        RECT 70.775 27.855 71.365 28.175 ;
        RECT 70.775 27.735 70.945 27.855 ;
        RECT 68.310 27.165 68.640 27.545 ;
        RECT 68.845 27.335 69.080 27.695 ;
        RECT 69.250 27.165 69.580 27.525 ;
        RECT 69.750 27.335 69.920 27.695 ;
        RECT 70.170 27.335 70.945 27.735 ;
        RECT 71.115 27.165 71.365 27.650 ;
        RECT 71.535 27.335 71.795 28.315 ;
        RECT 73.990 28.970 74.390 29.525 ;
        RECT 74.635 29.335 74.965 29.695 ;
        RECT 75.135 29.275 76.145 29.525 ;
        RECT 75.135 29.165 75.305 29.275 ;
        RECT 75.975 29.185 76.145 29.275 ;
        RECT 74.565 28.995 75.305 29.165 ;
        RECT 76.480 29.165 76.650 29.525 ;
        RECT 76.820 29.335 77.150 29.695 ;
        RECT 77.320 29.165 77.490 29.525 ;
        RECT 77.660 29.290 77.990 29.695 ;
        RECT 73.990 28.295 74.320 28.970 ;
        RECT 74.565 28.785 74.735 28.995 ;
        RECT 74.490 28.455 74.735 28.785 ;
        RECT 75.770 28.825 76.265 29.015 ;
        RECT 76.480 28.995 77.490 29.165 ;
        RECT 78.260 29.165 78.430 29.525 ;
        RECT 78.600 29.335 78.930 29.695 ;
        RECT 79.100 29.165 79.270 29.525 ;
        RECT 78.260 28.995 79.270 29.165 ;
        RECT 79.520 29.145 80.120 29.525 ;
        RECT 80.385 29.315 80.715 29.695 ;
        RECT 79.520 28.975 80.715 29.145 ;
        RECT 79.520 28.845 79.760 28.975 ;
        RECT 74.905 28.505 75.345 28.745 ;
        RECT 75.770 28.655 76.435 28.825 ;
        RECT 76.605 28.505 76.980 28.825 ;
        RECT 77.275 28.530 78.440 28.815 ;
        RECT 80.545 28.785 80.715 28.975 ;
        RECT 80.885 28.950 81.145 29.525 ;
        RECT 73.990 27.315 74.390 28.295 ;
        RECT 74.565 27.845 74.735 28.455 ;
        RECT 75.175 28.015 75.595 28.335 ;
        RECT 77.275 28.265 77.445 28.530 ;
        RECT 75.825 28.095 77.445 28.265 ;
        RECT 74.565 27.675 75.230 27.845 ;
        RECT 75.825 27.825 76.075 28.095 ;
        RECT 77.670 28.015 78.030 28.345 ;
        RECT 78.270 28.185 78.440 28.530 ;
        RECT 78.610 28.420 79.000 28.750 ;
        RECT 79.190 28.505 79.560 28.675 ;
        RECT 79.990 28.505 80.320 28.785 ;
        RECT 79.190 28.185 79.360 28.505 ;
        RECT 80.150 28.455 80.320 28.505 ;
        RECT 80.545 28.455 80.800 28.785 ;
        RECT 78.270 28.015 79.360 28.185 ;
        RECT 79.530 27.900 79.930 28.335 ;
        RECT 80.545 28.155 80.715 28.455 ;
        RECT 80.970 28.295 81.145 28.950 ;
        RECT 75.060 27.655 75.230 27.675 ;
        RECT 76.480 27.675 77.490 27.845 ;
        RECT 64.520 26.995 71.880 27.165 ;
        RECT 74.560 27.145 74.890 27.505 ;
        RECT 75.060 27.315 76.145 27.655 ;
        RECT 76.480 27.315 76.650 27.675 ;
        RECT 76.820 27.145 77.150 27.505 ;
        RECT 77.320 27.315 77.490 27.675 ;
        RECT 78.195 27.675 79.270 27.845 ;
        RECT 80.125 27.835 80.715 28.155 ;
        RECT 80.125 27.715 80.295 27.835 ;
        RECT 77.660 27.145 77.990 27.525 ;
        RECT 78.195 27.315 78.430 27.675 ;
        RECT 78.600 27.145 78.930 27.505 ;
        RECT 79.100 27.315 79.270 27.675 ;
        RECT 79.520 27.315 80.295 27.715 ;
        RECT 80.465 27.145 80.715 27.630 ;
        RECT 80.885 27.315 81.145 28.295 ;
        RECT 73.870 26.975 81.230 27.145 ;
        RECT 84.010 26.895 88.150 27.065 ;
        RECT 37.080 25.215 37.480 26.195 ;
        RECT 37.655 25.745 37.825 26.355 ;
        RECT 38.265 25.915 38.685 26.235 ;
        RECT 40.365 26.165 40.535 26.430 ;
        RECT 38.915 25.995 40.535 26.165 ;
        RECT 37.655 25.575 38.320 25.745 ;
        RECT 38.915 25.725 39.165 25.995 ;
        RECT 40.760 25.915 41.120 26.245 ;
        RECT 41.360 26.085 41.530 26.430 ;
        RECT 41.700 26.320 42.090 26.650 ;
        RECT 42.280 26.405 42.650 26.575 ;
        RECT 43.080 26.405 43.410 26.685 ;
        RECT 42.280 26.085 42.450 26.405 ;
        RECT 43.240 26.355 43.410 26.405 ;
        RECT 43.635 26.355 43.890 26.685 ;
        RECT 41.360 25.915 42.450 26.085 ;
        RECT 42.620 25.800 43.020 26.235 ;
        RECT 43.635 26.055 43.805 26.355 ;
        RECT 44.060 26.195 44.235 26.850 ;
        RECT 38.150 25.555 38.320 25.575 ;
        RECT 39.570 25.575 40.580 25.745 ;
        RECT 27.610 24.895 34.970 25.065 ;
        RECT 37.650 25.045 37.980 25.405 ;
        RECT 38.150 25.215 39.235 25.555 ;
        RECT 39.570 25.215 39.740 25.575 ;
        RECT 39.910 25.045 40.240 25.405 ;
        RECT 40.410 25.215 40.580 25.575 ;
        RECT 41.285 25.575 42.360 25.745 ;
        RECT 43.215 25.735 43.805 26.055 ;
        RECT 43.215 25.615 43.385 25.735 ;
        RECT 40.750 25.045 41.080 25.425 ;
        RECT 41.285 25.215 41.520 25.575 ;
        RECT 41.690 25.045 42.020 25.405 ;
        RECT 42.190 25.215 42.360 25.575 ;
        RECT 42.610 25.215 43.385 25.615 ;
        RECT 43.555 25.045 43.805 25.530 ;
        RECT 43.975 25.215 44.235 26.195 ;
        RECT 84.370 26.085 84.615 26.690 ;
        RECT 84.835 26.360 85.345 26.895 ;
        RECT 84.095 25.915 85.325 26.085 ;
        RECT 46.230 25.385 53.590 25.555 ;
        RECT 36.960 24.875 44.320 25.045 ;
        RECT 46.350 24.660 46.750 25.215 ;
        RECT 46.995 25.025 47.325 25.385 ;
        RECT 47.495 24.965 48.505 25.215 ;
        RECT 47.495 24.855 47.665 24.965 ;
        RECT 48.335 24.875 48.505 24.965 ;
        RECT 46.925 24.685 47.665 24.855 ;
        RECT 48.840 24.855 49.010 25.215 ;
        RECT 49.180 25.025 49.510 25.385 ;
        RECT 49.680 24.855 49.850 25.215 ;
        RECT 50.020 24.980 50.350 25.385 ;
        RECT 46.350 23.985 46.680 24.660 ;
        RECT 46.925 24.475 47.095 24.685 ;
        RECT 46.850 24.145 47.095 24.475 ;
        RECT 48.130 24.515 48.625 24.705 ;
        RECT 48.840 24.685 49.850 24.855 ;
        RECT 50.620 24.855 50.790 25.215 ;
        RECT 50.960 25.025 51.290 25.385 ;
        RECT 51.460 24.855 51.630 25.215 ;
        RECT 50.620 24.685 51.630 24.855 ;
        RECT 51.880 24.835 52.480 25.215 ;
        RECT 52.745 25.005 53.075 25.385 ;
        RECT 55.580 25.365 62.940 25.535 ;
        RECT 51.880 24.665 53.075 24.835 ;
        RECT 51.880 24.535 52.120 24.665 ;
        RECT 47.265 24.195 47.705 24.435 ;
        RECT 48.130 24.345 48.795 24.515 ;
        RECT 48.965 24.195 49.340 24.515 ;
        RECT 49.635 24.220 50.800 24.505 ;
        RECT 52.905 24.475 53.075 24.665 ;
        RECT 53.245 24.640 53.505 25.215 ;
        RECT 46.350 23.005 46.750 23.985 ;
        RECT 46.925 23.535 47.095 24.145 ;
        RECT 47.535 23.705 47.955 24.025 ;
        RECT 49.635 23.955 49.805 24.220 ;
        RECT 48.185 23.785 49.805 23.955 ;
        RECT 46.925 23.365 47.590 23.535 ;
        RECT 48.185 23.515 48.435 23.785 ;
        RECT 50.030 23.705 50.390 24.035 ;
        RECT 50.630 23.875 50.800 24.220 ;
        RECT 50.970 24.110 51.360 24.440 ;
        RECT 51.550 24.195 51.920 24.365 ;
        RECT 52.350 24.195 52.680 24.475 ;
        RECT 51.550 23.875 51.720 24.195 ;
        RECT 52.510 24.145 52.680 24.195 ;
        RECT 52.905 24.145 53.160 24.475 ;
        RECT 50.630 23.705 51.720 23.875 ;
        RECT 51.890 23.590 52.290 24.025 ;
        RECT 52.905 23.845 53.075 24.145 ;
        RECT 53.330 23.985 53.505 24.640 ;
        RECT 47.420 23.345 47.590 23.365 ;
        RECT 48.840 23.365 49.850 23.535 ;
        RECT 46.920 22.835 47.250 23.195 ;
        RECT 47.420 23.005 48.505 23.345 ;
        RECT 48.840 23.005 49.010 23.365 ;
        RECT 49.180 22.835 49.510 23.195 ;
        RECT 49.680 23.005 49.850 23.365 ;
        RECT 50.555 23.365 51.630 23.535 ;
        RECT 52.485 23.525 53.075 23.845 ;
        RECT 52.485 23.405 52.655 23.525 ;
        RECT 50.020 22.835 50.350 23.215 ;
        RECT 50.555 23.005 50.790 23.365 ;
        RECT 50.960 22.835 51.290 23.195 ;
        RECT 51.460 23.005 51.630 23.365 ;
        RECT 51.880 23.005 52.655 23.405 ;
        RECT 52.825 22.835 53.075 23.320 ;
        RECT 53.245 23.005 53.505 23.985 ;
        RECT 55.700 24.640 56.100 25.195 ;
        RECT 56.345 25.005 56.675 25.365 ;
        RECT 56.845 24.945 57.855 25.195 ;
        RECT 56.845 24.835 57.015 24.945 ;
        RECT 57.685 24.855 57.855 24.945 ;
        RECT 56.275 24.665 57.015 24.835 ;
        RECT 58.190 24.835 58.360 25.195 ;
        RECT 58.530 25.005 58.860 25.365 ;
        RECT 59.030 24.835 59.200 25.195 ;
        RECT 59.370 24.960 59.700 25.365 ;
        RECT 55.700 23.965 56.030 24.640 ;
        RECT 56.275 24.455 56.445 24.665 ;
        RECT 56.200 24.125 56.445 24.455 ;
        RECT 57.480 24.495 57.975 24.685 ;
        RECT 58.190 24.665 59.200 24.835 ;
        RECT 59.970 24.835 60.140 25.195 ;
        RECT 60.310 25.005 60.640 25.365 ;
        RECT 60.810 24.835 60.980 25.195 ;
        RECT 59.970 24.665 60.980 24.835 ;
        RECT 61.230 24.815 61.830 25.195 ;
        RECT 62.095 24.985 62.425 25.365 ;
        RECT 64.660 25.345 72.020 25.515 ;
        RECT 61.230 24.645 62.425 24.815 ;
        RECT 61.230 24.515 61.470 24.645 ;
        RECT 56.615 24.175 57.055 24.415 ;
        RECT 57.480 24.325 58.145 24.495 ;
        RECT 58.315 24.175 58.690 24.495 ;
        RECT 58.985 24.200 60.150 24.485 ;
        RECT 62.255 24.455 62.425 24.645 ;
        RECT 62.595 24.620 62.855 25.195 ;
        RECT 55.700 22.985 56.100 23.965 ;
        RECT 56.275 23.515 56.445 24.125 ;
        RECT 56.885 23.685 57.305 24.005 ;
        RECT 58.985 23.935 59.155 24.200 ;
        RECT 57.535 23.765 59.155 23.935 ;
        RECT 56.275 23.345 56.940 23.515 ;
        RECT 57.535 23.495 57.785 23.765 ;
        RECT 59.380 23.685 59.740 24.015 ;
        RECT 59.980 23.855 60.150 24.200 ;
        RECT 60.320 24.090 60.710 24.420 ;
        RECT 60.900 24.175 61.270 24.345 ;
        RECT 61.700 24.175 62.030 24.455 ;
        RECT 60.900 23.855 61.070 24.175 ;
        RECT 61.860 24.125 62.030 24.175 ;
        RECT 62.255 24.125 62.510 24.455 ;
        RECT 59.980 23.685 61.070 23.855 ;
        RECT 61.240 23.570 61.640 24.005 ;
        RECT 62.255 23.825 62.425 24.125 ;
        RECT 62.680 23.965 62.855 24.620 ;
        RECT 56.770 23.325 56.940 23.345 ;
        RECT 58.190 23.345 59.200 23.515 ;
        RECT 46.230 22.665 53.590 22.835 ;
        RECT 56.270 22.815 56.600 23.175 ;
        RECT 56.770 22.985 57.855 23.325 ;
        RECT 58.190 22.985 58.360 23.345 ;
        RECT 58.530 22.815 58.860 23.175 ;
        RECT 59.030 22.985 59.200 23.345 ;
        RECT 59.905 23.345 60.980 23.515 ;
        RECT 61.835 23.505 62.425 23.825 ;
        RECT 61.835 23.385 62.005 23.505 ;
        RECT 59.370 22.815 59.700 23.195 ;
        RECT 59.905 22.985 60.140 23.345 ;
        RECT 60.310 22.815 60.640 23.175 ;
        RECT 60.810 22.985 60.980 23.345 ;
        RECT 61.230 22.985 62.005 23.385 ;
        RECT 62.175 22.815 62.425 23.300 ;
        RECT 62.595 22.985 62.855 23.965 ;
        RECT 64.780 24.620 65.180 25.175 ;
        RECT 65.425 24.985 65.755 25.345 ;
        RECT 65.925 24.925 66.935 25.175 ;
        RECT 65.925 24.815 66.095 24.925 ;
        RECT 66.765 24.835 66.935 24.925 ;
        RECT 65.355 24.645 66.095 24.815 ;
        RECT 67.270 24.815 67.440 25.175 ;
        RECT 67.610 24.985 67.940 25.345 ;
        RECT 68.110 24.815 68.280 25.175 ;
        RECT 68.450 24.940 68.780 25.345 ;
        RECT 64.780 23.945 65.110 24.620 ;
        RECT 65.355 24.435 65.525 24.645 ;
        RECT 65.280 24.105 65.525 24.435 ;
        RECT 66.560 24.475 67.055 24.665 ;
        RECT 67.270 24.645 68.280 24.815 ;
        RECT 69.050 24.815 69.220 25.175 ;
        RECT 69.390 24.985 69.720 25.345 ;
        RECT 69.890 24.815 70.060 25.175 ;
        RECT 69.050 24.645 70.060 24.815 ;
        RECT 70.310 24.795 70.910 25.175 ;
        RECT 71.175 24.965 71.505 25.345 ;
        RECT 74.010 25.325 81.370 25.495 ;
        RECT 70.310 24.625 71.505 24.795 ;
        RECT 70.310 24.495 70.550 24.625 ;
        RECT 65.695 24.155 66.135 24.395 ;
        RECT 66.560 24.305 67.225 24.475 ;
        RECT 67.395 24.155 67.770 24.475 ;
        RECT 68.065 24.180 69.230 24.465 ;
        RECT 71.335 24.435 71.505 24.625 ;
        RECT 71.675 24.600 71.935 25.175 ;
        RECT 64.780 22.965 65.180 23.945 ;
        RECT 65.355 23.495 65.525 24.105 ;
        RECT 65.965 23.665 66.385 23.985 ;
        RECT 68.065 23.915 68.235 24.180 ;
        RECT 66.615 23.745 68.235 23.915 ;
        RECT 65.355 23.325 66.020 23.495 ;
        RECT 66.615 23.475 66.865 23.745 ;
        RECT 68.460 23.665 68.820 23.995 ;
        RECT 69.060 23.835 69.230 24.180 ;
        RECT 69.400 24.070 69.790 24.400 ;
        RECT 69.980 24.155 70.350 24.325 ;
        RECT 70.780 24.155 71.110 24.435 ;
        RECT 69.980 23.835 70.150 24.155 ;
        RECT 70.940 24.105 71.110 24.155 ;
        RECT 71.335 24.105 71.590 24.435 ;
        RECT 69.060 23.665 70.150 23.835 ;
        RECT 70.320 23.550 70.720 23.985 ;
        RECT 71.335 23.805 71.505 24.105 ;
        RECT 71.760 23.945 71.935 24.600 ;
        RECT 65.850 23.305 66.020 23.325 ;
        RECT 67.270 23.325 68.280 23.495 ;
        RECT 55.580 22.645 62.940 22.815 ;
        RECT 65.350 22.795 65.680 23.155 ;
        RECT 65.850 22.965 66.935 23.305 ;
        RECT 67.270 22.965 67.440 23.325 ;
        RECT 67.610 22.795 67.940 23.155 ;
        RECT 68.110 22.965 68.280 23.325 ;
        RECT 68.985 23.325 70.060 23.495 ;
        RECT 70.915 23.485 71.505 23.805 ;
        RECT 70.915 23.365 71.085 23.485 ;
        RECT 68.450 22.795 68.780 23.175 ;
        RECT 68.985 22.965 69.220 23.325 ;
        RECT 69.390 22.795 69.720 23.155 ;
        RECT 69.890 22.965 70.060 23.325 ;
        RECT 70.310 22.965 71.085 23.365 ;
        RECT 71.255 22.795 71.505 23.280 ;
        RECT 71.675 22.965 71.935 23.945 ;
        RECT 74.130 24.600 74.530 25.155 ;
        RECT 74.775 24.965 75.105 25.325 ;
        RECT 75.275 24.905 76.285 25.155 ;
        RECT 75.275 24.795 75.445 24.905 ;
        RECT 76.115 24.815 76.285 24.905 ;
        RECT 74.705 24.625 75.445 24.795 ;
        RECT 76.620 24.795 76.790 25.155 ;
        RECT 76.960 24.965 77.290 25.325 ;
        RECT 77.460 24.795 77.630 25.155 ;
        RECT 77.800 24.920 78.130 25.325 ;
        RECT 74.130 23.925 74.460 24.600 ;
        RECT 74.705 24.415 74.875 24.625 ;
        RECT 74.630 24.085 74.875 24.415 ;
        RECT 75.910 24.455 76.405 24.645 ;
        RECT 76.620 24.625 77.630 24.795 ;
        RECT 78.400 24.795 78.570 25.155 ;
        RECT 78.740 24.965 79.070 25.325 ;
        RECT 79.240 24.795 79.410 25.155 ;
        RECT 78.400 24.625 79.410 24.795 ;
        RECT 79.660 24.775 80.260 25.155 ;
        RECT 80.525 24.945 80.855 25.325 ;
        RECT 79.660 24.605 80.855 24.775 ;
        RECT 79.660 24.475 79.900 24.605 ;
        RECT 75.045 24.135 75.485 24.375 ;
        RECT 75.910 24.285 76.575 24.455 ;
        RECT 76.745 24.135 77.120 24.455 ;
        RECT 77.415 24.160 78.580 24.445 ;
        RECT 80.685 24.415 80.855 24.605 ;
        RECT 81.025 24.580 81.285 25.155 ;
        RECT 84.095 25.105 84.435 25.915 ;
        RECT 84.605 25.350 85.355 25.540 ;
        RECT 84.095 24.695 84.610 25.105 ;
        RECT 74.130 22.945 74.530 23.925 ;
        RECT 74.705 23.475 74.875 24.085 ;
        RECT 75.315 23.645 75.735 23.965 ;
        RECT 77.415 23.895 77.585 24.160 ;
        RECT 75.965 23.725 77.585 23.895 ;
        RECT 74.705 23.305 75.370 23.475 ;
        RECT 75.965 23.455 76.215 23.725 ;
        RECT 77.810 23.645 78.170 23.975 ;
        RECT 78.410 23.815 78.580 24.160 ;
        RECT 78.750 24.050 79.140 24.380 ;
        RECT 79.330 24.135 79.700 24.305 ;
        RECT 80.130 24.135 80.460 24.415 ;
        RECT 79.330 23.815 79.500 24.135 ;
        RECT 80.290 24.085 80.460 24.135 ;
        RECT 80.685 24.085 80.940 24.415 ;
        RECT 78.410 23.645 79.500 23.815 ;
        RECT 79.670 23.530 80.070 23.965 ;
        RECT 80.685 23.785 80.855 24.085 ;
        RECT 81.110 23.925 81.285 24.580 ;
        RECT 84.845 24.345 85.015 25.105 ;
        RECT 85.185 24.685 85.355 25.350 ;
        RECT 85.525 25.365 85.715 26.725 ;
        RECT 85.885 25.565 86.160 26.725 ;
        RECT 86.350 26.360 86.880 26.725 ;
        RECT 87.305 26.495 87.635 26.895 ;
        RECT 86.705 26.325 86.880 26.360 ;
        RECT 86.365 25.365 86.535 26.165 ;
        RECT 85.525 25.195 86.535 25.365 ;
        RECT 86.705 26.155 87.635 26.325 ;
        RECT 87.805 26.155 88.060 26.725 ;
        RECT 86.705 25.025 86.875 26.155 ;
        RECT 87.465 25.985 87.635 26.155 ;
        RECT 85.750 24.855 86.875 25.025 ;
        RECT 87.045 25.655 87.240 25.985 ;
        RECT 87.465 25.655 87.720 25.985 ;
        RECT 87.045 24.685 87.215 25.655 ;
        RECT 87.890 25.485 88.060 26.155 ;
        RECT 85.185 24.515 87.215 24.685 ;
        RECT 87.385 24.345 87.555 25.485 ;
        RECT 87.725 24.515 88.060 25.485 ;
        RECT 84.010 24.175 88.150 24.345 ;
        RECT 75.200 23.285 75.370 23.305 ;
        RECT 76.620 23.305 77.630 23.475 ;
        RECT 64.660 22.625 72.020 22.795 ;
        RECT 74.700 22.775 75.030 23.135 ;
        RECT 75.200 22.945 76.285 23.285 ;
        RECT 76.620 22.945 76.790 23.305 ;
        RECT 76.960 22.775 77.290 23.135 ;
        RECT 77.460 22.945 77.630 23.305 ;
        RECT 78.335 23.305 79.410 23.475 ;
        RECT 80.265 23.465 80.855 23.785 ;
        RECT 80.265 23.345 80.435 23.465 ;
        RECT 77.800 22.775 78.130 23.155 ;
        RECT 78.335 22.945 78.570 23.305 ;
        RECT 78.740 22.775 79.070 23.135 ;
        RECT 79.240 22.945 79.410 23.305 ;
        RECT 79.660 22.945 80.435 23.345 ;
        RECT 80.605 22.775 80.855 23.260 ;
        RECT 81.025 22.945 81.285 23.925 ;
        RECT 74.010 22.605 81.370 22.775 ;
        RECT 30.410 16.615 31.790 16.785 ;
        RECT 30.740 15.815 31.070 16.445 ;
        RECT 30.740 15.215 30.970 15.815 ;
        RECT 31.240 15.795 31.470 16.615 ;
        RECT 31.140 15.385 31.470 15.625 ;
        RECT 30.740 14.235 31.070 15.215 ;
        RECT 31.240 14.065 31.450 15.205 ;
        RECT 30.410 13.895 31.790 14.065 ;
        RECT 9.030 11.355 16.390 11.525 ;
        RECT 9.150 10.630 9.550 11.185 ;
        RECT 9.795 10.995 10.125 11.355 ;
        RECT 10.295 10.935 11.305 11.185 ;
        RECT 10.295 10.825 10.465 10.935 ;
        RECT 11.135 10.845 11.305 10.935 ;
        RECT 9.725 10.655 10.465 10.825 ;
        RECT 11.640 10.825 11.810 11.185 ;
        RECT 11.980 10.995 12.310 11.355 ;
        RECT 12.480 10.825 12.650 11.185 ;
        RECT 12.820 10.950 13.150 11.355 ;
        RECT 9.150 9.955 9.480 10.630 ;
        RECT 9.725 10.445 9.895 10.655 ;
        RECT 9.650 10.115 9.895 10.445 ;
        RECT 10.930 10.485 11.425 10.675 ;
        RECT 11.640 10.655 12.650 10.825 ;
        RECT 13.420 10.825 13.590 11.185 ;
        RECT 13.760 10.995 14.090 11.355 ;
        RECT 14.260 10.825 14.430 11.185 ;
        RECT 13.420 10.655 14.430 10.825 ;
        RECT 14.680 10.805 15.280 11.185 ;
        RECT 15.545 10.975 15.875 11.355 ;
        RECT 18.380 11.335 25.740 11.505 ;
        RECT 14.680 10.635 15.875 10.805 ;
        RECT 14.680 10.505 14.920 10.635 ;
        RECT 10.065 10.165 10.505 10.405 ;
        RECT 10.930 10.315 11.595 10.485 ;
        RECT 11.765 10.165 12.140 10.485 ;
        RECT 12.435 10.190 13.600 10.475 ;
        RECT 15.705 10.445 15.875 10.635 ;
        RECT 16.045 10.610 16.305 11.185 ;
        RECT 9.150 8.975 9.550 9.955 ;
        RECT 9.725 9.505 9.895 10.115 ;
        RECT 10.335 9.675 10.755 9.995 ;
        RECT 12.435 9.925 12.605 10.190 ;
        RECT 10.985 9.755 12.605 9.925 ;
        RECT 9.725 9.335 10.390 9.505 ;
        RECT 10.985 9.485 11.235 9.755 ;
        RECT 12.830 9.675 13.190 10.005 ;
        RECT 13.430 9.845 13.600 10.190 ;
        RECT 13.770 10.080 14.160 10.410 ;
        RECT 14.350 10.165 14.720 10.335 ;
        RECT 15.150 10.165 15.480 10.445 ;
        RECT 14.350 9.845 14.520 10.165 ;
        RECT 15.310 10.115 15.480 10.165 ;
        RECT 15.705 10.115 15.960 10.445 ;
        RECT 13.430 9.675 14.520 9.845 ;
        RECT 14.690 9.560 15.090 9.995 ;
        RECT 15.705 9.815 15.875 10.115 ;
        RECT 16.130 9.955 16.305 10.610 ;
        RECT 10.220 9.315 10.390 9.335 ;
        RECT 11.640 9.335 12.650 9.505 ;
        RECT 9.720 8.805 10.050 9.165 ;
        RECT 10.220 8.975 11.305 9.315 ;
        RECT 11.640 8.975 11.810 9.335 ;
        RECT 11.980 8.805 12.310 9.165 ;
        RECT 12.480 8.975 12.650 9.335 ;
        RECT 13.355 9.335 14.430 9.505 ;
        RECT 15.285 9.495 15.875 9.815 ;
        RECT 15.285 9.375 15.455 9.495 ;
        RECT 12.820 8.805 13.150 9.185 ;
        RECT 13.355 8.975 13.590 9.335 ;
        RECT 13.760 8.805 14.090 9.165 ;
        RECT 14.260 8.975 14.430 9.335 ;
        RECT 14.680 8.975 15.455 9.375 ;
        RECT 15.625 8.805 15.875 9.290 ;
        RECT 16.045 8.975 16.305 9.955 ;
        RECT 18.500 10.610 18.900 11.165 ;
        RECT 19.145 10.975 19.475 11.335 ;
        RECT 19.645 10.915 20.655 11.165 ;
        RECT 19.645 10.805 19.815 10.915 ;
        RECT 20.485 10.825 20.655 10.915 ;
        RECT 19.075 10.635 19.815 10.805 ;
        RECT 20.990 10.805 21.160 11.165 ;
        RECT 21.330 10.975 21.660 11.335 ;
        RECT 21.830 10.805 22.000 11.165 ;
        RECT 22.170 10.930 22.500 11.335 ;
        RECT 18.500 9.935 18.830 10.610 ;
        RECT 19.075 10.425 19.245 10.635 ;
        RECT 19.000 10.095 19.245 10.425 ;
        RECT 20.280 10.465 20.775 10.655 ;
        RECT 20.990 10.635 22.000 10.805 ;
        RECT 22.770 10.805 22.940 11.165 ;
        RECT 23.110 10.975 23.440 11.335 ;
        RECT 23.610 10.805 23.780 11.165 ;
        RECT 22.770 10.635 23.780 10.805 ;
        RECT 24.030 10.785 24.630 11.165 ;
        RECT 24.895 10.955 25.225 11.335 ;
        RECT 27.460 11.315 34.820 11.485 ;
        RECT 24.030 10.615 25.225 10.785 ;
        RECT 24.030 10.485 24.270 10.615 ;
        RECT 19.415 10.145 19.855 10.385 ;
        RECT 20.280 10.295 20.945 10.465 ;
        RECT 21.115 10.145 21.490 10.465 ;
        RECT 21.785 10.170 22.950 10.455 ;
        RECT 25.055 10.425 25.225 10.615 ;
        RECT 25.395 10.590 25.655 11.165 ;
        RECT 18.500 8.955 18.900 9.935 ;
        RECT 19.075 9.485 19.245 10.095 ;
        RECT 19.685 9.655 20.105 9.975 ;
        RECT 21.785 9.905 21.955 10.170 ;
        RECT 20.335 9.735 21.955 9.905 ;
        RECT 19.075 9.315 19.740 9.485 ;
        RECT 20.335 9.465 20.585 9.735 ;
        RECT 22.180 9.655 22.540 9.985 ;
        RECT 22.780 9.825 22.950 10.170 ;
        RECT 23.120 10.060 23.510 10.390 ;
        RECT 23.700 10.145 24.070 10.315 ;
        RECT 24.500 10.145 24.830 10.425 ;
        RECT 23.700 9.825 23.870 10.145 ;
        RECT 24.660 10.095 24.830 10.145 ;
        RECT 25.055 10.095 25.310 10.425 ;
        RECT 22.780 9.655 23.870 9.825 ;
        RECT 24.040 9.540 24.440 9.975 ;
        RECT 25.055 9.795 25.225 10.095 ;
        RECT 25.480 9.935 25.655 10.590 ;
        RECT 19.570 9.295 19.740 9.315 ;
        RECT 20.990 9.315 22.000 9.485 ;
        RECT 9.030 8.635 16.390 8.805 ;
        RECT 19.070 8.785 19.400 9.145 ;
        RECT 19.570 8.955 20.655 9.295 ;
        RECT 20.990 8.955 21.160 9.315 ;
        RECT 21.330 8.785 21.660 9.145 ;
        RECT 21.830 8.955 22.000 9.315 ;
        RECT 22.705 9.315 23.780 9.485 ;
        RECT 24.635 9.475 25.225 9.795 ;
        RECT 24.635 9.355 24.805 9.475 ;
        RECT 22.170 8.785 22.500 9.165 ;
        RECT 22.705 8.955 22.940 9.315 ;
        RECT 23.110 8.785 23.440 9.145 ;
        RECT 23.610 8.955 23.780 9.315 ;
        RECT 24.030 8.955 24.805 9.355 ;
        RECT 24.975 8.785 25.225 9.270 ;
        RECT 25.395 8.955 25.655 9.935 ;
        RECT 27.580 10.590 27.980 11.145 ;
        RECT 28.225 10.955 28.555 11.315 ;
        RECT 28.725 10.895 29.735 11.145 ;
        RECT 28.725 10.785 28.895 10.895 ;
        RECT 29.565 10.805 29.735 10.895 ;
        RECT 28.155 10.615 28.895 10.785 ;
        RECT 30.070 10.785 30.240 11.145 ;
        RECT 30.410 10.955 30.740 11.315 ;
        RECT 30.910 10.785 31.080 11.145 ;
        RECT 31.250 10.910 31.580 11.315 ;
        RECT 27.580 9.915 27.910 10.590 ;
        RECT 28.155 10.405 28.325 10.615 ;
        RECT 28.080 10.075 28.325 10.405 ;
        RECT 29.360 10.445 29.855 10.635 ;
        RECT 30.070 10.615 31.080 10.785 ;
        RECT 31.850 10.785 32.020 11.145 ;
        RECT 32.190 10.955 32.520 11.315 ;
        RECT 32.690 10.785 32.860 11.145 ;
        RECT 31.850 10.615 32.860 10.785 ;
        RECT 33.110 10.765 33.710 11.145 ;
        RECT 33.975 10.935 34.305 11.315 ;
        RECT 36.810 11.295 44.170 11.465 ;
        RECT 33.110 10.595 34.305 10.765 ;
        RECT 33.110 10.465 33.350 10.595 ;
        RECT 28.495 10.125 28.935 10.365 ;
        RECT 29.360 10.275 30.025 10.445 ;
        RECT 30.195 10.125 30.570 10.445 ;
        RECT 30.865 10.150 32.030 10.435 ;
        RECT 34.135 10.405 34.305 10.595 ;
        RECT 34.475 10.570 34.735 11.145 ;
        RECT 27.580 8.935 27.980 9.915 ;
        RECT 28.155 9.465 28.325 10.075 ;
        RECT 28.765 9.635 29.185 9.955 ;
        RECT 30.865 9.885 31.035 10.150 ;
        RECT 29.415 9.715 31.035 9.885 ;
        RECT 28.155 9.295 28.820 9.465 ;
        RECT 29.415 9.445 29.665 9.715 ;
        RECT 31.260 9.635 31.620 9.965 ;
        RECT 31.860 9.805 32.030 10.150 ;
        RECT 32.200 10.040 32.590 10.370 ;
        RECT 32.780 10.125 33.150 10.295 ;
        RECT 33.580 10.125 33.910 10.405 ;
        RECT 32.780 9.805 32.950 10.125 ;
        RECT 33.740 10.075 33.910 10.125 ;
        RECT 34.135 10.075 34.390 10.405 ;
        RECT 31.860 9.635 32.950 9.805 ;
        RECT 33.120 9.520 33.520 9.955 ;
        RECT 34.135 9.775 34.305 10.075 ;
        RECT 34.560 9.915 34.735 10.570 ;
        RECT 28.650 9.275 28.820 9.295 ;
        RECT 30.070 9.295 31.080 9.465 ;
        RECT 18.380 8.615 25.740 8.785 ;
        RECT 28.150 8.765 28.480 9.125 ;
        RECT 28.650 8.935 29.735 9.275 ;
        RECT 30.070 8.935 30.240 9.295 ;
        RECT 30.410 8.765 30.740 9.125 ;
        RECT 30.910 8.935 31.080 9.295 ;
        RECT 31.785 9.295 32.860 9.465 ;
        RECT 33.715 9.455 34.305 9.775 ;
        RECT 33.715 9.335 33.885 9.455 ;
        RECT 31.250 8.765 31.580 9.145 ;
        RECT 31.785 8.935 32.020 9.295 ;
        RECT 32.190 8.765 32.520 9.125 ;
        RECT 32.690 8.935 32.860 9.295 ;
        RECT 33.110 8.935 33.885 9.335 ;
        RECT 34.055 8.765 34.305 9.250 ;
        RECT 34.475 8.935 34.735 9.915 ;
        RECT 36.930 10.570 37.330 11.125 ;
        RECT 37.575 10.935 37.905 11.295 ;
        RECT 38.075 10.875 39.085 11.125 ;
        RECT 38.075 10.765 38.245 10.875 ;
        RECT 38.915 10.785 39.085 10.875 ;
        RECT 37.505 10.595 38.245 10.765 ;
        RECT 39.420 10.765 39.590 11.125 ;
        RECT 39.760 10.935 40.090 11.295 ;
        RECT 40.260 10.765 40.430 11.125 ;
        RECT 40.600 10.890 40.930 11.295 ;
        RECT 36.930 9.895 37.260 10.570 ;
        RECT 37.505 10.385 37.675 10.595 ;
        RECT 37.430 10.055 37.675 10.385 ;
        RECT 38.710 10.425 39.205 10.615 ;
        RECT 39.420 10.595 40.430 10.765 ;
        RECT 41.200 10.765 41.370 11.125 ;
        RECT 41.540 10.935 41.870 11.295 ;
        RECT 42.040 10.765 42.210 11.125 ;
        RECT 41.200 10.595 42.210 10.765 ;
        RECT 42.460 10.745 43.060 11.125 ;
        RECT 43.325 10.915 43.655 11.295 ;
        RECT 45.880 11.285 53.240 11.455 ;
        RECT 42.460 10.575 43.655 10.745 ;
        RECT 42.460 10.445 42.700 10.575 ;
        RECT 37.845 10.105 38.285 10.345 ;
        RECT 38.710 10.255 39.375 10.425 ;
        RECT 39.545 10.105 39.920 10.425 ;
        RECT 40.215 10.130 41.380 10.415 ;
        RECT 43.485 10.385 43.655 10.575 ;
        RECT 43.825 10.550 44.085 11.125 ;
        RECT 36.930 8.915 37.330 9.895 ;
        RECT 37.505 9.445 37.675 10.055 ;
        RECT 38.115 9.615 38.535 9.935 ;
        RECT 40.215 9.865 40.385 10.130 ;
        RECT 38.765 9.695 40.385 9.865 ;
        RECT 37.505 9.275 38.170 9.445 ;
        RECT 38.765 9.425 39.015 9.695 ;
        RECT 40.610 9.615 40.970 9.945 ;
        RECT 41.210 9.785 41.380 10.130 ;
        RECT 41.550 10.020 41.940 10.350 ;
        RECT 42.130 10.105 42.500 10.275 ;
        RECT 42.930 10.105 43.260 10.385 ;
        RECT 42.130 9.785 42.300 10.105 ;
        RECT 43.090 10.055 43.260 10.105 ;
        RECT 43.485 10.055 43.740 10.385 ;
        RECT 41.210 9.615 42.300 9.785 ;
        RECT 42.470 9.500 42.870 9.935 ;
        RECT 43.485 9.755 43.655 10.055 ;
        RECT 43.910 9.895 44.085 10.550 ;
        RECT 38.000 9.255 38.170 9.275 ;
        RECT 39.420 9.275 40.430 9.445 ;
        RECT 27.460 8.595 34.820 8.765 ;
        RECT 37.500 8.745 37.830 9.105 ;
        RECT 38.000 8.915 39.085 9.255 ;
        RECT 39.420 8.915 39.590 9.275 ;
        RECT 39.760 8.745 40.090 9.105 ;
        RECT 40.260 8.915 40.430 9.275 ;
        RECT 41.135 9.275 42.210 9.445 ;
        RECT 43.065 9.435 43.655 9.755 ;
        RECT 43.065 9.315 43.235 9.435 ;
        RECT 40.600 8.745 40.930 9.125 ;
        RECT 41.135 8.915 41.370 9.275 ;
        RECT 41.540 8.745 41.870 9.105 ;
        RECT 42.040 8.915 42.210 9.275 ;
        RECT 42.460 8.915 43.235 9.315 ;
        RECT 43.405 8.745 43.655 9.230 ;
        RECT 43.825 8.915 44.085 9.895 ;
        RECT 46.000 10.560 46.400 11.115 ;
        RECT 46.645 10.925 46.975 11.285 ;
        RECT 47.145 10.865 48.155 11.115 ;
        RECT 47.145 10.755 47.315 10.865 ;
        RECT 47.985 10.775 48.155 10.865 ;
        RECT 46.575 10.585 47.315 10.755 ;
        RECT 48.490 10.755 48.660 11.115 ;
        RECT 48.830 10.925 49.160 11.285 ;
        RECT 49.330 10.755 49.500 11.115 ;
        RECT 49.670 10.880 50.000 11.285 ;
        RECT 46.000 9.885 46.330 10.560 ;
        RECT 46.575 10.375 46.745 10.585 ;
        RECT 46.500 10.045 46.745 10.375 ;
        RECT 47.780 10.415 48.275 10.605 ;
        RECT 48.490 10.585 49.500 10.755 ;
        RECT 50.270 10.755 50.440 11.115 ;
        RECT 50.610 10.925 50.940 11.285 ;
        RECT 51.110 10.755 51.280 11.115 ;
        RECT 50.270 10.585 51.280 10.755 ;
        RECT 51.530 10.735 52.130 11.115 ;
        RECT 52.395 10.905 52.725 11.285 ;
        RECT 55.230 11.265 62.590 11.435 ;
        RECT 51.530 10.565 52.725 10.735 ;
        RECT 51.530 10.435 51.770 10.565 ;
        RECT 46.915 10.095 47.355 10.335 ;
        RECT 47.780 10.245 48.445 10.415 ;
        RECT 48.615 10.095 48.990 10.415 ;
        RECT 49.285 10.120 50.450 10.405 ;
        RECT 52.555 10.375 52.725 10.565 ;
        RECT 52.895 10.540 53.155 11.115 ;
        RECT 46.000 8.905 46.400 9.885 ;
        RECT 46.575 9.435 46.745 10.045 ;
        RECT 47.185 9.605 47.605 9.925 ;
        RECT 49.285 9.855 49.455 10.120 ;
        RECT 47.835 9.685 49.455 9.855 ;
        RECT 46.575 9.265 47.240 9.435 ;
        RECT 47.835 9.415 48.085 9.685 ;
        RECT 49.680 9.605 50.040 9.935 ;
        RECT 50.280 9.775 50.450 10.120 ;
        RECT 50.620 10.010 51.010 10.340 ;
        RECT 51.200 10.095 51.570 10.265 ;
        RECT 52.000 10.095 52.330 10.375 ;
        RECT 51.200 9.775 51.370 10.095 ;
        RECT 52.160 10.045 52.330 10.095 ;
        RECT 52.555 10.045 52.810 10.375 ;
        RECT 50.280 9.605 51.370 9.775 ;
        RECT 51.540 9.490 51.940 9.925 ;
        RECT 52.555 9.745 52.725 10.045 ;
        RECT 52.980 9.885 53.155 10.540 ;
        RECT 47.070 9.245 47.240 9.265 ;
        RECT 48.490 9.265 49.500 9.435 ;
        RECT 36.810 8.575 44.170 8.745 ;
        RECT 46.570 8.735 46.900 9.095 ;
        RECT 47.070 8.905 48.155 9.245 ;
        RECT 48.490 8.905 48.660 9.265 ;
        RECT 48.830 8.735 49.160 9.095 ;
        RECT 49.330 8.905 49.500 9.265 ;
        RECT 50.205 9.265 51.280 9.435 ;
        RECT 52.135 9.425 52.725 9.745 ;
        RECT 52.135 9.305 52.305 9.425 ;
        RECT 49.670 8.735 50.000 9.115 ;
        RECT 50.205 8.905 50.440 9.265 ;
        RECT 50.610 8.735 50.940 9.095 ;
        RECT 51.110 8.905 51.280 9.265 ;
        RECT 51.530 8.905 52.305 9.305 ;
        RECT 52.475 8.735 52.725 9.220 ;
        RECT 52.895 8.905 53.155 9.885 ;
        RECT 55.350 10.540 55.750 11.095 ;
        RECT 55.995 10.905 56.325 11.265 ;
        RECT 56.495 10.845 57.505 11.095 ;
        RECT 56.495 10.735 56.665 10.845 ;
        RECT 57.335 10.755 57.505 10.845 ;
        RECT 55.925 10.565 56.665 10.735 ;
        RECT 57.840 10.735 58.010 11.095 ;
        RECT 58.180 10.905 58.510 11.265 ;
        RECT 58.680 10.735 58.850 11.095 ;
        RECT 59.020 10.860 59.350 11.265 ;
        RECT 55.350 9.865 55.680 10.540 ;
        RECT 55.925 10.355 56.095 10.565 ;
        RECT 55.850 10.025 56.095 10.355 ;
        RECT 57.130 10.395 57.625 10.585 ;
        RECT 57.840 10.565 58.850 10.735 ;
        RECT 59.620 10.735 59.790 11.095 ;
        RECT 59.960 10.905 60.290 11.265 ;
        RECT 60.460 10.735 60.630 11.095 ;
        RECT 59.620 10.565 60.630 10.735 ;
        RECT 60.880 10.715 61.480 11.095 ;
        RECT 61.745 10.885 62.075 11.265 ;
        RECT 64.310 11.245 71.670 11.415 ;
        RECT 60.880 10.545 62.075 10.715 ;
        RECT 60.880 10.415 61.120 10.545 ;
        RECT 56.265 10.075 56.705 10.315 ;
        RECT 57.130 10.225 57.795 10.395 ;
        RECT 57.965 10.075 58.340 10.395 ;
        RECT 58.635 10.100 59.800 10.385 ;
        RECT 61.905 10.355 62.075 10.545 ;
        RECT 62.245 10.520 62.505 11.095 ;
        RECT 55.350 8.885 55.750 9.865 ;
        RECT 55.925 9.415 56.095 10.025 ;
        RECT 56.535 9.585 56.955 9.905 ;
        RECT 58.635 9.835 58.805 10.100 ;
        RECT 57.185 9.665 58.805 9.835 ;
        RECT 55.925 9.245 56.590 9.415 ;
        RECT 57.185 9.395 57.435 9.665 ;
        RECT 59.030 9.585 59.390 9.915 ;
        RECT 59.630 9.755 59.800 10.100 ;
        RECT 59.970 9.990 60.360 10.320 ;
        RECT 60.550 10.075 60.920 10.245 ;
        RECT 61.350 10.075 61.680 10.355 ;
        RECT 60.550 9.755 60.720 10.075 ;
        RECT 61.510 10.025 61.680 10.075 ;
        RECT 61.905 10.025 62.160 10.355 ;
        RECT 59.630 9.585 60.720 9.755 ;
        RECT 60.890 9.470 61.290 9.905 ;
        RECT 61.905 9.725 62.075 10.025 ;
        RECT 62.330 9.865 62.505 10.520 ;
        RECT 56.420 9.225 56.590 9.245 ;
        RECT 57.840 9.245 58.850 9.415 ;
        RECT 45.880 8.565 53.240 8.735 ;
        RECT 55.920 8.715 56.250 9.075 ;
        RECT 56.420 8.885 57.505 9.225 ;
        RECT 57.840 8.885 58.010 9.245 ;
        RECT 58.180 8.715 58.510 9.075 ;
        RECT 58.680 8.885 58.850 9.245 ;
        RECT 59.555 9.245 60.630 9.415 ;
        RECT 61.485 9.405 62.075 9.725 ;
        RECT 61.485 9.285 61.655 9.405 ;
        RECT 59.020 8.715 59.350 9.095 ;
        RECT 59.555 8.885 59.790 9.245 ;
        RECT 59.960 8.715 60.290 9.075 ;
        RECT 60.460 8.885 60.630 9.245 ;
        RECT 60.880 8.885 61.655 9.285 ;
        RECT 61.825 8.715 62.075 9.200 ;
        RECT 62.245 8.885 62.505 9.865 ;
        RECT 64.430 10.520 64.830 11.075 ;
        RECT 65.075 10.885 65.405 11.245 ;
        RECT 65.575 10.825 66.585 11.075 ;
        RECT 65.575 10.715 65.745 10.825 ;
        RECT 66.415 10.735 66.585 10.825 ;
        RECT 65.005 10.545 65.745 10.715 ;
        RECT 66.920 10.715 67.090 11.075 ;
        RECT 67.260 10.885 67.590 11.245 ;
        RECT 67.760 10.715 67.930 11.075 ;
        RECT 68.100 10.840 68.430 11.245 ;
        RECT 64.430 9.845 64.760 10.520 ;
        RECT 65.005 10.335 65.175 10.545 ;
        RECT 64.930 10.005 65.175 10.335 ;
        RECT 66.210 10.375 66.705 10.565 ;
        RECT 66.920 10.545 67.930 10.715 ;
        RECT 68.700 10.715 68.870 11.075 ;
        RECT 69.040 10.885 69.370 11.245 ;
        RECT 69.540 10.715 69.710 11.075 ;
        RECT 68.700 10.545 69.710 10.715 ;
        RECT 69.960 10.695 70.560 11.075 ;
        RECT 70.825 10.865 71.155 11.245 ;
        RECT 73.660 11.225 81.020 11.395 ;
        RECT 69.960 10.525 71.155 10.695 ;
        RECT 69.960 10.395 70.200 10.525 ;
        RECT 65.345 10.055 65.785 10.295 ;
        RECT 66.210 10.205 66.875 10.375 ;
        RECT 67.045 10.055 67.420 10.375 ;
        RECT 67.715 10.080 68.880 10.365 ;
        RECT 70.985 10.335 71.155 10.525 ;
        RECT 71.325 10.500 71.585 11.075 ;
        RECT 64.430 8.865 64.830 9.845 ;
        RECT 65.005 9.395 65.175 10.005 ;
        RECT 65.615 9.565 66.035 9.885 ;
        RECT 67.715 9.815 67.885 10.080 ;
        RECT 66.265 9.645 67.885 9.815 ;
        RECT 65.005 9.225 65.670 9.395 ;
        RECT 66.265 9.375 66.515 9.645 ;
        RECT 68.110 9.565 68.470 9.895 ;
        RECT 68.710 9.735 68.880 10.080 ;
        RECT 69.050 9.970 69.440 10.300 ;
        RECT 69.630 10.055 70.000 10.225 ;
        RECT 70.430 10.055 70.760 10.335 ;
        RECT 69.630 9.735 69.800 10.055 ;
        RECT 70.590 10.005 70.760 10.055 ;
        RECT 70.985 10.005 71.240 10.335 ;
        RECT 68.710 9.565 69.800 9.735 ;
        RECT 69.970 9.450 70.370 9.885 ;
        RECT 70.985 9.705 71.155 10.005 ;
        RECT 71.410 9.845 71.585 10.500 ;
        RECT 65.500 9.205 65.670 9.225 ;
        RECT 66.920 9.225 67.930 9.395 ;
        RECT 55.230 8.545 62.590 8.715 ;
        RECT 65.000 8.695 65.330 9.055 ;
        RECT 65.500 8.865 66.585 9.205 ;
        RECT 66.920 8.865 67.090 9.225 ;
        RECT 67.260 8.695 67.590 9.055 ;
        RECT 67.760 8.865 67.930 9.225 ;
        RECT 68.635 9.225 69.710 9.395 ;
        RECT 70.565 9.385 71.155 9.705 ;
        RECT 70.565 9.265 70.735 9.385 ;
        RECT 68.100 8.695 68.430 9.075 ;
        RECT 68.635 8.865 68.870 9.225 ;
        RECT 69.040 8.695 69.370 9.055 ;
        RECT 69.540 8.865 69.710 9.225 ;
        RECT 69.960 8.865 70.735 9.265 ;
        RECT 70.905 8.695 71.155 9.180 ;
        RECT 71.325 8.865 71.585 9.845 ;
        RECT 73.780 10.500 74.180 11.055 ;
        RECT 74.425 10.865 74.755 11.225 ;
        RECT 74.925 10.805 75.935 11.055 ;
        RECT 74.925 10.695 75.095 10.805 ;
        RECT 75.765 10.715 75.935 10.805 ;
        RECT 74.355 10.525 75.095 10.695 ;
        RECT 76.270 10.695 76.440 11.055 ;
        RECT 76.610 10.865 76.940 11.225 ;
        RECT 77.110 10.695 77.280 11.055 ;
        RECT 77.450 10.820 77.780 11.225 ;
        RECT 73.780 9.825 74.110 10.500 ;
        RECT 74.355 10.315 74.525 10.525 ;
        RECT 74.280 9.985 74.525 10.315 ;
        RECT 75.560 10.355 76.055 10.545 ;
        RECT 76.270 10.525 77.280 10.695 ;
        RECT 78.050 10.695 78.220 11.055 ;
        RECT 78.390 10.865 78.720 11.225 ;
        RECT 78.890 10.695 79.060 11.055 ;
        RECT 78.050 10.525 79.060 10.695 ;
        RECT 79.310 10.675 79.910 11.055 ;
        RECT 80.175 10.845 80.505 11.225 ;
        RECT 79.310 10.505 80.505 10.675 ;
        RECT 79.310 10.375 79.550 10.505 ;
        RECT 74.695 10.035 75.135 10.275 ;
        RECT 75.560 10.185 76.225 10.355 ;
        RECT 76.395 10.035 76.770 10.355 ;
        RECT 77.065 10.060 78.230 10.345 ;
        RECT 80.335 10.315 80.505 10.505 ;
        RECT 80.675 10.480 80.935 11.055 ;
        RECT 73.780 8.845 74.180 9.825 ;
        RECT 74.355 9.375 74.525 9.985 ;
        RECT 74.965 9.545 75.385 9.865 ;
        RECT 77.065 9.795 77.235 10.060 ;
        RECT 75.615 9.625 77.235 9.795 ;
        RECT 74.355 9.205 75.020 9.375 ;
        RECT 75.615 9.355 75.865 9.625 ;
        RECT 77.460 9.545 77.820 9.875 ;
        RECT 78.060 9.715 78.230 10.060 ;
        RECT 78.400 9.950 78.790 10.280 ;
        RECT 78.980 10.035 79.350 10.205 ;
        RECT 79.780 10.035 80.110 10.315 ;
        RECT 78.980 9.715 79.150 10.035 ;
        RECT 79.940 9.985 80.110 10.035 ;
        RECT 80.335 9.985 80.590 10.315 ;
        RECT 78.060 9.545 79.150 9.715 ;
        RECT 79.320 9.430 79.720 9.865 ;
        RECT 80.335 9.685 80.505 9.985 ;
        RECT 80.760 9.825 80.935 10.480 ;
        RECT 74.850 9.185 75.020 9.205 ;
        RECT 76.270 9.205 77.280 9.375 ;
        RECT 64.310 8.525 71.670 8.695 ;
        RECT 74.350 8.675 74.680 9.035 ;
        RECT 74.850 8.845 75.935 9.185 ;
        RECT 76.270 8.845 76.440 9.205 ;
        RECT 76.610 8.675 76.940 9.035 ;
        RECT 77.110 8.845 77.280 9.205 ;
        RECT 77.985 9.205 79.060 9.375 ;
        RECT 79.915 9.365 80.505 9.685 ;
        RECT 79.915 9.245 80.085 9.365 ;
        RECT 77.450 8.675 77.780 9.055 ;
        RECT 77.985 8.845 78.220 9.205 ;
        RECT 78.390 8.675 78.720 9.035 ;
        RECT 78.890 8.845 79.060 9.205 ;
        RECT 79.310 8.845 80.085 9.245 ;
        RECT 80.255 8.675 80.505 9.160 ;
        RECT 80.675 8.845 80.935 9.825 ;
        RECT 73.660 8.505 81.020 8.675 ;
      LAYER met1 ;
        RECT 47.150 88.730 48.530 89.210 ;
        RECT 33.015 87.485 47.695 87.935 ;
        RECT 47.865 87.485 68.665 87.935 ;
        RECT 47.150 86.010 48.530 86.490 ;
        RECT 45.225 85.270 57.410 85.275 ;
        RECT 45.180 84.885 57.410 85.270 ;
        RECT 45.180 83.500 45.620 84.885 ;
        RECT 22.340 82.690 25.560 83.170 ;
        RECT 22.730 81.190 23.030 82.690 ;
        RECT 29.730 82.020 30.740 82.190 ;
        RECT 25.160 81.690 31.295 82.020 ;
        RECT 29.730 81.560 30.740 81.690 ;
        RECT 23.180 81.260 23.730 81.540 ;
        RECT 23.350 80.450 23.505 81.260 ;
        RECT 22.340 79.970 25.560 80.450 ;
        RECT 22.830 78.970 25.130 79.450 ;
        RECT 22.870 77.570 23.250 77.930 ;
        RECT 23.880 77.850 24.150 78.970 ;
        RECT 30.965 78.165 31.295 81.690 ;
        RECT 33.040 78.420 36.260 78.900 ;
        RECT 22.920 76.730 23.190 77.570 ;
        RECT 23.830 77.540 24.170 77.850 ;
        RECT 30.965 77.835 35.235 78.165 ;
        RECT 33.955 77.820 34.285 77.835 ;
        RECT 24.790 77.180 25.220 77.550 ;
        RECT 25.970 77.290 34.280 77.580 ;
        RECT 25.970 77.260 34.285 77.290 ;
        RECT 23.830 76.730 24.170 76.740 ;
        RECT 22.830 76.250 25.130 76.730 ;
        RECT 22.390 74.870 25.610 75.350 ;
        RECT 22.780 73.370 23.080 74.870 ;
        RECT 25.970 74.710 26.290 77.260 ;
        RECT 32.890 76.710 33.410 77.120 ;
        RECT 33.955 76.950 34.285 77.260 ;
        RECT 34.450 76.570 34.740 76.650 ;
        RECT 28.750 75.920 31.050 76.400 ;
        RECT 31.740 76.350 34.740 76.570 ;
        RECT 31.750 75.780 32.150 76.350 ;
        RECT 34.450 76.320 34.740 76.350 ;
        RECT 34.905 76.330 35.235 77.835 ;
        RECT 35.890 77.200 36.170 77.220 ;
        RECT 35.890 76.950 37.000 77.200 ;
        RECT 35.890 76.930 36.170 76.950 ;
        RECT 25.200 74.390 26.290 74.710 ;
        RECT 26.450 75.400 30.100 75.660 ;
        RECT 30.520 75.490 32.150 75.780 ;
        RECT 33.040 75.700 36.260 76.180 ;
        RECT 23.230 73.440 23.780 73.720 ;
        RECT 23.400 72.630 23.555 73.440 ;
        RECT 22.390 72.150 25.610 72.630 ;
        RECT 22.880 71.150 25.180 71.630 ;
        RECT 22.920 69.750 23.300 70.120 ;
        RECT 23.940 70.030 24.170 71.150 ;
        RECT 22.960 68.910 23.230 69.750 ;
        RECT 23.880 69.720 24.220 70.030 ;
        RECT 24.830 69.100 25.690 69.570 ;
        RECT 22.880 68.430 25.180 68.910 ;
        RECT 22.350 66.530 25.570 67.010 ;
        RECT 26.450 66.830 26.710 75.400 ;
        RECT 29.840 74.780 30.100 75.400 ;
        RECT 28.850 74.755 29.530 74.760 ;
        RECT 27.810 74.390 29.530 74.755 ;
        RECT 29.700 74.450 30.100 74.780 ;
        RECT 27.810 74.365 29.225 74.390 ;
        RECT 27.810 69.855 28.200 74.365 ;
        RECT 28.750 73.200 31.050 73.680 ;
        RECT 29.120 71.090 32.340 71.570 ;
        RECT 36.735 70.885 36.985 76.950 ;
        RECT 38.210 71.010 40.970 71.490 ;
        RECT 36.735 70.860 36.990 70.885 ;
        RECT 36.735 70.625 39.970 70.860 ;
        RECT 36.950 70.620 39.970 70.625 ;
        RECT 45.180 70.480 45.630 83.500 ;
        RECT 47.150 82.610 50.370 83.090 ;
        RECT 47.540 81.110 47.840 82.610 ;
        RECT 54.540 81.940 55.550 82.110 ;
        RECT 49.970 81.610 56.105 81.940 ;
        RECT 54.540 81.480 55.550 81.610 ;
        RECT 47.990 81.180 48.540 81.460 ;
        RECT 48.160 80.370 48.315 81.180 ;
        RECT 47.150 79.890 50.370 80.370 ;
        RECT 47.640 78.890 49.940 79.370 ;
        RECT 47.680 77.490 48.060 77.850 ;
        RECT 48.690 77.770 48.960 78.890 ;
        RECT 55.775 78.085 56.105 81.610 ;
        RECT 57.850 78.340 61.070 78.820 ;
        RECT 47.730 76.650 48.000 77.490 ;
        RECT 48.640 77.460 48.980 77.770 ;
        RECT 55.775 77.755 60.045 78.085 ;
        RECT 58.765 77.740 59.095 77.755 ;
        RECT 49.600 77.100 50.030 77.470 ;
        RECT 50.780 77.210 59.090 77.500 ;
        RECT 50.780 77.180 59.095 77.210 ;
        RECT 48.640 76.650 48.980 76.660 ;
        RECT 47.640 76.170 49.940 76.650 ;
        RECT 47.200 74.790 50.420 75.270 ;
        RECT 47.590 73.290 47.890 74.790 ;
        RECT 50.780 74.630 51.100 77.180 ;
        RECT 57.700 76.630 58.220 77.040 ;
        RECT 58.765 76.870 59.095 77.180 ;
        RECT 59.260 76.490 59.550 76.570 ;
        RECT 53.560 75.840 55.860 76.320 ;
        RECT 56.550 76.270 59.550 76.490 ;
        RECT 56.560 75.700 56.960 76.270 ;
        RECT 59.260 76.240 59.550 76.270 ;
        RECT 59.715 76.250 60.045 77.755 ;
        RECT 60.700 77.120 60.980 77.140 ;
        RECT 60.700 76.870 61.810 77.120 ;
        RECT 60.700 76.850 60.980 76.870 ;
        RECT 50.010 74.310 51.100 74.630 ;
        RECT 51.260 75.320 54.910 75.580 ;
        RECT 55.330 75.410 56.960 75.700 ;
        RECT 57.850 75.620 61.070 76.100 ;
        RECT 48.040 73.360 48.590 73.640 ;
        RECT 48.210 72.550 48.365 73.360 ;
        RECT 47.200 72.070 50.420 72.550 ;
        RECT 47.690 71.070 49.990 71.550 ;
        RECT 37.230 70.150 40.170 70.450 ;
        RECT 29.115 69.855 29.505 70.145 ;
        RECT 37.230 70.090 37.600 70.150 ;
        RECT 27.810 69.465 29.505 69.855 ;
        RECT 22.740 65.030 23.040 66.530 ;
        RECT 26.450 66.480 26.880 66.830 ;
        RECT 26.450 66.140 26.710 66.480 ;
        RECT 25.180 65.880 26.710 66.140 ;
        RECT 27.810 65.425 28.200 69.465 ;
        RECT 30.010 68.990 30.360 69.680 ;
        RECT 30.500 69.000 30.840 69.930 ;
        RECT 31.010 69.020 31.370 69.940 ;
        RECT 31.900 68.990 33.330 69.360 ;
        RECT 33.970 69.220 36.270 69.700 ;
        RECT 37.230 69.650 37.590 70.090 ;
        RECT 32.925 68.925 33.330 68.990 ;
        RECT 37.230 68.930 37.580 69.650 ;
        RECT 38.180 69.280 38.620 69.870 ;
        RECT 38.780 69.790 39.480 69.960 ;
        RECT 39.810 69.860 40.170 70.150 ;
        RECT 40.590 70.090 45.630 70.480 ;
        RECT 38.780 69.450 39.470 69.790 ;
        RECT 39.700 69.520 40.170 69.860 ;
        RECT 47.730 69.670 48.110 70.040 ;
        RECT 48.750 69.950 48.980 71.070 ;
        RECT 29.120 68.370 32.340 68.850 ;
        RECT 32.925 68.555 35.315 68.925 ;
        RECT 35.600 68.570 37.580 68.930 ;
        RECT 47.770 68.830 48.040 69.670 ;
        RECT 48.690 69.640 49.030 69.950 ;
        RECT 49.640 69.020 50.500 69.490 ;
        RECT 32.720 67.515 34.465 67.885 ;
        RECT 29.740 66.880 32.040 67.360 ;
        RECT 30.600 66.340 31.090 66.720 ;
        RECT 32.720 66.490 33.090 67.515 ;
        RECT 34.945 67.445 35.315 68.555 ;
        RECT 38.210 68.290 40.970 68.770 ;
        RECT 47.690 68.350 49.990 68.830 ;
        RECT 33.970 66.500 36.270 66.980 ;
        RECT 31.660 66.120 33.090 66.490 ;
        RECT 47.160 66.450 50.380 66.930 ;
        RECT 51.260 66.750 51.520 75.320 ;
        RECT 54.650 74.700 54.910 75.320 ;
        RECT 53.660 74.675 54.340 74.680 ;
        RECT 52.620 74.310 54.340 74.675 ;
        RECT 54.510 74.370 54.910 74.700 ;
        RECT 52.620 74.285 54.035 74.310 ;
        RECT 52.620 69.775 53.010 74.285 ;
        RECT 53.560 73.120 55.860 73.600 ;
        RECT 53.930 71.010 57.150 71.490 ;
        RECT 61.545 70.805 61.795 76.870 ;
        RECT 68.215 73.485 68.665 87.485 ;
        RECT 80.935 84.265 93.285 84.315 ;
        RECT 80.935 84.235 102.850 84.265 ;
        RECT 80.935 84.165 117.395 84.235 ;
        RECT 80.935 81.835 81.085 84.165 ;
        RECT 92.560 84.115 117.395 84.165 ;
        RECT 99.975 84.085 117.395 84.115 ;
        RECT 106.035 84.030 106.185 84.085 ;
        RECT 81.680 83.230 83.060 83.710 ;
        RECT 85.520 83.180 86.900 83.660 ;
        RECT 89.890 83.190 91.270 83.670 ;
        RECT 92.960 83.180 94.340 83.660 ;
        RECT 96.800 83.130 98.180 83.610 ;
        RECT 101.170 83.140 102.550 83.620 ;
        RECT 106.780 83.150 108.160 83.630 ;
        RECT 110.620 83.100 112.000 83.580 ;
        RECT 114.990 83.110 116.370 83.590 ;
        RECT 82.000 81.835 82.330 82.100 ;
        RECT 80.935 81.685 82.330 81.835 ;
        RECT 82.480 81.690 86.170 82.060 ;
        RECT 82.000 81.680 82.330 81.685 ;
        RECT 86.320 81.640 90.530 82.090 ;
        RECT 90.690 81.950 91.000 82.080 ;
        RECT 90.690 81.940 91.570 81.950 ;
        RECT 93.280 81.940 93.610 82.050 ;
        RECT 90.690 81.740 93.610 81.940 ;
        RECT 90.970 81.710 93.610 81.740 ;
        RECT 92.560 81.635 93.610 81.710 ;
        RECT 93.760 81.640 97.450 82.010 ;
        RECT 93.280 81.630 93.610 81.635 ;
        RECT 97.600 81.590 101.810 82.040 ;
        RECT 101.970 81.960 102.280 82.030 ;
        RECT 107.090 81.960 107.430 82.020 ;
        RECT 101.970 81.690 107.430 81.960 ;
        RECT 102.200 81.680 107.430 81.690 ;
        RECT 107.090 81.600 107.430 81.680 ;
        RECT 107.580 81.610 111.270 81.980 ;
        RECT 111.420 81.560 115.630 82.010 ;
        RECT 115.790 81.870 116.100 82.000 ;
        RECT 117.245 81.870 117.395 84.085 ;
        RECT 115.790 81.720 117.395 81.870 ;
        RECT 115.790 81.660 116.100 81.720 ;
        RECT 81.680 80.510 83.060 80.990 ;
        RECT 85.520 80.460 86.900 80.940 ;
        RECT 89.890 80.470 91.270 80.950 ;
        RECT 92.960 80.460 94.340 80.940 ;
        RECT 96.800 80.410 98.180 80.890 ;
        RECT 101.170 80.420 102.550 80.900 ;
        RECT 106.780 80.430 108.160 80.910 ;
        RECT 110.620 80.380 112.000 80.860 ;
        RECT 114.990 80.390 116.370 80.870 ;
        RECT 116.865 78.035 117.015 81.720 ;
        RECT 116.860 78.030 117.015 78.035 ;
        RECT 114.875 77.885 117.015 78.030 ;
        RECT 114.875 73.745 115.025 77.885 ;
        RECT 117.420 73.920 127.080 74.400 ;
        RECT 114.875 73.595 118.655 73.745 ;
        RECT 68.215 73.035 113.985 73.485 ;
        RECT 118.505 73.070 118.655 73.595 ;
        RECT 63.020 70.930 65.780 71.410 ;
        RECT 61.545 70.780 61.800 70.805 ;
        RECT 61.545 70.545 64.780 70.780 ;
        RECT 61.760 70.540 64.780 70.545 ;
        RECT 68.215 70.490 68.665 73.035 ;
        RECT 113.090 72.995 113.985 73.035 ;
        RECT 113.090 72.545 117.905 72.995 ;
        RECT 113.090 72.540 113.680 72.545 ;
        RECT 118.220 72.450 118.660 73.070 ;
        RECT 120.690 72.890 120.990 73.630 ;
        RECT 121.685 73.380 121.975 73.425 ;
        RECT 124.915 73.380 125.205 73.425 ;
        RECT 121.685 73.240 125.205 73.380 ;
        RECT 121.685 73.195 121.975 73.240 ;
        RECT 124.915 73.195 125.205 73.240 ;
        RECT 119.810 72.700 120.100 72.745 ;
        RECT 121.650 72.700 121.940 72.745 ;
        RECT 119.810 72.560 121.940 72.700 ;
        RECT 119.810 72.515 120.100 72.560 ;
        RECT 121.650 72.515 121.940 72.560 ;
        RECT 122.220 72.510 122.550 73.100 ;
        RECT 122.750 72.510 123.020 73.100 ;
        RECT 118.890 72.360 119.180 72.405 ;
        RECT 123.420 72.360 123.850 73.090 ;
        RECT 123.995 72.700 124.285 72.745 ;
        RECT 125.835 72.700 126.125 72.745 ;
        RECT 126.740 72.730 141.150 73.050 ;
        RECT 123.995 72.560 126.125 72.700 ;
        RECT 123.995 72.515 124.285 72.560 ;
        RECT 125.835 72.515 126.125 72.560 ;
        RECT 124.410 72.360 124.700 72.405 ;
        RECT 125.330 72.360 125.620 72.405 ;
        RECT 118.890 72.220 125.620 72.360 ;
        RECT 118.890 72.175 119.180 72.220 ;
        RECT 123.420 72.170 123.850 72.220 ;
        RECT 124.410 72.175 124.700 72.220 ;
        RECT 125.330 72.175 125.620 72.220 ;
        RECT 117.420 71.200 127.080 71.680 ;
        RECT 65.710 70.400 68.665 70.490 ;
        RECT 62.040 70.070 64.980 70.370 ;
        RECT 53.925 69.775 54.315 70.065 ;
        RECT 62.040 70.010 62.410 70.070 ;
        RECT 52.620 69.385 54.315 69.775 ;
        RECT 23.190 65.100 23.740 65.380 ;
        RECT 23.360 64.290 23.515 65.100 ;
        RECT 27.810 65.035 30.405 65.425 ;
        RECT 22.350 63.810 25.570 64.290 ;
        RECT 22.840 62.810 25.140 63.290 ;
        RECT 22.880 61.410 23.260 61.820 ;
        RECT 23.880 61.690 24.130 62.810 ;
        RECT 22.950 60.570 23.210 61.410 ;
        RECT 23.840 61.380 24.180 61.690 ;
        RECT 24.800 61.530 25.550 62.020 ;
        RECT 27.810 60.605 28.200 65.035 ;
        RECT 30.880 64.850 31.290 65.770 ;
        RECT 47.550 64.950 47.850 66.450 ;
        RECT 51.260 66.400 51.690 66.750 ;
        RECT 51.260 66.060 51.520 66.400 ;
        RECT 49.990 65.800 51.520 66.060 ;
        RECT 52.620 65.345 53.010 69.385 ;
        RECT 54.820 68.910 55.170 69.600 ;
        RECT 55.310 68.920 55.650 69.850 ;
        RECT 55.820 68.940 56.180 69.860 ;
        RECT 56.710 68.910 58.140 69.280 ;
        RECT 58.780 69.140 61.080 69.620 ;
        RECT 62.040 69.570 62.400 70.010 ;
        RECT 57.735 68.845 58.140 68.910 ;
        RECT 62.040 68.850 62.390 69.570 ;
        RECT 62.990 69.200 63.430 69.790 ;
        RECT 63.590 69.710 64.290 69.880 ;
        RECT 64.620 69.780 64.980 70.070 ;
        RECT 65.400 70.040 68.665 70.400 ;
        RECT 65.400 70.010 68.630 70.040 ;
        RECT 63.590 69.370 64.280 69.710 ;
        RECT 64.510 69.440 64.980 69.780 ;
        RECT 53.930 68.290 57.150 68.770 ;
        RECT 57.735 68.475 60.125 68.845 ;
        RECT 60.410 68.490 62.390 68.850 ;
        RECT 57.530 67.435 59.275 67.805 ;
        RECT 54.550 66.800 56.850 67.280 ;
        RECT 55.410 66.260 55.900 66.640 ;
        RECT 57.530 66.410 57.900 67.435 ;
        RECT 59.755 67.365 60.125 68.475 ;
        RECT 63.020 68.210 65.780 68.690 ;
        RECT 58.780 66.420 61.080 66.900 ;
        RECT 56.470 66.040 57.900 66.410 ;
        RECT 48.000 65.020 48.550 65.300 ;
        RECT 29.740 64.160 32.040 64.640 ;
        RECT 48.170 64.210 48.325 65.020 ;
        RECT 52.620 64.955 55.215 65.345 ;
        RECT 47.160 63.730 50.380 64.210 ;
        RECT 47.650 62.730 49.950 63.210 ;
        RECT 29.720 61.780 32.020 62.260 ;
        RECT 47.690 61.330 48.070 61.740 ;
        RECT 48.690 61.610 48.940 62.730 ;
        RECT 31.670 60.750 32.010 61.090 ;
        RECT 22.840 60.090 25.140 60.570 ;
        RECT 27.810 60.215 30.475 60.605 ;
        RECT 30.710 60.300 31.060 60.630 ;
        RECT 47.760 60.490 48.020 61.330 ;
        RECT 48.650 61.300 48.990 61.610 ;
        RECT 49.610 61.450 50.360 61.940 ;
        RECT 52.620 60.525 53.010 64.955 ;
        RECT 55.690 64.770 56.100 65.690 ;
        RECT 54.550 64.080 56.850 64.560 ;
        RECT 54.530 61.700 56.830 62.180 ;
        RECT 56.480 60.670 56.820 61.010 ;
        RECT 22.400 58.710 25.620 59.190 ;
        RECT 22.790 57.210 23.090 58.710 ;
        RECT 27.810 58.350 28.200 60.215 ;
        RECT 47.650 60.010 49.950 60.490 ;
        RECT 52.620 60.135 55.285 60.525 ;
        RECT 55.520 60.220 55.870 60.550 ;
        RECT 29.720 59.060 32.020 59.540 ;
        RECT 47.210 58.630 50.430 59.110 ;
        RECT 25.210 57.960 28.200 58.350 ;
        RECT 23.240 57.280 23.790 57.560 ;
        RECT 23.410 56.470 23.565 57.280 ;
        RECT 47.600 57.130 47.900 58.630 ;
        RECT 52.620 58.270 53.010 60.135 ;
        RECT 54.530 58.980 56.830 59.460 ;
        RECT 50.020 57.880 53.010 58.270 ;
        RECT 48.050 57.200 48.600 57.480 ;
        RECT 22.400 55.990 25.620 56.470 ;
        RECT 48.220 56.390 48.375 57.200 ;
        RECT 47.210 55.910 50.430 56.390 ;
        RECT 22.890 54.990 25.190 55.470 ;
        RECT 22.930 53.590 23.310 53.930 ;
        RECT 23.880 53.650 24.240 54.990 ;
        RECT 47.700 54.910 50.000 55.390 ;
        RECT 23.030 52.750 23.280 53.590 ;
        RECT 23.890 53.540 24.230 53.650 ;
        RECT 24.850 53.260 26.010 53.810 ;
        RECT 47.740 53.510 48.120 53.850 ;
        RECT 48.690 53.570 49.050 54.910 ;
        RECT 23.890 52.750 24.230 52.770 ;
        RECT 22.890 52.270 25.190 52.750 ;
        RECT 47.840 52.670 48.090 53.510 ;
        RECT 48.700 53.460 49.040 53.570 ;
        RECT 49.660 53.180 50.820 53.730 ;
        RECT 48.700 52.670 49.040 52.690 ;
        RECT 47.700 52.190 50.000 52.670 ;
        RECT 30.560 32.760 31.940 33.240 ;
        RECT 30.670 31.660 31.140 31.990 ;
        RECT 31.310 31.690 31.640 31.990 ;
        RECT 30.560 30.040 31.940 30.520 ;
        RECT 46.090 29.600 53.450 30.080 ;
        RECT 47.070 28.720 47.360 28.765 ;
        RECT 47.500 28.720 47.640 29.600 ;
        RECT 55.440 29.580 62.800 30.060 ;
        RECT 47.990 29.060 48.280 29.105 ;
        RECT 51.690 29.060 51.980 29.105 ;
        RECT 47.990 28.920 51.980 29.060 ;
        RECT 47.990 28.875 48.280 28.920 ;
        RECT 51.690 28.875 51.980 28.920 ;
        RECT 48.910 28.720 49.200 28.765 ;
        RECT 50.770 28.720 51.060 28.765 ;
        RECT 52.150 28.720 52.440 28.765 ;
        RECT 47.070 28.580 52.440 28.720 ;
        RECT 47.070 28.535 47.360 28.580 ;
        RECT 48.910 28.535 49.200 28.580 ;
        RECT 50.770 28.535 51.060 28.580 ;
        RECT 52.150 28.535 52.440 28.580 ;
        RECT 56.420 28.700 56.710 28.745 ;
        RECT 56.850 28.700 56.990 29.580 ;
        RECT 64.520 29.560 71.880 30.040 ;
        RECT 57.340 29.040 57.630 29.085 ;
        RECT 61.040 29.040 61.330 29.085 ;
        RECT 57.340 28.900 61.330 29.040 ;
        RECT 57.340 28.855 57.630 28.900 ;
        RECT 61.040 28.855 61.330 28.900 ;
        RECT 58.260 28.700 58.550 28.745 ;
        RECT 60.120 28.700 60.410 28.745 ;
        RECT 61.500 28.700 61.790 28.745 ;
        RECT 56.420 28.560 61.790 28.700 ;
        RECT 56.420 28.515 56.710 28.560 ;
        RECT 58.260 28.515 58.550 28.560 ;
        RECT 60.120 28.515 60.410 28.560 ;
        RECT 61.500 28.515 61.790 28.560 ;
        RECT 65.500 28.680 65.790 28.725 ;
        RECT 65.930 28.680 66.070 29.560 ;
        RECT 73.870 29.540 81.230 30.020 ;
        RECT 66.420 29.020 66.710 29.065 ;
        RECT 70.120 29.020 70.410 29.065 ;
        RECT 66.420 28.880 70.410 29.020 ;
        RECT 66.420 28.835 66.710 28.880 ;
        RECT 70.120 28.835 70.410 28.880 ;
        RECT 67.340 28.680 67.630 28.725 ;
        RECT 69.200 28.680 69.490 28.725 ;
        RECT 70.580 28.680 70.870 28.725 ;
        RECT 65.500 28.540 70.870 28.680 ;
        RECT 65.500 28.495 65.790 28.540 ;
        RECT 67.340 28.495 67.630 28.540 ;
        RECT 69.200 28.495 69.490 28.540 ;
        RECT 70.580 28.495 70.870 28.540 ;
        RECT 74.850 28.660 75.140 28.705 ;
        RECT 75.280 28.660 75.420 29.540 ;
        RECT 75.770 29.000 76.060 29.045 ;
        RECT 79.470 29.000 79.760 29.045 ;
        RECT 75.770 28.860 79.760 29.000 ;
        RECT 75.770 28.815 76.060 28.860 ;
        RECT 79.470 28.815 79.760 28.860 ;
        RECT 140.830 28.870 141.150 72.730 ;
        RECT 76.690 28.660 76.980 28.705 ;
        RECT 78.550 28.660 78.840 28.705 ;
        RECT 79.930 28.660 80.220 28.705 ;
        RECT 74.850 28.520 80.220 28.660 ;
        RECT 140.830 28.550 152.160 28.870 ;
        RECT 74.850 28.475 75.140 28.520 ;
        RECT 76.690 28.475 76.980 28.520 ;
        RECT 78.550 28.475 78.840 28.520 ;
        RECT 79.930 28.475 80.220 28.520 ;
        RECT 47.530 28.380 47.820 28.425 ;
        RECT 49.830 28.380 50.120 28.425 ;
        RECT 51.690 28.380 51.980 28.425 ;
        RECT 47.530 28.240 51.980 28.380 ;
        RECT 47.530 28.195 47.820 28.240 ;
        RECT 49.830 28.195 50.120 28.240 ;
        RECT 9.180 27.500 16.540 27.980 ;
        RECT 10.160 26.620 10.450 26.665 ;
        RECT 10.590 26.620 10.730 27.500 ;
        RECT 18.530 27.480 25.890 27.960 ;
        RECT 11.080 26.960 11.370 27.005 ;
        RECT 14.780 26.960 15.070 27.005 ;
        RECT 11.080 26.820 15.070 26.960 ;
        RECT 11.080 26.775 11.370 26.820 ;
        RECT 14.780 26.775 15.070 26.820 ;
        RECT 12.000 26.620 12.290 26.665 ;
        RECT 13.860 26.620 14.150 26.665 ;
        RECT 15.240 26.620 15.530 26.665 ;
        RECT 10.160 26.480 15.530 26.620 ;
        RECT 10.160 26.435 10.450 26.480 ;
        RECT 12.000 26.435 12.290 26.480 ;
        RECT 13.860 26.435 14.150 26.480 ;
        RECT 15.240 26.435 15.530 26.480 ;
        RECT 19.510 26.600 19.800 26.645 ;
        RECT 19.940 26.600 20.080 27.480 ;
        RECT 27.610 27.460 34.970 27.940 ;
        RECT 20.430 26.940 20.720 26.985 ;
        RECT 24.130 26.940 24.420 26.985 ;
        RECT 20.430 26.800 24.420 26.940 ;
        RECT 20.430 26.755 20.720 26.800 ;
        RECT 24.130 26.755 24.420 26.800 ;
        RECT 21.350 26.600 21.640 26.645 ;
        RECT 23.210 26.600 23.500 26.645 ;
        RECT 24.590 26.600 24.880 26.645 ;
        RECT 19.510 26.460 24.880 26.600 ;
        RECT 19.510 26.415 19.800 26.460 ;
        RECT 21.350 26.415 21.640 26.460 ;
        RECT 23.210 26.415 23.500 26.460 ;
        RECT 24.590 26.415 24.880 26.460 ;
        RECT 28.590 26.580 28.880 26.625 ;
        RECT 29.020 26.580 29.160 27.460 ;
        RECT 36.960 27.440 44.320 27.920 ;
        RECT 48.020 27.810 48.350 28.100 ;
        RECT 29.510 26.920 29.800 26.965 ;
        RECT 33.210 26.920 33.500 26.965 ;
        RECT 29.510 26.780 33.500 26.920 ;
        RECT 29.510 26.735 29.800 26.780 ;
        RECT 33.210 26.735 33.500 26.780 ;
        RECT 30.430 26.580 30.720 26.625 ;
        RECT 32.290 26.580 32.580 26.625 ;
        RECT 33.670 26.580 33.960 26.625 ;
        RECT 28.590 26.440 33.960 26.580 ;
        RECT 28.590 26.395 28.880 26.440 ;
        RECT 30.430 26.395 30.720 26.440 ;
        RECT 32.290 26.395 32.580 26.440 ;
        RECT 33.670 26.395 33.960 26.440 ;
        RECT 37.940 26.560 38.230 26.605 ;
        RECT 38.370 26.560 38.510 27.440 ;
        RECT 50.300 27.360 50.440 28.240 ;
        RECT 51.690 28.195 51.980 28.240 ;
        RECT 56.880 28.360 57.170 28.405 ;
        RECT 59.180 28.360 59.470 28.405 ;
        RECT 61.040 28.360 61.330 28.405 ;
        RECT 56.880 28.220 61.330 28.360 ;
        RECT 56.880 28.175 57.170 28.220 ;
        RECT 59.180 28.175 59.470 28.220 ;
        RECT 53.060 28.020 53.360 28.150 ;
        RECT 57.360 28.020 57.660 28.070 ;
        RECT 53.060 27.830 57.660 28.020 ;
        RECT 53.060 27.770 53.360 27.830 ;
        RECT 57.360 27.760 57.660 27.830 ;
        RECT 38.860 26.900 39.150 26.945 ;
        RECT 42.560 26.900 42.850 26.945 ;
        RECT 38.860 26.760 42.850 26.900 ;
        RECT 46.090 26.880 53.450 27.360 ;
        RECT 59.650 27.340 59.790 28.220 ;
        RECT 61.040 28.175 61.330 28.220 ;
        RECT 65.960 28.340 66.250 28.385 ;
        RECT 68.260 28.340 68.550 28.385 ;
        RECT 70.120 28.340 70.410 28.385 ;
        RECT 65.960 28.200 70.410 28.340 ;
        RECT 65.960 28.155 66.250 28.200 ;
        RECT 68.260 28.155 68.550 28.200 ;
        RECT 62.460 28.010 62.720 28.130 ;
        RECT 66.440 28.010 66.740 28.060 ;
        RECT 62.460 27.820 66.740 28.010 ;
        RECT 62.460 27.750 62.720 27.820 ;
        RECT 55.440 26.860 62.800 27.340 ;
        RECT 68.730 27.320 68.870 28.200 ;
        RECT 70.120 28.155 70.410 28.200 ;
        RECT 75.310 28.320 75.600 28.365 ;
        RECT 77.610 28.320 77.900 28.365 ;
        RECT 79.470 28.320 79.760 28.365 ;
        RECT 75.310 28.180 79.760 28.320 ;
        RECT 75.310 28.135 75.600 28.180 ;
        RECT 77.610 28.135 77.900 28.180 ;
        RECT 71.490 27.980 71.790 28.110 ;
        RECT 75.790 27.980 76.090 28.030 ;
        RECT 71.490 27.790 76.090 27.980 ;
        RECT 71.490 27.730 71.790 27.790 ;
        RECT 75.790 27.720 76.090 27.790 ;
        RECT 64.520 26.840 71.880 27.320 ;
        RECT 78.080 27.300 78.220 28.180 ;
        RECT 79.470 28.135 79.760 28.180 ;
        RECT 80.830 27.980 81.140 28.040 ;
        RECT 80.830 27.820 83.610 27.980 ;
        RECT 80.830 27.770 81.140 27.820 ;
        RECT 73.870 26.820 81.230 27.300 ;
        RECT 38.860 26.715 39.150 26.760 ;
        RECT 42.560 26.715 42.850 26.760 ;
        RECT 39.780 26.560 40.070 26.605 ;
        RECT 41.640 26.560 41.930 26.605 ;
        RECT 43.020 26.560 43.310 26.605 ;
        RECT 37.940 26.420 43.310 26.560 ;
        RECT 37.940 26.375 38.230 26.420 ;
        RECT 39.780 26.375 40.070 26.420 ;
        RECT 41.640 26.375 41.930 26.420 ;
        RECT 43.020 26.375 43.310 26.420 ;
        RECT 83.450 26.510 83.610 27.820 ;
        RECT 84.010 26.740 88.150 27.220 ;
        RECT 83.450 26.350 86.160 26.510 ;
        RECT 10.620 26.280 10.910 26.325 ;
        RECT 12.920 26.280 13.210 26.325 ;
        RECT 14.780 26.280 15.070 26.325 ;
        RECT 10.620 26.140 15.070 26.280 ;
        RECT 10.620 26.095 10.910 26.140 ;
        RECT 12.920 26.095 13.210 26.140 ;
        RECT 11.110 25.710 11.440 26.000 ;
        RECT 13.390 25.260 13.530 26.140 ;
        RECT 14.780 26.095 15.070 26.140 ;
        RECT 19.970 26.260 20.260 26.305 ;
        RECT 22.270 26.260 22.560 26.305 ;
        RECT 24.130 26.260 24.420 26.305 ;
        RECT 19.970 26.120 24.420 26.260 ;
        RECT 19.970 26.075 20.260 26.120 ;
        RECT 22.270 26.075 22.560 26.120 ;
        RECT 16.150 25.920 16.450 26.050 ;
        RECT 20.450 25.920 20.750 25.970 ;
        RECT 16.150 25.730 20.750 25.920 ;
        RECT 16.150 25.670 16.450 25.730 ;
        RECT 20.450 25.660 20.750 25.730 ;
        RECT 9.180 24.780 16.540 25.260 ;
        RECT 22.740 25.240 22.880 26.120 ;
        RECT 24.130 26.075 24.420 26.120 ;
        RECT 29.050 26.240 29.340 26.285 ;
        RECT 31.350 26.240 31.640 26.285 ;
        RECT 33.210 26.240 33.500 26.285 ;
        RECT 29.050 26.100 33.500 26.240 ;
        RECT 25.500 25.910 25.820 26.100 ;
        RECT 29.050 26.055 29.340 26.100 ;
        RECT 31.350 26.055 31.640 26.100 ;
        RECT 29.530 25.910 29.830 25.960 ;
        RECT 25.500 25.720 29.830 25.910 ;
        RECT 25.500 25.620 25.820 25.720 ;
        RECT 18.530 24.760 25.890 25.240 ;
        RECT 31.820 25.220 31.960 26.100 ;
        RECT 33.210 26.055 33.500 26.100 ;
        RECT 38.400 26.220 38.690 26.265 ;
        RECT 40.700 26.220 40.990 26.265 ;
        RECT 42.560 26.220 42.850 26.265 ;
        RECT 38.400 26.080 42.850 26.220 ;
        RECT 38.400 26.035 38.690 26.080 ;
        RECT 40.700 26.035 40.990 26.080 ;
        RECT 34.580 25.880 34.880 26.010 ;
        RECT 38.880 25.880 39.180 25.930 ;
        RECT 34.580 25.690 39.180 25.880 ;
        RECT 34.580 25.630 34.880 25.690 ;
        RECT 38.880 25.620 39.180 25.690 ;
        RECT 27.610 24.740 34.970 25.220 ;
        RECT 41.170 25.200 41.310 26.080 ;
        RECT 42.560 26.035 42.850 26.080 ;
        RECT 45.530 26.050 82.950 26.210 ;
        RECT 43.920 25.880 44.230 25.940 ;
        RECT 45.530 25.880 45.690 26.050 ;
        RECT 43.920 25.720 45.690 25.880 ;
        RECT 43.920 25.670 44.230 25.720 ;
        RECT 46.230 25.230 53.590 25.710 ;
        RECT 36.960 24.720 44.320 25.200 ;
        RECT 47.210 24.350 47.500 24.395 ;
        RECT 47.640 24.350 47.780 25.230 ;
        RECT 55.580 25.210 62.940 25.690 ;
        RECT 48.130 24.690 48.420 24.735 ;
        RECT 51.830 24.690 52.120 24.735 ;
        RECT 48.130 24.550 52.120 24.690 ;
        RECT 48.130 24.505 48.420 24.550 ;
        RECT 51.830 24.505 52.120 24.550 ;
        RECT 49.050 24.350 49.340 24.395 ;
        RECT 50.910 24.350 51.200 24.395 ;
        RECT 52.290 24.350 52.580 24.395 ;
        RECT 47.210 24.210 52.580 24.350 ;
        RECT 47.210 24.165 47.500 24.210 ;
        RECT 49.050 24.165 49.340 24.210 ;
        RECT 50.910 24.165 51.200 24.210 ;
        RECT 52.290 24.165 52.580 24.210 ;
        RECT 56.560 24.330 56.850 24.375 ;
        RECT 56.990 24.330 57.130 25.210 ;
        RECT 64.660 25.190 72.020 25.670 ;
        RECT 57.480 24.670 57.770 24.715 ;
        RECT 61.180 24.670 61.470 24.715 ;
        RECT 57.480 24.530 61.470 24.670 ;
        RECT 57.480 24.485 57.770 24.530 ;
        RECT 61.180 24.485 61.470 24.530 ;
        RECT 58.400 24.330 58.690 24.375 ;
        RECT 60.260 24.330 60.550 24.375 ;
        RECT 61.640 24.330 61.930 24.375 ;
        RECT 56.560 24.190 61.930 24.330 ;
        RECT 56.560 24.145 56.850 24.190 ;
        RECT 58.400 24.145 58.690 24.190 ;
        RECT 60.260 24.145 60.550 24.190 ;
        RECT 61.640 24.145 61.930 24.190 ;
        RECT 65.640 24.310 65.930 24.355 ;
        RECT 66.070 24.310 66.210 25.190 ;
        RECT 74.010 25.170 81.370 25.650 ;
        RECT 82.605 25.540 82.950 26.050 ;
        RECT 85.490 25.670 85.740 26.210 ;
        RECT 84.630 25.540 84.900 25.600 ;
        RECT 82.605 25.350 85.360 25.540 ;
        RECT 84.630 25.270 84.900 25.350 ;
        RECT 66.560 24.650 66.850 24.695 ;
        RECT 70.260 24.650 70.550 24.695 ;
        RECT 66.560 24.510 70.550 24.650 ;
        RECT 66.560 24.465 66.850 24.510 ;
        RECT 70.260 24.465 70.550 24.510 ;
        RECT 67.480 24.310 67.770 24.355 ;
        RECT 69.340 24.310 69.630 24.355 ;
        RECT 70.720 24.310 71.010 24.355 ;
        RECT 65.640 24.170 71.010 24.310 ;
        RECT 65.640 24.125 65.930 24.170 ;
        RECT 67.480 24.125 67.770 24.170 ;
        RECT 69.340 24.125 69.630 24.170 ;
        RECT 70.720 24.125 71.010 24.170 ;
        RECT 74.990 24.290 75.280 24.335 ;
        RECT 75.420 24.290 75.560 25.170 ;
        RECT 85.540 25.120 85.700 25.670 ;
        RECT 85.890 25.570 86.160 26.350 ;
        RECT 85.890 25.550 86.080 25.570 ;
        RECT 82.790 24.960 85.700 25.120 ;
        RECT 75.910 24.630 76.200 24.675 ;
        RECT 79.610 24.630 79.900 24.675 ;
        RECT 75.910 24.490 79.900 24.630 ;
        RECT 75.910 24.445 76.200 24.490 ;
        RECT 79.610 24.445 79.900 24.490 ;
        RECT 76.830 24.290 77.120 24.335 ;
        RECT 78.690 24.290 78.980 24.335 ;
        RECT 80.070 24.290 80.360 24.335 ;
        RECT 74.990 24.150 80.360 24.290 ;
        RECT 74.990 24.105 75.280 24.150 ;
        RECT 76.830 24.105 77.120 24.150 ;
        RECT 78.690 24.105 78.980 24.150 ;
        RECT 80.070 24.105 80.360 24.150 ;
        RECT 47.670 24.010 47.960 24.055 ;
        RECT 49.970 24.010 50.260 24.055 ;
        RECT 51.830 24.010 52.120 24.055 ;
        RECT 47.670 23.870 52.120 24.010 ;
        RECT 47.670 23.825 47.960 23.870 ;
        RECT 49.970 23.825 50.260 23.870 ;
        RECT 48.160 23.440 48.490 23.730 ;
        RECT 50.440 22.990 50.580 23.870 ;
        RECT 51.830 23.825 52.120 23.870 ;
        RECT 57.020 23.990 57.310 24.035 ;
        RECT 59.320 23.990 59.610 24.035 ;
        RECT 61.180 23.990 61.470 24.035 ;
        RECT 57.020 23.850 61.470 23.990 ;
        RECT 57.020 23.805 57.310 23.850 ;
        RECT 59.320 23.805 59.610 23.850 ;
        RECT 53.200 23.650 53.500 23.780 ;
        RECT 57.500 23.650 57.800 23.700 ;
        RECT 53.200 23.460 57.800 23.650 ;
        RECT 53.200 23.400 53.500 23.460 ;
        RECT 57.500 23.390 57.800 23.460 ;
        RECT 46.230 22.510 53.590 22.990 ;
        RECT 59.790 22.970 59.930 23.850 ;
        RECT 61.180 23.805 61.470 23.850 ;
        RECT 66.100 23.970 66.390 24.015 ;
        RECT 68.400 23.970 68.690 24.015 ;
        RECT 70.260 23.970 70.550 24.015 ;
        RECT 66.100 23.830 70.550 23.970 ;
        RECT 66.100 23.785 66.390 23.830 ;
        RECT 68.400 23.785 68.690 23.830 ;
        RECT 62.590 23.640 62.860 23.710 ;
        RECT 66.580 23.640 66.880 23.690 ;
        RECT 62.590 23.450 66.880 23.640 ;
        RECT 62.590 23.350 62.860 23.450 ;
        RECT 55.580 22.490 62.940 22.970 ;
        RECT 68.870 22.950 69.010 23.830 ;
        RECT 70.260 23.785 70.550 23.830 ;
        RECT 75.450 23.950 75.740 23.995 ;
        RECT 77.750 23.950 78.040 23.995 ;
        RECT 79.610 23.950 79.900 23.995 ;
        RECT 75.450 23.810 79.900 23.950 ;
        RECT 75.450 23.765 75.740 23.810 ;
        RECT 77.750 23.765 78.040 23.810 ;
        RECT 71.630 23.610 71.930 23.740 ;
        RECT 75.930 23.610 76.230 23.660 ;
        RECT 71.630 23.420 76.230 23.610 ;
        RECT 71.630 23.360 71.930 23.420 ;
        RECT 75.930 23.350 76.230 23.420 ;
        RECT 64.660 22.470 72.020 22.950 ;
        RECT 78.220 22.930 78.360 23.810 ;
        RECT 79.610 23.765 79.900 23.810 ;
        RECT 80.970 23.610 81.280 23.670 ;
        RECT 82.790 23.610 82.950 24.960 ;
        RECT 87.730 24.720 88.060 25.490 ;
        RECT 84.010 24.020 88.150 24.500 ;
        RECT 80.970 23.450 82.950 23.610 ;
        RECT 80.970 23.400 81.280 23.450 ;
        RECT 74.010 22.450 81.370 22.930 ;
        RECT 30.410 16.460 31.790 16.940 ;
        RECT 30.520 15.360 30.990 15.690 ;
        RECT 31.160 15.390 31.490 15.690 ;
        RECT 30.410 13.740 31.790 14.220 ;
        RECT 9.030 11.200 16.390 11.680 ;
        RECT 10.010 10.320 10.300 10.365 ;
        RECT 10.440 10.320 10.580 11.200 ;
        RECT 18.380 11.180 25.740 11.660 ;
        RECT 10.930 10.660 11.220 10.705 ;
        RECT 14.630 10.660 14.920 10.705 ;
        RECT 10.930 10.520 14.920 10.660 ;
        RECT 10.930 10.475 11.220 10.520 ;
        RECT 14.630 10.475 14.920 10.520 ;
        RECT 11.850 10.320 12.140 10.365 ;
        RECT 13.710 10.320 14.000 10.365 ;
        RECT 15.090 10.320 15.380 10.365 ;
        RECT 10.010 10.180 15.380 10.320 ;
        RECT 10.010 10.135 10.300 10.180 ;
        RECT 11.850 10.135 12.140 10.180 ;
        RECT 13.710 10.135 14.000 10.180 ;
        RECT 15.090 10.135 15.380 10.180 ;
        RECT 19.360 10.300 19.650 10.345 ;
        RECT 19.790 10.300 19.930 11.180 ;
        RECT 27.460 11.160 34.820 11.640 ;
        RECT 20.280 10.640 20.570 10.685 ;
        RECT 23.980 10.640 24.270 10.685 ;
        RECT 20.280 10.500 24.270 10.640 ;
        RECT 20.280 10.455 20.570 10.500 ;
        RECT 23.980 10.455 24.270 10.500 ;
        RECT 21.200 10.300 21.490 10.345 ;
        RECT 23.060 10.300 23.350 10.345 ;
        RECT 24.440 10.300 24.730 10.345 ;
        RECT 19.360 10.160 24.730 10.300 ;
        RECT 19.360 10.115 19.650 10.160 ;
        RECT 21.200 10.115 21.490 10.160 ;
        RECT 23.060 10.115 23.350 10.160 ;
        RECT 24.440 10.115 24.730 10.160 ;
        RECT 28.440 10.280 28.730 10.325 ;
        RECT 28.870 10.280 29.010 11.160 ;
        RECT 36.810 11.140 44.170 11.620 ;
        RECT 29.360 10.620 29.650 10.665 ;
        RECT 33.060 10.620 33.350 10.665 ;
        RECT 29.360 10.480 33.350 10.620 ;
        RECT 29.360 10.435 29.650 10.480 ;
        RECT 33.060 10.435 33.350 10.480 ;
        RECT 30.280 10.280 30.570 10.325 ;
        RECT 32.140 10.280 32.430 10.325 ;
        RECT 33.520 10.280 33.810 10.325 ;
        RECT 28.440 10.140 33.810 10.280 ;
        RECT 28.440 10.095 28.730 10.140 ;
        RECT 30.280 10.095 30.570 10.140 ;
        RECT 32.140 10.095 32.430 10.140 ;
        RECT 33.520 10.095 33.810 10.140 ;
        RECT 37.790 10.260 38.080 10.305 ;
        RECT 38.220 10.260 38.360 11.140 ;
        RECT 45.880 11.130 53.240 11.610 ;
        RECT 38.710 10.600 39.000 10.645 ;
        RECT 42.410 10.600 42.700 10.645 ;
        RECT 38.710 10.460 42.700 10.600 ;
        RECT 38.710 10.415 39.000 10.460 ;
        RECT 42.410 10.415 42.700 10.460 ;
        RECT 39.630 10.260 39.920 10.305 ;
        RECT 41.490 10.260 41.780 10.305 ;
        RECT 42.870 10.260 43.160 10.305 ;
        RECT 37.790 10.120 43.160 10.260 ;
        RECT 37.790 10.075 38.080 10.120 ;
        RECT 39.630 10.075 39.920 10.120 ;
        RECT 41.490 10.075 41.780 10.120 ;
        RECT 42.870 10.075 43.160 10.120 ;
        RECT 46.860 10.250 47.150 10.295 ;
        RECT 47.290 10.250 47.430 11.130 ;
        RECT 55.230 11.110 62.590 11.590 ;
        RECT 47.780 10.590 48.070 10.635 ;
        RECT 51.480 10.590 51.770 10.635 ;
        RECT 47.780 10.450 51.770 10.590 ;
        RECT 47.780 10.405 48.070 10.450 ;
        RECT 51.480 10.405 51.770 10.450 ;
        RECT 48.700 10.250 48.990 10.295 ;
        RECT 50.560 10.250 50.850 10.295 ;
        RECT 51.940 10.250 52.230 10.295 ;
        RECT 46.860 10.110 52.230 10.250 ;
        RECT 46.860 10.065 47.150 10.110 ;
        RECT 48.700 10.065 48.990 10.110 ;
        RECT 50.560 10.065 50.850 10.110 ;
        RECT 51.940 10.065 52.230 10.110 ;
        RECT 56.210 10.230 56.500 10.275 ;
        RECT 56.640 10.230 56.780 11.110 ;
        RECT 64.310 11.090 71.670 11.570 ;
        RECT 57.130 10.570 57.420 10.615 ;
        RECT 60.830 10.570 61.120 10.615 ;
        RECT 57.130 10.430 61.120 10.570 ;
        RECT 57.130 10.385 57.420 10.430 ;
        RECT 60.830 10.385 61.120 10.430 ;
        RECT 58.050 10.230 58.340 10.275 ;
        RECT 59.910 10.230 60.200 10.275 ;
        RECT 61.290 10.230 61.580 10.275 ;
        RECT 56.210 10.090 61.580 10.230 ;
        RECT 56.210 10.045 56.500 10.090 ;
        RECT 58.050 10.045 58.340 10.090 ;
        RECT 59.910 10.045 60.200 10.090 ;
        RECT 61.290 10.045 61.580 10.090 ;
        RECT 65.290 10.210 65.580 10.255 ;
        RECT 65.720 10.210 65.860 11.090 ;
        RECT 73.660 11.070 81.020 11.550 ;
        RECT 66.210 10.550 66.500 10.595 ;
        RECT 69.910 10.550 70.200 10.595 ;
        RECT 66.210 10.410 70.200 10.550 ;
        RECT 66.210 10.365 66.500 10.410 ;
        RECT 69.910 10.365 70.200 10.410 ;
        RECT 67.130 10.210 67.420 10.255 ;
        RECT 68.990 10.210 69.280 10.255 ;
        RECT 70.370 10.210 70.660 10.255 ;
        RECT 65.290 10.070 70.660 10.210 ;
        RECT 65.290 10.025 65.580 10.070 ;
        RECT 67.130 10.025 67.420 10.070 ;
        RECT 68.990 10.025 69.280 10.070 ;
        RECT 70.370 10.025 70.660 10.070 ;
        RECT 74.640 10.190 74.930 10.235 ;
        RECT 75.070 10.190 75.210 11.070 ;
        RECT 75.560 10.530 75.850 10.575 ;
        RECT 79.260 10.530 79.550 10.575 ;
        RECT 75.560 10.390 79.550 10.530 ;
        RECT 75.560 10.345 75.850 10.390 ;
        RECT 79.260 10.345 79.550 10.390 ;
        RECT 76.480 10.190 76.770 10.235 ;
        RECT 78.340 10.190 78.630 10.235 ;
        RECT 79.720 10.190 80.010 10.235 ;
        RECT 74.640 10.050 80.010 10.190 ;
        RECT 10.470 9.980 10.760 10.025 ;
        RECT 12.770 9.980 13.060 10.025 ;
        RECT 14.630 9.980 14.920 10.025 ;
        RECT 74.640 10.005 74.930 10.050 ;
        RECT 76.480 10.005 76.770 10.050 ;
        RECT 78.340 10.005 78.630 10.050 ;
        RECT 79.720 10.005 80.010 10.050 ;
        RECT 10.470 9.840 14.920 9.980 ;
        RECT 10.470 9.795 10.760 9.840 ;
        RECT 12.770 9.795 13.060 9.840 ;
        RECT 10.960 9.410 11.290 9.700 ;
        RECT 13.240 8.960 13.380 9.840 ;
        RECT 14.630 9.795 14.920 9.840 ;
        RECT 19.820 9.960 20.110 10.005 ;
        RECT 22.120 9.960 22.410 10.005 ;
        RECT 23.980 9.960 24.270 10.005 ;
        RECT 19.820 9.820 24.270 9.960 ;
        RECT 19.820 9.775 20.110 9.820 ;
        RECT 22.120 9.775 22.410 9.820 ;
        RECT 16.000 9.620 16.300 9.750 ;
        RECT 20.300 9.620 20.600 9.670 ;
        RECT 16.000 9.430 20.600 9.620 ;
        RECT 16.000 9.370 16.300 9.430 ;
        RECT 20.300 9.360 20.600 9.430 ;
        RECT 9.030 8.480 16.390 8.960 ;
        RECT 22.590 8.940 22.730 9.820 ;
        RECT 23.980 9.775 24.270 9.820 ;
        RECT 28.900 9.940 29.190 9.985 ;
        RECT 31.200 9.940 31.490 9.985 ;
        RECT 33.060 9.940 33.350 9.985 ;
        RECT 28.900 9.800 33.350 9.940 ;
        RECT 28.900 9.755 29.190 9.800 ;
        RECT 31.200 9.755 31.490 9.800 ;
        RECT 25.390 9.610 25.650 9.700 ;
        RECT 29.380 9.610 29.680 9.660 ;
        RECT 25.390 9.420 29.680 9.610 ;
        RECT 25.390 9.370 25.650 9.420 ;
        RECT 18.380 8.460 25.740 8.940 ;
        RECT 31.670 8.920 31.810 9.800 ;
        RECT 33.060 9.755 33.350 9.800 ;
        RECT 38.250 9.920 38.540 9.965 ;
        RECT 40.550 9.920 40.840 9.965 ;
        RECT 42.410 9.920 42.700 9.965 ;
        RECT 38.250 9.780 42.700 9.920 ;
        RECT 38.250 9.735 38.540 9.780 ;
        RECT 40.550 9.735 40.840 9.780 ;
        RECT 34.430 9.580 34.730 9.710 ;
        RECT 38.730 9.580 39.030 9.630 ;
        RECT 34.430 9.390 39.030 9.580 ;
        RECT 34.430 9.330 34.730 9.390 ;
        RECT 38.730 9.320 39.030 9.390 ;
        RECT 27.460 8.440 34.820 8.920 ;
        RECT 41.020 8.900 41.160 9.780 ;
        RECT 42.410 9.735 42.700 9.780 ;
        RECT 47.320 9.910 47.610 9.955 ;
        RECT 49.620 9.910 49.910 9.955 ;
        RECT 51.480 9.910 51.770 9.955 ;
        RECT 47.320 9.770 51.770 9.910 ;
        RECT 47.320 9.725 47.610 9.770 ;
        RECT 49.620 9.725 49.910 9.770 ;
        RECT 43.770 9.580 44.080 9.640 ;
        RECT 47.810 9.580 48.140 9.630 ;
        RECT 43.770 9.420 48.140 9.580 ;
        RECT 43.770 9.370 44.080 9.420 ;
        RECT 47.810 9.380 48.140 9.420 ;
        RECT 36.810 8.420 44.170 8.900 ;
        RECT 50.090 8.890 50.230 9.770 ;
        RECT 51.480 9.725 51.770 9.770 ;
        RECT 56.670 9.890 56.960 9.935 ;
        RECT 58.970 9.890 59.260 9.935 ;
        RECT 60.830 9.890 61.120 9.935 ;
        RECT 56.670 9.750 61.120 9.890 ;
        RECT 56.670 9.705 56.960 9.750 ;
        RECT 58.970 9.705 59.260 9.750 ;
        RECT 52.850 9.550 53.150 9.680 ;
        RECT 57.150 9.550 57.450 9.600 ;
        RECT 52.850 9.360 57.450 9.550 ;
        RECT 52.850 9.300 53.150 9.360 ;
        RECT 57.150 9.290 57.450 9.360 ;
        RECT 45.880 8.410 53.240 8.890 ;
        RECT 59.440 8.870 59.580 9.750 ;
        RECT 60.830 9.705 61.120 9.750 ;
        RECT 65.750 9.870 66.040 9.915 ;
        RECT 68.050 9.870 68.340 9.915 ;
        RECT 69.910 9.870 70.200 9.915 ;
        RECT 65.750 9.730 70.200 9.870 ;
        RECT 65.750 9.685 66.040 9.730 ;
        RECT 68.050 9.685 68.340 9.730 ;
        RECT 62.220 9.540 62.500 9.650 ;
        RECT 66.230 9.540 66.530 9.590 ;
        RECT 62.220 9.350 66.530 9.540 ;
        RECT 62.220 9.320 62.500 9.350 ;
        RECT 55.230 8.390 62.590 8.870 ;
        RECT 68.520 8.850 68.660 9.730 ;
        RECT 69.910 9.685 70.200 9.730 ;
        RECT 75.100 9.850 75.390 9.895 ;
        RECT 77.400 9.850 77.690 9.895 ;
        RECT 79.260 9.850 79.550 9.895 ;
        RECT 75.100 9.710 79.550 9.850 ;
        RECT 75.100 9.665 75.390 9.710 ;
        RECT 77.400 9.665 77.690 9.710 ;
        RECT 71.280 9.510 71.580 9.640 ;
        RECT 75.580 9.510 75.880 9.560 ;
        RECT 71.280 9.320 75.880 9.510 ;
        RECT 71.280 9.260 71.580 9.320 ;
        RECT 75.580 9.250 75.880 9.320 ;
        RECT 64.310 8.370 71.670 8.850 ;
        RECT 77.870 8.830 78.010 9.710 ;
        RECT 79.260 9.665 79.550 9.710 ;
        RECT 80.680 9.340 82.050 9.650 ;
        RECT 73.660 8.350 81.020 8.830 ;
        RECT 151.840 4.310 152.160 28.550 ;
        RECT 151.150 3.190 152.710 4.310 ;
      LAYER met2 ;
        RECT 47.150 88.730 48.530 89.220 ;
        RECT 32.315 87.935 32.725 87.940 ;
        RECT 32.315 87.930 33.795 87.935 ;
        RECT 32.315 87.525 33.800 87.930 ;
        RECT 22.360 82.680 23.660 83.180 ;
        RECT 29.730 81.560 30.740 82.190 ;
        RECT 24.430 79.970 25.530 80.450 ;
        RECT 22.810 78.960 24.690 79.400 ;
        RECT 24.790 77.360 25.330 77.550 ;
        RECT 24.790 77.180 27.290 77.360 ;
        RECT 24.180 76.270 25.140 76.750 ;
        RECT 22.380 74.890 23.750 75.350 ;
        RECT 24.730 72.170 25.590 72.620 ;
        RECT 22.880 71.160 24.350 71.600 ;
        RECT 27.110 70.490 27.290 77.180 ;
        RECT 28.740 73.200 29.540 73.680 ;
        RECT 30.050 72.550 30.390 81.560 ;
        RECT 32.315 77.120 32.725 87.525 ;
        RECT 33.020 87.490 33.800 87.525 ;
        RECT 47.160 86.010 48.530 86.510 ;
        RECT 57.005 85.270 57.415 85.275 ;
        RECT 57.000 85.165 57.530 85.270 ;
        RECT 57.000 83.810 57.535 85.165 ;
        RECT 47.170 82.600 48.470 83.100 ;
        RECT 54.540 81.480 55.550 82.110 ;
        RECT 49.240 79.890 50.340 80.370 ;
        RECT 33.040 78.420 34.470 78.900 ;
        RECT 47.620 78.880 49.500 79.320 ;
        RECT 49.600 77.280 50.140 77.470 ;
        RECT 32.315 76.710 33.410 77.120 ;
        RECT 49.600 77.100 52.100 77.280 ;
        RECT 30.540 75.920 31.270 76.400 ;
        RECT 48.990 76.190 49.950 76.670 ;
        RECT 35.230 75.700 36.260 76.190 ;
        RECT 47.190 74.810 48.560 75.270 ;
        RECT 30.050 72.210 30.840 72.550 ;
        RECT 27.110 70.310 30.160 70.490 ;
        RECT 29.980 69.680 30.160 70.310 ;
        RECT 24.840 69.400 25.690 69.560 ;
        RECT 29.980 69.400 30.360 69.680 ;
        RECT 24.840 69.160 28.570 69.400 ;
        RECT 29.970 69.160 30.360 69.400 ;
        RECT 24.840 69.090 25.690 69.160 ;
        RECT 24.100 68.420 25.200 68.900 ;
        RECT 28.320 67.960 28.560 69.160 ;
        RECT 30.010 68.970 30.360 69.160 ;
        RECT 30.500 68.960 30.840 72.210 ;
        RECT 38.175 72.435 42.655 72.905 ;
        RECT 31.610 71.090 32.350 71.580 ;
        RECT 31.005 69.005 31.375 69.925 ;
        RECT 33.970 69.210 34.730 69.690 ;
        RECT 38.175 69.285 38.645 72.435 ;
        RECT 39.200 71.020 40.360 71.480 ;
        RECT 38.790 69.450 39.480 69.960 ;
        RECT 29.120 68.360 29.870 68.850 ;
        RECT 31.005 68.635 31.715 69.005 ;
        RECT 28.320 67.720 30.870 67.960 ;
        RECT 22.340 66.550 23.690 66.980 ;
        RECT 29.750 66.890 30.420 67.350 ;
        RECT 30.630 66.860 30.870 67.720 ;
        RECT 26.800 66.830 28.830 66.840 ;
        RECT 26.450 66.480 28.830 66.830 ;
        RECT 28.470 65.850 28.830 66.480 ;
        RECT 30.600 66.340 31.090 66.860 ;
        RECT 31.345 65.860 31.715 68.635 ;
        RECT 38.210 68.290 38.720 68.770 ;
        RECT 35.480 66.500 36.240 66.980 ;
        RECT 30.700 65.850 31.715 65.860 ;
        RECT 28.470 65.490 31.715 65.850 ;
        RECT 30.930 64.720 31.290 65.490 ;
        RECT 24.610 63.830 25.560 64.270 ;
        RECT 29.740 64.170 30.500 64.640 ;
        RECT 22.870 62.800 23.900 63.270 ;
        RECT 24.800 61.690 25.550 62.020 ;
        RECT 31.150 61.780 32.010 62.260 ;
        RECT 24.800 61.530 30.950 61.690 ;
        RECT 30.790 60.630 30.950 61.530 ;
        RECT 38.890 61.090 39.230 69.450 ;
        RECT 31.670 60.750 39.230 61.090 ;
        RECT 24.290 60.110 25.120 60.580 ;
        RECT 30.710 60.300 31.060 60.630 ;
        RECT 22.550 58.730 23.450 59.170 ;
        RECT 29.720 59.060 30.500 59.540 ;
        RECT 24.690 56.020 25.590 56.460 ;
        RECT 22.900 54.980 23.880 55.460 ;
        RECT 42.185 53.810 42.655 72.435 ;
        RECT 49.540 72.090 50.400 72.540 ;
        RECT 47.690 71.080 49.160 71.520 ;
        RECT 51.920 70.410 52.100 77.100 ;
        RECT 53.550 73.120 54.350 73.600 ;
        RECT 54.860 72.470 55.200 81.480 ;
        RECT 57.125 77.040 57.535 83.810 ;
        RECT 81.730 83.230 82.790 83.690 ;
        RECT 85.580 83.200 86.640 83.660 ;
        RECT 90.040 83.200 91.100 83.660 ;
        RECT 93.010 83.180 94.070 83.640 ;
        RECT 96.860 83.150 97.920 83.610 ;
        RECT 101.320 83.150 102.380 83.610 ;
        RECT 106.830 83.150 107.890 83.610 ;
        RECT 110.680 83.120 111.740 83.580 ;
        RECT 115.140 83.120 116.200 83.580 ;
        RECT 81.680 80.510 82.740 80.970 ;
        RECT 85.630 80.470 86.690 80.930 ;
        RECT 89.980 80.470 91.040 80.930 ;
        RECT 92.960 80.460 94.020 80.920 ;
        RECT 96.910 80.420 97.970 80.880 ;
        RECT 101.260 80.420 102.320 80.880 ;
        RECT 106.780 80.430 107.840 80.890 ;
        RECT 110.730 80.390 111.790 80.850 ;
        RECT 115.080 80.390 116.140 80.850 ;
        RECT 57.850 78.340 59.280 78.820 ;
        RECT 57.125 76.630 58.220 77.040 ;
        RECT 55.350 75.840 56.080 76.320 ;
        RECT 60.040 75.620 61.070 76.110 ;
        RECT 129.880 74.760 136.950 75.100 ;
        RECT 121.560 73.940 122.710 74.400 ;
        RECT 129.880 73.630 130.220 74.760 ;
        RECT 134.740 73.630 135.860 73.970 ;
        RECT 120.690 73.290 130.220 73.630 ;
        RECT 132.040 73.290 135.880 73.630 ;
        RECT 65.710 72.825 67.170 72.905 ;
        RECT 54.860 72.130 55.650 72.470 ;
        RECT 51.920 70.230 54.970 70.410 ;
        RECT 54.790 69.600 54.970 70.230 ;
        RECT 49.650 69.320 50.500 69.480 ;
        RECT 54.790 69.320 55.170 69.600 ;
        RECT 49.650 69.080 53.380 69.320 ;
        RECT 54.780 69.080 55.170 69.320 ;
        RECT 49.650 69.010 50.500 69.080 ;
        RECT 48.910 68.340 50.010 68.820 ;
        RECT 53.130 67.880 53.370 69.080 ;
        RECT 54.820 68.890 55.170 69.080 ;
        RECT 55.310 68.880 55.650 72.130 ;
        RECT 62.985 72.355 67.465 72.825 ;
        RECT 120.690 72.440 120.990 73.290 ;
        RECT 56.420 71.010 57.160 71.500 ;
        RECT 55.815 68.925 56.185 69.845 ;
        RECT 58.780 69.130 59.540 69.610 ;
        RECT 62.985 69.205 63.455 72.355 ;
        RECT 64.010 70.940 65.170 71.400 ;
        RECT 63.600 69.370 64.290 69.880 ;
        RECT 53.930 68.280 54.680 68.770 ;
        RECT 55.815 68.555 56.525 68.925 ;
        RECT 53.130 67.640 55.680 67.880 ;
        RECT 47.150 66.470 48.500 66.900 ;
        RECT 54.560 66.810 55.230 67.270 ;
        RECT 55.440 66.780 55.680 67.640 ;
        RECT 51.610 66.750 53.640 66.760 ;
        RECT 51.260 66.400 53.640 66.750 ;
        RECT 53.280 65.770 53.640 66.400 ;
        RECT 55.410 66.260 55.900 66.780 ;
        RECT 56.155 65.780 56.525 68.555 ;
        RECT 63.020 68.210 63.530 68.690 ;
        RECT 60.290 66.420 61.050 66.900 ;
        RECT 55.510 65.770 56.525 65.780 ;
        RECT 53.280 65.410 56.525 65.770 ;
        RECT 55.740 64.640 56.100 65.410 ;
        RECT 49.420 63.750 50.370 64.190 ;
        RECT 54.550 64.090 55.310 64.560 ;
        RECT 47.680 62.720 48.710 63.190 ;
        RECT 49.610 61.610 50.360 61.940 ;
        RECT 55.960 61.700 56.820 62.180 ;
        RECT 49.610 61.450 55.760 61.610 ;
        RECT 55.600 60.550 55.760 61.450 ;
        RECT 63.700 61.010 64.040 69.370 ;
        RECT 56.480 60.670 64.040 61.010 ;
        RECT 49.100 60.030 49.930 60.500 ;
        RECT 55.520 60.220 55.870 60.550 ;
        RECT 47.360 58.650 48.260 59.090 ;
        RECT 54.530 58.980 55.310 59.460 ;
        RECT 49.500 55.940 50.400 56.380 ;
        RECT 47.710 54.900 48.690 55.380 ;
        RECT 66.705 53.810 67.465 72.355 ;
        RECT 119.250 71.200 121.060 71.670 ;
        RECT 122.240 70.560 122.520 73.100 ;
        RECT 122.240 70.280 122.510 70.560 ;
        RECT 24.850 53.340 42.655 53.810 ;
        RECT 65.710 53.730 67.465 53.810 ;
        RECT 24.850 53.260 26.010 53.340 ;
        RECT 49.660 53.260 67.465 53.730 ;
        RECT 116.290 70.000 122.510 70.280 ;
        RECT 49.660 53.180 50.820 53.260 ;
        RECT 24.280 52.290 25.180 52.730 ;
        RECT 49.090 52.210 49.990 52.650 ;
        RECT 30.560 32.790 31.940 33.240 ;
        RECT 27.925 31.990 28.255 32.020 ;
        RECT 11.110 31.660 31.140 31.990 ;
        RECT 31.310 31.970 65.780 31.990 ;
        RECT 116.290 31.970 116.570 70.000 ;
        RECT 122.730 66.450 123.030 73.110 ;
        RECT 123.420 72.570 123.880 73.120 ;
        RECT 132.040 72.570 132.380 73.290 ;
        RECT 134.740 73.020 135.860 73.290 ;
        RECT 123.420 72.180 132.380 72.570 ;
        RECT 136.610 72.570 136.950 74.760 ;
        RECT 136.610 72.550 138.020 72.570 ;
        RECT 136.610 72.180 138.650 72.550 ;
        RECT 132.040 72.160 132.380 72.180 ;
        RECT 137.560 71.680 138.650 72.180 ;
        RECT 31.310 31.690 116.570 31.970 ;
        RECT 121.260 66.150 123.040 66.450 ;
        RECT 11.110 25.710 11.450 31.660 ;
        RECT 30.550 30.090 31.370 30.520 ;
        RECT 12.550 27.510 13.450 27.980 ;
        RECT 21.890 27.490 22.790 27.960 ;
        RECT 30.510 27.470 31.410 27.940 ;
        RECT 40.050 27.450 40.950 27.920 ;
        RECT 48.020 27.810 48.360 30.090 ;
        RECT 49.540 29.610 50.440 30.080 ;
        RECT 59.000 29.550 59.910 30.030 ;
        RECT 67.850 29.570 68.760 30.050 ;
        RECT 77.320 29.560 78.220 30.020 ;
        RECT 51.710 26.890 52.620 27.370 ;
        RECT 56.560 26.860 57.470 27.340 ;
        RECT 70.080 26.830 70.990 27.310 ;
        RECT 74.680 26.810 75.590 27.290 ;
        RECT 85.790 26.740 86.690 27.220 ;
        RECT 88.465 25.875 88.740 31.690 ;
        RECT 12.600 24.780 13.500 25.250 ;
        RECT 46.640 25.230 47.540 25.710 ;
        RECT 21.890 24.760 22.790 25.230 ;
        RECT 30.460 24.750 31.360 25.220 ;
        RECT 61.040 25.200 61.950 25.680 ;
        RECT 40.020 24.730 40.920 25.200 ;
        RECT 65.350 25.190 66.260 25.670 ;
        RECT 79.330 25.180 80.240 25.650 ;
        RECT 88.480 25.490 88.720 25.875 ;
        RECT 87.740 25.250 88.720 25.490 ;
        RECT 87.740 24.710 88.060 25.250 ;
        RECT 48.160 22.510 48.500 24.010 ;
        RECT 85.810 23.990 86.710 24.470 ;
        RECT 49.670 22.490 50.570 22.970 ;
        RECT 59.140 22.480 60.050 22.960 ;
        RECT 68.150 22.470 69.060 22.950 ;
        RECT 77.800 22.440 78.710 22.920 ;
        RECT 30.410 16.460 31.770 16.930 ;
        RECT 121.260 15.690 121.560 66.150 ;
        RECT 10.960 15.360 30.990 15.690 ;
        RECT 31.160 15.390 121.560 15.690 ;
        RECT 10.960 9.410 11.300 15.360 ;
        RECT 30.400 13.760 31.500 14.210 ;
        RECT 12.700 11.210 13.600 11.680 ;
        RECT 21.670 11.180 22.570 11.650 ;
        RECT 30.770 11.160 31.670 11.630 ;
        RECT 39.960 11.140 40.860 11.610 ;
        RECT 49.020 11.130 49.920 11.600 ;
        RECT 58.100 11.120 59.000 11.590 ;
        RECT 67.670 11.090 68.570 11.560 ;
        RECT 77.350 11.080 78.250 11.550 ;
        RECT 81.530 9.330 81.880 15.390 ;
        RECT 12.690 8.500 13.590 8.970 ;
        RECT 21.670 8.460 22.570 8.930 ;
        RECT 30.950 8.450 31.850 8.920 ;
        RECT 39.970 8.420 40.870 8.890 ;
        RECT 49.230 8.410 50.130 8.880 ;
        RECT 58.080 8.390 58.980 8.860 ;
        RECT 67.520 8.370 68.420 8.840 ;
        RECT 77.260 8.360 78.160 8.830 ;
        RECT 151.150 3.190 152.710 4.310 ;
      LAYER met3 ;
        RECT 4.070 88.610 119.355 89.680 ;
        RECT 93.995 88.600 95.065 88.610 ;
        RECT 1.000 85.190 66.530 86.650 ;
        RECT 1.000 85.110 105.760 85.190 ;
        RECT 1.000 84.050 116.380 85.110 ;
        RECT 1.000 84.040 66.530 84.050 ;
        RECT 20.180 83.140 21.400 84.040 ;
        RECT 20.180 82.680 24.220 83.140 ;
        RECT 20.180 79.420 21.400 82.680 ;
        RECT 24.400 79.970 27.920 80.410 ;
        RECT 26.710 79.560 27.920 79.970 ;
        RECT 20.180 78.960 24.690 79.420 ;
        RECT 20.180 75.330 21.400 78.960 ;
        RECT 26.700 76.720 27.920 79.560 ;
        RECT 24.170 76.280 27.920 76.720 ;
        RECT 31.600 78.900 32.510 84.040 ;
        RECT 31.600 78.420 34.480 78.900 ;
        RECT 31.600 76.390 32.510 78.420 ;
        RECT 20.180 74.870 24.500 75.330 ;
        RECT 20.180 71.620 21.400 74.870 ;
        RECT 26.700 73.690 27.920 76.280 ;
        RECT 30.440 75.900 32.510 76.390 ;
        RECT 26.700 73.210 30.130 73.690 ;
        RECT 26.700 72.610 27.920 73.210 ;
        RECT 24.710 72.170 27.920 72.610 ;
        RECT 20.180 71.160 24.400 71.620 ;
        RECT 20.180 67.020 21.400 71.160 ;
        RECT 26.700 68.880 27.920 72.170 ;
        RECT 31.600 72.165 32.510 75.900 ;
        RECT 35.250 75.700 37.760 76.180 ;
        RECT 31.605 72.150 32.510 72.165 ;
        RECT 31.605 71.670 33.420 72.150 ;
        RECT 31.605 71.640 32.510 71.670 ;
        RECT 31.600 71.065 32.510 71.640 ;
        RECT 32.945 69.690 33.420 71.670 ;
        RECT 32.920 69.230 34.740 69.690 ;
        RECT 24.110 68.860 27.920 68.880 ;
        RECT 24.110 68.440 30.430 68.860 ;
        RECT 26.700 68.380 30.430 68.440 ;
        RECT 20.180 66.560 24.420 67.020 ;
        RECT 20.180 63.290 21.400 66.560 ;
        RECT 26.700 64.640 27.920 68.380 ;
        RECT 32.945 67.350 33.420 69.230 ;
        RECT 29.740 66.890 33.420 67.350 ;
        RECT 36.740 68.760 37.760 75.700 ;
        RECT 39.190 70.940 40.360 84.040 ;
        RECT 44.700 83.860 46.210 84.040 ;
        RECT 56.120 83.860 57.320 84.040 ;
        RECT 63.710 83.860 65.170 84.040 ;
        RECT 44.990 83.060 46.210 83.860 ;
        RECT 44.990 82.600 49.030 83.060 ;
        RECT 44.990 79.340 46.210 82.600 ;
        RECT 49.210 79.890 52.730 80.330 ;
        RECT 51.520 79.480 52.730 79.890 ;
        RECT 44.990 78.880 49.500 79.340 ;
        RECT 44.990 75.250 46.210 78.880 ;
        RECT 51.510 76.640 52.730 79.480 ;
        RECT 48.980 76.200 52.730 76.640 ;
        RECT 56.410 78.820 57.320 83.860 ;
        RECT 56.410 78.340 59.290 78.820 ;
        RECT 56.410 76.310 57.320 78.340 ;
        RECT 44.990 74.790 49.310 75.250 ;
        RECT 44.990 71.540 46.210 74.790 ;
        RECT 51.510 73.610 52.730 76.200 ;
        RECT 55.250 75.820 57.320 76.310 ;
        RECT 51.510 73.130 54.940 73.610 ;
        RECT 51.510 72.530 52.730 73.130 ;
        RECT 49.520 72.090 52.730 72.530 ;
        RECT 44.990 71.080 49.210 71.540 ;
        RECT 36.740 68.280 38.730 68.760 ;
        RECT 36.740 66.970 37.760 68.280 ;
        RECT 26.700 64.270 30.490 64.640 ;
        RECT 24.630 64.160 30.490 64.270 ;
        RECT 24.630 63.830 27.920 64.160 ;
        RECT 20.180 62.830 24.760 63.290 ;
        RECT 20.180 59.200 21.400 62.830 ;
        RECT 26.700 60.550 27.920 63.830 ;
        RECT 32.945 62.270 33.420 66.890 ;
        RECT 35.460 66.490 37.760 66.970 ;
        RECT 30.965 61.795 33.420 62.270 ;
        RECT 24.250 60.110 27.920 60.550 ;
        RECT 26.700 59.530 27.920 60.110 ;
        RECT 20.180 58.740 24.190 59.200 ;
        RECT 26.700 59.050 30.500 59.530 ;
        RECT 20.180 55.450 21.400 58.740 ;
        RECT 26.700 56.470 27.920 59.050 ;
        RECT 24.680 56.000 27.920 56.470 ;
        RECT 20.180 54.990 24.520 55.450 ;
        RECT 20.180 54.980 21.400 54.990 ;
        RECT 26.700 52.770 27.920 56.000 ;
        RECT 24.260 52.240 27.920 52.770 ;
        RECT 26.700 49.410 27.920 52.240 ;
        RECT 36.740 49.410 37.760 66.490 ;
        RECT 44.990 66.940 46.210 71.080 ;
        RECT 51.510 68.800 52.730 72.090 ;
        RECT 56.410 72.085 57.320 75.820 ;
        RECT 60.060 75.620 62.570 76.100 ;
        RECT 56.415 72.070 57.320 72.085 ;
        RECT 56.415 71.590 58.230 72.070 ;
        RECT 56.415 71.560 57.320 71.590 ;
        RECT 56.410 70.985 57.320 71.560 ;
        RECT 57.755 69.610 58.230 71.590 ;
        RECT 57.730 69.150 59.550 69.610 ;
        RECT 48.920 68.780 52.730 68.800 ;
        RECT 48.920 68.360 55.240 68.780 ;
        RECT 51.510 68.300 55.240 68.360 ;
        RECT 44.990 66.480 49.230 66.940 ;
        RECT 44.990 63.210 46.210 66.480 ;
        RECT 51.510 64.560 52.730 68.300 ;
        RECT 57.755 67.270 58.230 69.150 ;
        RECT 54.550 66.810 58.230 67.270 ;
        RECT 61.550 68.680 62.570 75.620 ;
        RECT 64.000 70.860 65.170 83.860 ;
        RECT 75.990 77.030 77.130 84.050 ;
        RECT 81.700 83.260 82.840 84.050 ;
        RECT 85.540 83.210 86.680 84.050 ;
        RECT 89.990 83.190 91.130 84.050 ;
        RECT 92.260 84.000 102.710 84.050 ;
        RECT 92.980 83.210 94.120 84.000 ;
        RECT 96.820 83.160 97.960 84.000 ;
        RECT 101.270 83.140 102.410 84.000 ;
        RECT 104.950 83.970 116.380 84.050 ;
        RECT 106.800 83.180 107.940 83.970 ;
        RECT 110.640 83.130 111.780 83.970 ;
        RECT 115.090 83.110 116.230 83.970 ;
        RECT 81.665 80.135 82.735 80.995 ;
        RECT 85.635 80.135 86.705 80.925 ;
        RECT 89.965 80.135 91.035 80.955 ;
        RECT 80.985 80.090 91.500 80.135 ;
        RECT 80.985 80.085 92.550 80.090 ;
        RECT 92.945 80.085 94.015 80.945 ;
        RECT 96.915 80.085 97.985 80.875 ;
        RECT 101.245 80.085 102.315 80.905 ;
        RECT 106.765 80.085 107.835 80.915 ;
        RECT 80.985 80.055 107.835 80.085 ;
        RECT 110.735 80.055 111.805 80.845 ;
        RECT 115.065 80.135 116.135 80.875 ;
        RECT 118.285 80.135 119.355 88.610 ;
        RECT 113.135 80.055 119.355 80.135 ;
        RECT 80.985 80.050 108.550 80.055 ;
        RECT 108.950 80.050 109.830 80.055 ;
        RECT 80.985 80.030 109.830 80.050 ;
        RECT 110.470 80.030 119.355 80.055 ;
        RECT 80.985 79.480 119.355 80.030 ;
        RECT 80.985 79.065 119.370 79.480 ;
        RECT 91.460 79.015 119.370 79.065 ;
        RECT 102.985 78.985 119.370 79.015 ;
        RECT 116.350 78.970 119.370 78.985 ;
        RECT 75.990 75.890 122.680 77.030 ;
        RECT 121.550 75.750 122.680 75.890 ;
        RECT 121.550 73.950 122.690 75.750 ;
        RECT 134.780 73.020 135.870 73.940 ;
        RECT 137.560 71.680 138.650 72.550 ;
        RECT 119.260 70.640 121.060 71.670 ;
        RECT 119.260 69.730 121.020 70.640 ;
        RECT 61.550 68.200 63.540 68.680 ;
        RECT 75.550 68.630 121.020 69.730 ;
        RECT 61.550 66.890 62.570 68.200 ;
        RECT 51.510 64.190 55.300 64.560 ;
        RECT 49.440 64.080 55.300 64.190 ;
        RECT 49.440 63.750 52.730 64.080 ;
        RECT 44.990 62.750 49.570 63.210 ;
        RECT 44.990 59.120 46.210 62.750 ;
        RECT 51.510 60.470 52.730 63.750 ;
        RECT 57.755 62.190 58.230 66.810 ;
        RECT 60.270 66.410 62.570 66.890 ;
        RECT 55.775 61.715 58.230 62.190 ;
        RECT 49.060 60.030 52.730 60.470 ;
        RECT 51.510 59.450 52.730 60.030 ;
        RECT 44.990 58.660 49.000 59.120 ;
        RECT 51.510 58.970 55.310 59.450 ;
        RECT 44.990 55.370 46.210 58.660 ;
        RECT 51.510 56.390 52.730 58.970 ;
        RECT 49.490 55.920 52.730 56.390 ;
        RECT 44.990 54.910 49.330 55.370 ;
        RECT 44.990 54.900 46.210 54.910 ;
        RECT 51.510 52.690 52.730 55.920 ;
        RECT 49.070 52.160 52.730 52.690 ;
        RECT 4.000 49.320 43.820 49.410 ;
        RECT 51.510 49.320 52.730 52.160 ;
        RECT 61.550 49.320 62.570 66.410 ;
        RECT 75.550 67.930 121.040 68.630 ;
        RECT 75.550 49.450 77.350 67.930 ;
        RECT 65.710 49.320 77.350 49.450 ;
        RECT 4.000 47.650 77.350 49.320 ;
        RECT 4.000 46.880 66.265 47.650 ;
        RECT 30.540 32.780 33.230 33.680 ;
        RECT 1.860 29.770 31.370 30.540 ;
        RECT 32.330 29.070 33.230 32.780 ;
        RECT 44.260 30.210 86.690 31.110 ;
        RECT 44.260 29.070 45.160 30.210 ;
        RECT 4.010 28.170 45.160 29.070 ;
        RECT 12.560 27.530 13.460 28.170 ;
        RECT 21.890 27.480 22.790 28.170 ;
        RECT 30.520 27.450 31.420 28.170 ;
        RECT 40.050 27.460 40.950 28.170 ;
        RECT 12.600 24.250 13.500 25.240 ;
        RECT 46.640 25.230 47.540 30.210 ;
        RECT 49.540 29.620 50.440 30.210 ;
        RECT 58.990 29.590 59.890 30.210 ;
        RECT 50.860 26.500 58.200 27.400 ;
        RECT 21.900 24.250 22.800 25.230 ;
        RECT 30.460 24.250 31.360 25.190 ;
        RECT 40.010 24.250 40.910 25.210 ;
        RECT 0.990 23.350 45.160 24.250 ;
        RECT 44.260 22.480 45.160 23.350 ;
        RECT 44.260 21.880 45.170 22.480 ;
        RECT 49.660 21.880 50.560 22.990 ;
        RECT 53.880 21.880 54.780 26.500 ;
        RECT 63.150 26.080 64.050 30.210 ;
        RECT 67.850 29.580 68.750 30.210 ;
        RECT 77.320 29.560 78.220 30.210 ;
        RECT 79.330 30.180 80.230 30.210 ;
        RECT 69.140 26.390 76.210 27.290 ;
        RECT 60.220 25.180 66.900 26.080 ;
        RECT 59.140 21.880 60.040 22.970 ;
        RECT 68.180 21.880 69.080 22.940 ;
        RECT 72.510 21.880 73.410 26.390 ;
        RECT 79.330 25.650 80.230 29.390 ;
        RECT 85.790 26.770 86.690 30.210 ;
        RECT 79.330 25.170 80.240 25.650 ;
        RECT 77.780 21.880 78.680 22.910 ;
        RECT 85.810 21.880 86.710 24.440 ;
        RECT 44.260 20.980 86.710 21.880 ;
        RECT 30.410 16.140 33.280 17.040 ;
        RECT 1.470 13.320 31.490 14.290 ;
        RECT 32.380 12.770 33.280 16.140 ;
        RECT 3.970 11.870 81.100 12.770 ;
        RECT 12.700 11.220 13.600 11.870 ;
        RECT 21.680 11.180 22.580 11.870 ;
        RECT 30.770 11.170 31.670 11.870 ;
        RECT 39.960 11.160 40.860 11.870 ;
        RECT 49.020 11.130 49.920 11.870 ;
        RECT 58.100 11.120 59.000 11.870 ;
        RECT 67.670 11.120 68.570 11.870 ;
        RECT 77.350 11.400 78.250 11.870 ;
        RECT 77.340 11.080 78.250 11.400 ;
        RECT 12.710 7.950 13.610 8.950 ;
        RECT 21.670 7.950 22.570 8.960 ;
        RECT 30.950 7.950 31.850 8.920 ;
        RECT 39.980 7.950 40.880 8.900 ;
        RECT 49.220 7.950 50.120 8.870 ;
        RECT 58.080 7.950 58.980 8.900 ;
        RECT 67.530 7.950 68.430 8.860 ;
        RECT 77.280 7.950 78.180 8.830 ;
        RECT 1.050 7.050 78.180 7.950 ;
        RECT 151.150 3.190 152.710 4.310 ;
      LAYER met4 ;
        RECT 135.550 73.940 135.850 224.760 ;
        RECT 134.780 73.020 135.870 73.940 ;
        RECT 138.310 72.550 138.610 224.760 ;
        RECT 137.560 71.680 138.650 72.550 ;
        RECT 151.150 3.190 152.710 4.310 ;
        RECT 151.810 1.000 152.710 3.190 ;
  END
END tt_um_ohmy90_adders
END LIBRARY

