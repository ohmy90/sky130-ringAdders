magic
tech sky130A
magscale 1 2
timestamp 1755109194
<< nwell >>
rect 18558 41910 18879 43548
rect 18542 40198 18863 41562
rect 18550 38770 18871 39766
rect 18564 37692 18885 38504
rect 18576 36726 18897 37350
rect 18584 36022 18905 36466
rect 18608 33162 18929 35078
rect 18608 30880 18929 32796
rect 18612 28634 18933 30550
rect 18604 26448 18925 28364
rect 18608 24202 18929 26118
rect 7632 23089 9548 23410
rect 9878 23093 11794 23414
rect 12064 23085 13980 23406
rect 14310 23089 16226 23410
rect 16592 23089 18508 23410
rect 9392 17212 9820 17533
rect 15443 17064 15881 17385
rect 16229 17102 16659 17423
rect 17095 17104 17533 17425
rect 17873 17094 18301 17415
rect 18989 17096 19423 17417
rect 19855 17098 20297 17419
rect 20625 17088 21065 17409
rect 21327 17086 21771 17407
rect 22111 17088 22553 17409
rect 22969 17078 23411 17399
rect 4338 16303 5150 16624
rect 9204 16307 10016 16628
rect 16208 16411 16650 16732
rect 17066 16401 17508 16722
rect 17848 16403 18292 16724
rect 18554 16401 18994 16722
rect 19322 16391 19764 16712
rect 20196 16393 20630 16714
rect 21318 16395 21746 16716
rect 22086 16385 22524 16706
rect 22960 16387 23390 16708
rect 4438 15559 5064 15880
rect 6570 15449 7382 15770
rect 9304 15563 9930 15884
rect 4348 14739 5160 15060
rect 5712 14949 6340 15270
rect 11436 15453 12248 15774
rect 9214 14743 10026 15064
rect 10578 14953 11206 15274
rect 23446 14549 25546 14870
rect 4448 13995 5074 14316
rect 5694 13983 6506 14304
rect 7684 13967 8404 14288
rect 9312 13999 9940 14320
rect 10560 13987 11372 14308
rect 12550 13971 13270 14292
rect 6756 13609 7380 13930
rect 11622 13613 12248 13934
rect 4340 13071 5152 13392
rect 5818 13141 6446 13462
rect 9206 13075 10018 13396
rect 10684 13145 11312 13466
rect 4440 12327 5066 12648
rect 5814 12121 6442 12442
rect 9304 12331 9932 12652
rect 10680 12125 11308 12446
rect 4350 11507 5162 11828
rect 9216 11511 10028 11832
rect 4448 10763 5076 11084
rect 9314 10767 9942 11088
rect 6074 6018 6508 6339
rect 9890 5386 11528 5707
rect 11950 5374 13590 5695
rect 13908 5382 15548 5703
rect 15904 5388 17542 5709
rect 1708 4966 3346 5287
rect 3842 4958 5480 5279
rect 5792 4958 7432 5279
rect 7794 4964 9434 5285
rect 10008 4512 11648 4833
rect 18264 4814 19260 5135
rect 12190 4468 13826 4789
rect 14190 4462 15828 4783
rect 16214 4444 17850 4765
rect 5956 2758 6396 3079
rect 1678 1706 3316 2027
rect 3748 1702 5386 2023
rect 5704 1702 7338 2023
rect 7702 1708 9340 2029
rect 9658 1708 11292 2029
rect 11646 1708 13284 2029
rect 13600 1708 15236 2029
rect 15662 1708 17300 2029
<< pwell >>
rect 18945 43421 19102 43507
rect 18937 42011 19119 43408
rect 18937 41977 19157 42011
rect 18937 41962 19119 41977
rect 18929 41435 19086 41521
rect 18921 40299 19103 41431
rect 18921 40270 19141 40299
rect 19107 40265 19141 40270
rect 18937 39639 19094 39725
rect 18929 38871 19111 39616
rect 18929 38842 19149 38871
rect 19115 38837 19149 38842
rect 18951 38377 19108 38463
rect 18943 37793 19125 38373
rect 18943 37759 19163 37793
rect 18943 37741 19125 37759
rect 18963 37223 19120 37309
rect 18955 36827 19137 37213
rect 18955 36793 19175 36827
rect 18955 36775 19137 36793
rect 18971 36339 19128 36425
rect 18963 36123 19145 36333
rect 18963 36089 19183 36123
rect 18963 36063 19145 36089
rect 18995 34951 19152 35037
rect 18987 34394 19169 34947
rect 19033 34086 19169 34394
rect 18989 33904 19169 34086
rect 19033 33263 19169 33904
rect 19033 33229 19207 33263
rect 19033 33201 19169 33229
rect 18995 32669 19152 32755
rect 18987 32112 19169 32665
rect 19033 31804 19169 32112
rect 18989 31622 19169 31804
rect 19033 30981 19169 31622
rect 19033 30947 19207 30981
rect 19033 30919 19169 30947
rect 18999 30423 19156 30509
rect 18991 29866 19173 30419
rect 19037 29558 19173 29866
rect 18993 29376 19173 29558
rect 19037 28735 19173 29376
rect 19037 28701 19211 28735
rect 19037 28673 19173 28701
rect 18991 28237 19148 28323
rect 18983 27680 19165 28233
rect 19029 27372 19165 27680
rect 18985 27190 19165 27372
rect 19029 26549 19165 27190
rect 19029 26515 19203 26549
rect 19029 26487 19165 26515
rect 18995 25991 19152 26077
rect 18987 25434 19169 25987
rect 19033 25126 19169 25434
rect 18989 24944 19169 25126
rect 19033 24303 19169 24944
rect 19033 24269 19207 24303
rect 19033 24241 19169 24269
rect 8374 22985 8556 23029
rect 8864 22985 9417 23031
rect 7671 22849 9417 22985
rect 9421 22866 9507 23023
rect 10620 22989 10802 23033
rect 11110 22989 11663 23035
rect 9917 22853 11663 22989
rect 11667 22870 11753 23027
rect 12806 22981 12988 23025
rect 13296 22981 13849 23027
rect 7699 22811 7733 22849
rect 9945 22815 9979 22853
rect 12103 22845 13849 22981
rect 13853 22862 13939 23019
rect 15052 22985 15234 23029
rect 15542 22985 16095 23031
rect 14349 22849 16095 22985
rect 16099 22866 16185 23023
rect 17334 22985 17516 23029
rect 17824 22985 18377 23031
rect 16631 22849 18377 22985
rect 18381 22866 18467 23023
rect 12131 22807 12165 22845
rect 14377 22811 14411 22849
rect 16659 22811 16693 22849
rect 9643 17777 9677 17811
rect 9643 17773 9664 17777
rect 9478 17591 9664 17773
rect 9693 17599 9779 17756
rect 16558 17667 16592 17701
rect 17432 17669 17466 17703
rect 16558 17663 16579 17667
rect 17432 17665 17453 17669
rect 15780 17629 15814 17663
rect 15780 17625 15801 17629
rect 15484 17451 15570 17608
rect 15615 17443 15801 17625
rect 16270 17489 16356 17646
rect 16393 17481 16579 17663
rect 17136 17491 17222 17648
rect 17267 17483 17453 17665
rect 18200 17659 18234 17693
rect 19322 17661 19356 17695
rect 20196 17663 20230 17697
rect 18200 17655 18221 17659
rect 19322 17657 19343 17661
rect 20196 17659 20217 17663
rect 17914 17481 18000 17638
rect 18035 17473 18221 17655
rect 19030 17483 19116 17640
rect 19157 17475 19343 17657
rect 19896 17485 19982 17642
rect 20031 17477 20217 17659
rect 20964 17653 20998 17687
rect 20964 17649 20985 17653
rect 20666 17475 20752 17632
rect 20799 17467 20985 17649
rect 21578 17651 21612 17685
rect 22452 17653 22486 17687
rect 21578 17647 21599 17651
rect 22452 17649 22473 17653
rect 21413 17465 21599 17647
rect 21644 17473 21730 17630
rect 22152 17475 22238 17632
rect 22287 17467 22473 17649
rect 23220 17643 23254 17677
rect 23220 17639 23241 17643
rect 23055 17457 23241 17639
rect 23284 17465 23370 17622
rect 4379 16080 4465 16237
rect 4477 16063 5111 16245
rect 9245 16084 9331 16241
rect 9343 16067 9977 16249
rect 16249 16188 16335 16345
rect 16378 16171 16564 16353
rect 16378 16167 16399 16171
rect 16365 16133 16399 16167
rect 17146 16161 17332 16343
rect 17381 16178 17467 16335
rect 17889 16180 17975 16337
rect 18020 16163 18206 16345
rect 17146 16157 17167 16161
rect 18020 16159 18041 16163
rect 17133 16123 17167 16157
rect 18007 16125 18041 16159
rect 18634 16161 18820 16343
rect 18867 16178 18953 16335
rect 18634 16157 18655 16161
rect 18621 16123 18655 16157
rect 19402 16151 19588 16333
rect 19637 16168 19723 16325
rect 20276 16153 20462 16335
rect 20503 16170 20589 16327
rect 21398 16155 21584 16337
rect 21619 16172 21705 16329
rect 19402 16147 19423 16151
rect 20276 16149 20297 16153
rect 21398 16151 21419 16155
rect 19389 16113 19423 16147
rect 20263 16115 20297 16149
rect 21385 16117 21419 16151
rect 22166 16145 22352 16327
rect 22397 16162 22483 16319
rect 23040 16147 23226 16329
rect 23263 16164 23349 16321
rect 22166 16141 22187 16145
rect 23040 16143 23061 16147
rect 22153 16107 22187 16141
rect 23027 16109 23061 16143
rect 4497 16025 4531 16063
rect 9363 16029 9397 16067
rect 4479 15336 4565 15493
rect 4795 15483 4985 15501
rect 4599 15319 4985 15483
rect 7024 15345 7251 15391
rect 4599 15315 4629 15319
rect 4595 15281 4629 15315
rect 6609 15209 7251 15345
rect 7255 15226 7341 15383
rect 9345 15340 9431 15497
rect 9661 15487 9851 15505
rect 9465 15323 9851 15487
rect 11890 15349 12117 15395
rect 9465 15319 9495 15323
rect 9461 15285 9495 15319
rect 6637 15171 6671 15209
rect 5979 14873 6169 14891
rect 5783 14709 6169 14873
rect 6213 14726 6299 14883
rect 11475 15213 12117 15349
rect 12121 15230 12207 15387
rect 11503 15175 11537 15213
rect 10845 14877 11035 14895
rect 10649 14713 11035 14877
rect 11079 14730 11165 14887
rect 10649 14709 10679 14713
rect 5783 14705 5813 14709
rect 4389 14516 4475 14673
rect 4487 14499 5121 14681
rect 5779 14671 5813 14705
rect 9255 14520 9341 14677
rect 9353 14503 9987 14685
rect 10645 14675 10679 14709
rect 4507 14461 4541 14499
rect 9373 14465 9407 14503
rect 24126 14488 24396 14495
rect 23938 14479 24396 14488
rect 23750 14445 24396 14479
rect 25011 14491 25195 14495
rect 25011 14445 25415 14491
rect 23485 14359 25415 14445
rect 23485 14352 24124 14359
rect 23485 14343 23936 14352
rect 23485 14309 23837 14343
rect 24396 14309 25415 14359
rect 25419 14326 25505 14483
rect 23513 14271 23547 14309
rect 4489 13772 4575 13929
rect 4805 13919 4995 13937
rect 4609 13755 4995 13919
rect 5735 13760 5821 13917
rect 6240 13879 6467 13925
rect 4609 13751 4639 13755
rect 4605 13717 4639 13751
rect 5825 13743 6467 13879
rect 5853 13705 5887 13743
rect 8084 13869 8273 13909
rect 7723 13733 8273 13869
rect 8277 13744 8363 13901
rect 9353 13776 9439 13933
rect 9671 13923 9861 13941
rect 9475 13759 9861 13923
rect 10601 13764 10687 13921
rect 11106 13883 11333 13929
rect 9475 13755 9505 13759
rect 7752 13689 7786 13733
rect 8084 13727 8273 13733
rect 9471 13721 9505 13755
rect 10691 13747 11333 13883
rect 10719 13709 10753 13747
rect 12950 13873 13139 13913
rect 12589 13737 13139 13873
rect 13143 13748 13229 13905
rect 12618 13693 12652 13737
rect 12950 13731 13139 13737
rect 7005 13505 7191 13551
rect 6824 13369 7191 13505
rect 7253 13386 7339 13543
rect 11871 13509 12057 13555
rect 6824 13365 6857 13369
rect 6823 13331 6857 13365
rect 4381 12848 4467 13005
rect 4479 12831 5113 13013
rect 5859 12918 5945 13075
rect 6223 13037 6407 13083
rect 11690 13373 12057 13509
rect 12121 13390 12207 13547
rect 11690 13369 11723 13373
rect 11689 13335 11723 13369
rect 5949 12901 6407 13037
rect 5977 12863 6011 12901
rect 9247 12852 9333 13009
rect 9345 12835 9979 13017
rect 10725 12922 10811 13079
rect 11089 13041 11273 13087
rect 10815 12905 11273 13041
rect 10843 12867 10877 12905
rect 4499 12793 4533 12831
rect 9365 12797 9399 12835
rect 4481 12104 4567 12261
rect 4797 12251 4987 12269
rect 4601 12087 4987 12251
rect 9345 12108 9431 12265
rect 9663 12255 9853 12273
rect 9467 12091 9853 12255
rect 9467 12087 9497 12091
rect 4601 12083 4631 12087
rect 4597 12049 4631 12083
rect 5855 11898 5941 12055
rect 6173 12045 6363 12063
rect 9463 12053 9497 12087
rect 5977 11881 6363 12045
rect 10721 11902 10807 12059
rect 11039 12049 11229 12067
rect 10843 11885 11229 12049
rect 10843 11881 10873 11885
rect 5977 11877 6007 11881
rect 5973 11843 6007 11877
rect 10839 11847 10873 11881
rect 4391 11284 4477 11441
rect 4489 11267 5123 11449
rect 9257 11288 9343 11445
rect 9355 11271 9989 11453
rect 4509 11229 4543 11267
rect 9375 11233 9409 11271
rect 4489 10540 4575 10697
rect 4807 10687 4997 10705
rect 4611 10523 4997 10687
rect 9355 10544 9441 10701
rect 9673 10691 9863 10709
rect 9477 10527 9863 10691
rect 9477 10523 9507 10527
rect 4611 10519 4641 10523
rect 4607 10485 4641 10519
rect 9473 10489 9507 10523
rect 6325 6583 6359 6617
rect 6325 6579 6346 6583
rect 6160 6397 6346 6579
rect 6381 6405 6467 6562
rect 11426 5947 11460 5985
rect 9931 5773 10017 5930
rect 10054 5811 11489 5947
rect 13488 5935 13522 5973
rect 15446 5943 15480 5981
rect 17440 5949 17474 5987
rect 10054 5765 10240 5811
rect 11303 5765 11489 5811
rect 11991 5761 12077 5918
rect 12116 5799 13551 5935
rect 12116 5753 12302 5799
rect 13365 5753 13551 5799
rect 13949 5769 14035 5926
rect 14074 5807 15509 5943
rect 14074 5761 14260 5807
rect 15323 5761 15509 5807
rect 15945 5775 16031 5932
rect 16068 5813 17503 5949
rect 16068 5767 16254 5813
rect 17317 5767 17503 5813
rect 3244 5527 3278 5565
rect 1749 5353 1835 5510
rect 1872 5391 3307 5527
rect 5378 5519 5412 5557
rect 7330 5519 7364 5557
rect 9332 5525 9366 5563
rect 1872 5345 2058 5391
rect 3121 5345 3307 5391
rect 3883 5345 3969 5502
rect 4006 5383 5441 5519
rect 4006 5337 4192 5383
rect 5255 5337 5441 5383
rect 5833 5345 5919 5502
rect 5958 5383 7393 5519
rect 5958 5337 6144 5383
rect 7207 5337 7393 5383
rect 7835 5351 7921 5508
rect 7960 5389 9395 5525
rect 7960 5343 8146 5389
rect 9209 5343 9395 5389
rect 19012 5375 19046 5413
rect 18349 5239 19129 5375
rect 18943 5193 19129 5239
rect 19133 5201 19219 5358
rect 11454 5073 11488 5111
rect 10082 4937 11517 5073
rect 10082 4891 10268 4937
rect 11331 4891 11517 4937
rect 11521 4899 11607 5056
rect 13724 5029 13758 5067
rect 12231 4855 12317 5012
rect 12352 4893 13787 5029
rect 15726 5023 15760 5061
rect 12352 4847 12538 4893
rect 13601 4847 13787 4893
rect 14231 4849 14317 5006
rect 14354 4887 15789 5023
rect 17748 5005 17782 5043
rect 14354 4841 14540 4887
rect 15603 4841 15789 4887
rect 16255 4831 16341 4988
rect 16376 4869 17811 5005
rect 16376 4823 16562 4869
rect 17625 4823 17811 4869
rect 6295 3323 6329 3357
rect 6295 3319 6316 3323
rect 5997 3145 6083 3302
rect 6130 3137 6316 3319
rect 3214 2267 3248 2305
rect 1719 2093 1805 2250
rect 1842 2131 3277 2267
rect 5284 2263 5318 2301
rect 7236 2263 7270 2301
rect 9238 2269 9272 2307
rect 11190 2269 11224 2307
rect 13182 2269 13216 2307
rect 15134 2269 15168 2307
rect 17198 2269 17232 2307
rect 1842 2085 2028 2131
rect 3091 2085 3277 2131
rect 3789 2089 3875 2246
rect 3912 2127 5347 2263
rect 3912 2081 4098 2127
rect 5161 2081 5347 2127
rect 5745 2089 5831 2246
rect 5864 2127 7299 2263
rect 5864 2081 6050 2127
rect 7113 2081 7299 2127
rect 7743 2095 7829 2252
rect 7866 2133 9301 2269
rect 7866 2087 8052 2133
rect 9115 2087 9301 2133
rect 9699 2095 9785 2252
rect 9818 2133 11253 2269
rect 9818 2087 10004 2133
rect 11067 2087 11253 2133
rect 11687 2095 11773 2252
rect 11810 2133 13245 2269
rect 11810 2087 11996 2133
rect 13059 2087 13245 2133
rect 13641 2095 13727 2252
rect 13762 2133 15197 2269
rect 13762 2087 13948 2133
rect 15011 2087 15197 2133
rect 15703 2095 15789 2252
rect 15826 2133 17261 2269
rect 15826 2087 16012 2133
rect 17075 2087 17261 2133
<< scnmos >>
rect 18963 43300 19093 43330
rect 18963 43216 19093 43246
rect 18963 43132 19093 43162
rect 18963 43048 19093 43078
rect 18963 42964 19093 42994
rect 18963 42880 19093 42910
rect 18963 42796 19093 42826
rect 18963 42712 19093 42742
rect 18963 42628 19093 42658
rect 18963 42544 19093 42574
rect 18963 42460 19093 42490
rect 18963 42376 19093 42406
rect 18963 42292 19093 42322
rect 18963 42208 19093 42238
rect 18963 42124 19093 42154
rect 18963 42040 19093 42070
rect 18947 41272 19077 41302
rect 18947 41188 19077 41218
rect 18947 41104 19077 41134
rect 18947 41020 19077 41050
rect 18947 40936 19077 40966
rect 18947 40852 19077 40882
rect 18947 40768 19077 40798
rect 18947 40684 19077 40714
rect 18947 40600 19077 40630
rect 18947 40516 19077 40546
rect 18947 40432 19077 40462
rect 18947 40348 19077 40378
rect 18955 39508 19085 39538
rect 18955 39424 19085 39454
rect 18955 39340 19085 39370
rect 18955 39256 19085 39286
rect 18955 39172 19085 39202
rect 18955 39088 19085 39118
rect 18955 39004 19085 39034
rect 18955 38920 19085 38950
rect 18969 38263 19099 38293
rect 18969 38179 19099 38209
rect 18969 38095 19099 38125
rect 18969 38011 19099 38041
rect 18969 37927 19099 37957
rect 18969 37843 19099 37873
rect 18981 37105 19111 37135
rect 18981 37021 19111 37051
rect 18981 36937 19111 36967
rect 18981 36853 19111 36883
rect 18989 36225 19119 36255
rect 18989 36141 19119 36171
rect 19013 34839 19143 34869
rect 19059 34744 19143 34774
rect 19013 34556 19143 34586
rect 19013 34472 19143 34502
rect 19059 34282 19143 34312
rect 19071 34187 19143 34217
rect 19071 34081 19143 34111
rect 19015 33980 19143 34010
rect 19059 33861 19143 33891
rect 19071 33762 19143 33792
rect 19071 33663 19143 33693
rect 19059 33551 19143 33581
rect 19059 33363 19143 33393
rect 19059 33279 19143 33309
rect 19013 32557 19143 32587
rect 19059 32462 19143 32492
rect 19013 32274 19143 32304
rect 19013 32190 19143 32220
rect 19059 32000 19143 32030
rect 19071 31905 19143 31935
rect 19071 31799 19143 31829
rect 19015 31698 19143 31728
rect 19059 31579 19143 31609
rect 19071 31480 19143 31510
rect 19071 31381 19143 31411
rect 19059 31269 19143 31299
rect 19059 31081 19143 31111
rect 19059 30997 19143 31027
rect 19017 30311 19147 30341
rect 19063 30216 19147 30246
rect 19017 30028 19147 30058
rect 19017 29944 19147 29974
rect 19063 29754 19147 29784
rect 19075 29659 19147 29689
rect 19075 29553 19147 29583
rect 19019 29452 19147 29482
rect 19063 29333 19147 29363
rect 19075 29234 19147 29264
rect 19075 29135 19147 29165
rect 19063 29023 19147 29053
rect 19063 28835 19147 28865
rect 19063 28751 19147 28781
rect 19009 28125 19139 28155
rect 19055 28030 19139 28060
rect 19009 27842 19139 27872
rect 19009 27758 19139 27788
rect 19055 27568 19139 27598
rect 19067 27473 19139 27503
rect 19067 27367 19139 27397
rect 19011 27266 19139 27296
rect 19055 27147 19139 27177
rect 19067 27048 19139 27078
rect 19067 26949 19139 26979
rect 19055 26837 19139 26867
rect 19055 26649 19139 26679
rect 19055 26565 19139 26595
rect 19013 25879 19143 25909
rect 19059 25784 19143 25814
rect 19013 25596 19143 25626
rect 19013 25512 19143 25542
rect 19059 25322 19143 25352
rect 19071 25227 19143 25257
rect 19071 25121 19143 25151
rect 19015 25020 19143 25050
rect 19059 24901 19143 24931
rect 19071 24802 19143 24832
rect 19071 24703 19143 24733
rect 19059 24591 19143 24621
rect 19059 24403 19143 24433
rect 19059 24319 19143 24349
rect 7749 22875 7779 22959
rect 7833 22875 7863 22959
rect 8021 22875 8051 22959
rect 8133 22875 8163 22947
rect 8232 22875 8262 22947
rect 8331 22875 8361 22959
rect 8450 22875 8480 23003
rect 8551 22875 8581 22947
rect 8657 22875 8687 22947
rect 8752 22875 8782 22959
rect 8942 22875 8972 23005
rect 9026 22875 9056 23005
rect 9214 22875 9244 22959
rect 9309 22875 9339 23005
rect 9995 22879 10025 22963
rect 10079 22879 10109 22963
rect 10267 22879 10297 22963
rect 10379 22879 10409 22951
rect 10478 22879 10508 22951
rect 10577 22879 10607 22963
rect 10696 22879 10726 23007
rect 10797 22879 10827 22951
rect 10903 22879 10933 22951
rect 10998 22879 11028 22963
rect 11188 22879 11218 23009
rect 11272 22879 11302 23009
rect 11460 22879 11490 22963
rect 11555 22879 11585 23009
rect 12181 22871 12211 22955
rect 12265 22871 12295 22955
rect 12453 22871 12483 22955
rect 12565 22871 12595 22943
rect 12664 22871 12694 22943
rect 12763 22871 12793 22955
rect 12882 22871 12912 22999
rect 12983 22871 13013 22943
rect 13089 22871 13119 22943
rect 13184 22871 13214 22955
rect 13374 22871 13404 23001
rect 13458 22871 13488 23001
rect 13646 22871 13676 22955
rect 13741 22871 13771 23001
rect 14427 22875 14457 22959
rect 14511 22875 14541 22959
rect 14699 22875 14729 22959
rect 14811 22875 14841 22947
rect 14910 22875 14940 22947
rect 15009 22875 15039 22959
rect 15128 22875 15158 23003
rect 15229 22875 15259 22947
rect 15335 22875 15365 22947
rect 15430 22875 15460 22959
rect 15620 22875 15650 23005
rect 15704 22875 15734 23005
rect 15892 22875 15922 22959
rect 15987 22875 16017 23005
rect 16709 22875 16739 22959
rect 16793 22875 16823 22959
rect 16981 22875 17011 22959
rect 17093 22875 17123 22947
rect 17192 22875 17222 22947
rect 17291 22875 17321 22959
rect 17410 22875 17440 23003
rect 17511 22875 17541 22947
rect 17617 22875 17647 22947
rect 17712 22875 17742 22959
rect 17902 22875 17932 23005
rect 17986 22875 18016 23005
rect 18174 22875 18204 22959
rect 18269 22875 18299 23005
rect 9556 17617 9586 17747
rect 15693 17469 15723 17599
rect 16471 17507 16501 17637
rect 17345 17509 17375 17639
rect 18113 17499 18143 17629
rect 19235 17501 19265 17631
rect 20109 17503 20139 17633
rect 20877 17493 20907 17623
rect 21491 17491 21521 17621
rect 22365 17493 22395 17623
rect 23133 17483 23163 17613
rect 4555 16089 4585 16219
rect 4639 16089 4669 16219
rect 4723 16089 4753 16219
rect 4807 16089 4837 16219
rect 4991 16089 5021 16219
rect 9421 16093 9451 16223
rect 9505 16093 9535 16223
rect 9589 16093 9619 16223
rect 9673 16093 9703 16223
rect 9857 16093 9887 16223
rect 16456 16197 16486 16327
rect 17224 16187 17254 16317
rect 18098 16189 18128 16319
rect 18712 16187 18742 16317
rect 19480 16177 19510 16307
rect 20354 16179 20384 16309
rect 21476 16181 21506 16311
rect 22244 16171 22274 16301
rect 23118 16173 23148 16303
rect 4681 15373 4711 15457
rect 4765 15373 4795 15457
rect 4873 15345 4903 15475
rect 9547 15377 9577 15461
rect 9631 15377 9661 15461
rect 6687 15235 6717 15319
rect 6775 15235 6805 15319
rect 6881 15235 6911 15319
rect 6977 15235 7007 15319
rect 7143 15235 7173 15365
rect 9739 15349 9769 15479
rect 11553 15239 11583 15323
rect 11641 15239 11671 15323
rect 11747 15239 11777 15323
rect 11843 15239 11873 15323
rect 12009 15239 12039 15369
rect 5865 14763 5895 14847
rect 5949 14763 5979 14847
rect 6057 14735 6087 14865
rect 10731 14767 10761 14851
rect 10815 14767 10845 14851
rect 10923 14739 10953 14869
rect 4565 14525 4595 14655
rect 4649 14525 4679 14655
rect 4733 14525 4763 14655
rect 4817 14525 4847 14655
rect 5001 14525 5031 14655
rect 9431 14529 9461 14659
rect 9515 14529 9545 14659
rect 9599 14529 9629 14659
rect 9683 14529 9713 14659
rect 9867 14529 9897 14659
rect 23563 14335 23593 14419
rect 23647 14335 23677 14419
rect 23731 14335 23761 14419
rect 23828 14369 23858 14453
rect 24016 14378 24046 14462
rect 24204 14385 24234 14469
rect 24288 14385 24318 14469
rect 24474 14335 24504 14419
rect 24558 14335 24588 14419
rect 24746 14335 24776 14419
rect 24934 14335 24964 14419
rect 25087 14385 25117 14469
rect 25307 14335 25337 14465
rect 4691 13809 4721 13893
rect 4775 13809 4805 13893
rect 4883 13781 4913 13911
rect 5903 13769 5933 13853
rect 5991 13769 6021 13853
rect 6097 13769 6127 13853
rect 6193 13769 6223 13853
rect 6359 13769 6389 13899
rect 7801 13759 7831 13843
rect 7897 13759 7927 13843
rect 7981 13759 8011 13843
rect 8065 13759 8095 13843
rect 8163 13753 8193 13883
rect 9557 13813 9587 13897
rect 9641 13813 9671 13897
rect 9749 13785 9779 13915
rect 10769 13773 10799 13857
rect 10857 13773 10887 13857
rect 10963 13773 10993 13857
rect 11059 13773 11089 13857
rect 11225 13773 11255 13903
rect 12667 13763 12697 13847
rect 12763 13763 12793 13847
rect 12847 13763 12877 13847
rect 12931 13763 12961 13847
rect 13029 13757 13059 13887
rect 6902 13395 6932 13479
rect 6986 13395 7016 13479
rect 7083 13395 7113 13525
rect 11768 13399 11798 13483
rect 11852 13399 11882 13483
rect 11949 13399 11979 13529
rect 4557 12857 4587 12987
rect 4641 12857 4671 12987
rect 4725 12857 4755 12987
rect 4809 12857 4839 12987
rect 4993 12857 5023 12987
rect 6027 12927 6057 13011
rect 6099 12927 6129 13011
rect 6171 12927 6201 13011
rect 6299 12927 6329 13057
rect 9423 12861 9453 12991
rect 9507 12861 9537 12991
rect 9591 12861 9621 12991
rect 9675 12861 9705 12991
rect 9859 12861 9889 12991
rect 10893 12931 10923 13015
rect 10965 12931 10995 13015
rect 11037 12931 11067 13015
rect 11165 12931 11195 13061
rect 4683 12141 4713 12225
rect 4767 12141 4797 12225
rect 4875 12113 4905 12243
rect 9549 12145 9579 12229
rect 9633 12145 9663 12229
rect 9741 12117 9771 12247
rect 6059 11935 6089 12019
rect 6143 11935 6173 12019
rect 6251 11907 6281 12037
rect 10925 11939 10955 12023
rect 11009 11939 11039 12023
rect 11117 11911 11147 12041
rect 4567 11293 4597 11423
rect 4651 11293 4681 11423
rect 4735 11293 4765 11423
rect 4819 11293 4849 11423
rect 5003 11293 5033 11423
rect 9433 11297 9463 11427
rect 9517 11297 9547 11427
rect 9601 11297 9631 11427
rect 9685 11297 9715 11427
rect 9869 11297 9899 11427
rect 4693 10577 4723 10661
rect 4777 10577 4807 10661
rect 4885 10549 4915 10679
rect 9559 10581 9589 10665
rect 9643 10581 9673 10665
rect 9751 10553 9781 10683
rect 6238 6423 6268 6553
rect 10132 5791 10162 5921
rect 10231 5837 10261 5921
rect 10327 5837 10357 5921
rect 10399 5837 10429 5921
rect 10495 5837 10525 5921
rect 10584 5837 10614 5921
rect 10668 5837 10698 5921
rect 10752 5837 10782 5921
rect 10940 5837 10970 5921
rect 11024 5837 11054 5921
rect 11108 5837 11138 5921
rect 11192 5837 11222 5921
rect 11282 5837 11312 5921
rect 1950 5371 1980 5501
rect 2049 5417 2079 5501
rect 2145 5417 2175 5501
rect 2217 5417 2247 5501
rect 2313 5417 2343 5501
rect 2402 5417 2432 5501
rect 2486 5417 2516 5501
rect 2570 5417 2600 5501
rect 2758 5417 2788 5501
rect 2842 5417 2872 5501
rect 2926 5417 2956 5501
rect 3010 5417 3040 5501
rect 3100 5417 3130 5501
rect 3199 5371 3229 5501
rect 4084 5363 4114 5493
rect 4183 5409 4213 5493
rect 4279 5409 4309 5493
rect 4351 5409 4381 5493
rect 4447 5409 4477 5493
rect 4536 5409 4566 5493
rect 4620 5409 4650 5493
rect 4704 5409 4734 5493
rect 4892 5409 4922 5493
rect 4976 5409 5006 5493
rect 5060 5409 5090 5493
rect 5144 5409 5174 5493
rect 5234 5409 5264 5493
rect 5333 5363 5363 5493
rect 6036 5363 6066 5493
rect 6135 5409 6165 5493
rect 6231 5409 6261 5493
rect 6303 5409 6333 5493
rect 6399 5409 6429 5493
rect 6488 5409 6518 5493
rect 6572 5409 6602 5493
rect 6656 5409 6686 5493
rect 6844 5409 6874 5493
rect 6928 5409 6958 5493
rect 7012 5409 7042 5493
rect 7096 5409 7126 5493
rect 7186 5409 7216 5493
rect 7285 5363 7315 5493
rect 8038 5369 8068 5499
rect 8137 5415 8167 5499
rect 8233 5415 8263 5499
rect 8305 5415 8335 5499
rect 8401 5415 8431 5499
rect 8490 5415 8520 5499
rect 8574 5415 8604 5499
rect 8658 5415 8688 5499
rect 8846 5415 8876 5499
rect 8930 5415 8960 5499
rect 9014 5415 9044 5499
rect 9098 5415 9128 5499
rect 9188 5415 9218 5499
rect 9287 5369 9317 5499
rect 11381 5791 11411 5921
rect 12194 5779 12224 5909
rect 12293 5825 12323 5909
rect 12389 5825 12419 5909
rect 12461 5825 12491 5909
rect 12557 5825 12587 5909
rect 12646 5825 12676 5909
rect 12730 5825 12760 5909
rect 12814 5825 12844 5909
rect 13002 5825 13032 5909
rect 13086 5825 13116 5909
rect 13170 5825 13200 5909
rect 13254 5825 13284 5909
rect 13344 5825 13374 5909
rect 13443 5779 13473 5909
rect 14152 5787 14182 5917
rect 14251 5833 14281 5917
rect 14347 5833 14377 5917
rect 14419 5833 14449 5917
rect 14515 5833 14545 5917
rect 14604 5833 14634 5917
rect 14688 5833 14718 5917
rect 14772 5833 14802 5917
rect 14960 5833 14990 5917
rect 15044 5833 15074 5917
rect 15128 5833 15158 5917
rect 15212 5833 15242 5917
rect 15302 5833 15332 5917
rect 15401 5787 15431 5917
rect 16146 5793 16176 5923
rect 16245 5839 16275 5923
rect 16341 5839 16371 5923
rect 16413 5839 16443 5923
rect 16509 5839 16539 5923
rect 16598 5839 16628 5923
rect 16682 5839 16712 5923
rect 16766 5839 16796 5923
rect 16954 5839 16984 5923
rect 17038 5839 17068 5923
rect 17122 5839 17152 5923
rect 17206 5839 17236 5923
rect 17296 5839 17326 5923
rect 17395 5793 17425 5923
rect 18427 5265 18457 5349
rect 18595 5265 18625 5349
rect 18691 5265 18721 5349
rect 18816 5265 18846 5349
rect 18912 5265 18942 5349
rect 10160 4917 10190 5047
rect 10259 4963 10289 5047
rect 10355 4963 10385 5047
rect 10427 4963 10457 5047
rect 10523 4963 10553 5047
rect 10612 4963 10642 5047
rect 10696 4963 10726 5047
rect 10780 4963 10810 5047
rect 10968 4963 10998 5047
rect 11052 4963 11082 5047
rect 11136 4963 11166 5047
rect 11220 4963 11250 5047
rect 11310 4963 11340 5047
rect 11409 4917 11439 5047
rect 12430 4873 12460 5003
rect 12529 4919 12559 5003
rect 12625 4919 12655 5003
rect 12697 4919 12727 5003
rect 12793 4919 12823 5003
rect 12882 4919 12912 5003
rect 12966 4919 12996 5003
rect 13050 4919 13080 5003
rect 13238 4919 13268 5003
rect 13322 4919 13352 5003
rect 13406 4919 13436 5003
rect 13490 4919 13520 5003
rect 13580 4919 13610 5003
rect 13679 4873 13709 5003
rect 19021 5219 19051 5349
rect 14432 4867 14462 4997
rect 14531 4913 14561 4997
rect 14627 4913 14657 4997
rect 14699 4913 14729 4997
rect 14795 4913 14825 4997
rect 14884 4913 14914 4997
rect 14968 4913 14998 4997
rect 15052 4913 15082 4997
rect 15240 4913 15270 4997
rect 15324 4913 15354 4997
rect 15408 4913 15438 4997
rect 15492 4913 15522 4997
rect 15582 4913 15612 4997
rect 15681 4867 15711 4997
rect 16454 4849 16484 4979
rect 16553 4895 16583 4979
rect 16649 4895 16679 4979
rect 16721 4895 16751 4979
rect 16817 4895 16847 4979
rect 16906 4895 16936 4979
rect 16990 4895 17020 4979
rect 17074 4895 17104 4979
rect 17262 4895 17292 4979
rect 17346 4895 17376 4979
rect 17430 4895 17460 4979
rect 17514 4895 17544 4979
rect 17604 4895 17634 4979
rect 17703 4849 17733 4979
rect 6208 3163 6238 3293
rect 1920 2111 1950 2241
rect 2019 2157 2049 2241
rect 2115 2157 2145 2241
rect 2187 2157 2217 2241
rect 2283 2157 2313 2241
rect 2372 2157 2402 2241
rect 2456 2157 2486 2241
rect 2540 2157 2570 2241
rect 2728 2157 2758 2241
rect 2812 2157 2842 2241
rect 2896 2157 2926 2241
rect 2980 2157 3010 2241
rect 3070 2157 3100 2241
rect 3169 2111 3199 2241
rect 3990 2107 4020 2237
rect 4089 2153 4119 2237
rect 4185 2153 4215 2237
rect 4257 2153 4287 2237
rect 4353 2153 4383 2237
rect 4442 2153 4472 2237
rect 4526 2153 4556 2237
rect 4610 2153 4640 2237
rect 4798 2153 4828 2237
rect 4882 2153 4912 2237
rect 4966 2153 4996 2237
rect 5050 2153 5080 2237
rect 5140 2153 5170 2237
rect 5239 2107 5269 2237
rect 5942 2107 5972 2237
rect 6041 2153 6071 2237
rect 6137 2153 6167 2237
rect 6209 2153 6239 2237
rect 6305 2153 6335 2237
rect 6394 2153 6424 2237
rect 6478 2153 6508 2237
rect 6562 2153 6592 2237
rect 6750 2153 6780 2237
rect 6834 2153 6864 2237
rect 6918 2153 6948 2237
rect 7002 2153 7032 2237
rect 7092 2153 7122 2237
rect 7191 2107 7221 2237
rect 7944 2113 7974 2243
rect 8043 2159 8073 2243
rect 8139 2159 8169 2243
rect 8211 2159 8241 2243
rect 8307 2159 8337 2243
rect 8396 2159 8426 2243
rect 8480 2159 8510 2243
rect 8564 2159 8594 2243
rect 8752 2159 8782 2243
rect 8836 2159 8866 2243
rect 8920 2159 8950 2243
rect 9004 2159 9034 2243
rect 9094 2159 9124 2243
rect 9193 2113 9223 2243
rect 9896 2113 9926 2243
rect 9995 2159 10025 2243
rect 10091 2159 10121 2243
rect 10163 2159 10193 2243
rect 10259 2159 10289 2243
rect 10348 2159 10378 2243
rect 10432 2159 10462 2243
rect 10516 2159 10546 2243
rect 10704 2159 10734 2243
rect 10788 2159 10818 2243
rect 10872 2159 10902 2243
rect 10956 2159 10986 2243
rect 11046 2159 11076 2243
rect 11145 2113 11175 2243
rect 11888 2113 11918 2243
rect 11987 2159 12017 2243
rect 12083 2159 12113 2243
rect 12155 2159 12185 2243
rect 12251 2159 12281 2243
rect 12340 2159 12370 2243
rect 12424 2159 12454 2243
rect 12508 2159 12538 2243
rect 12696 2159 12726 2243
rect 12780 2159 12810 2243
rect 12864 2159 12894 2243
rect 12948 2159 12978 2243
rect 13038 2159 13068 2243
rect 13137 2113 13167 2243
rect 13840 2113 13870 2243
rect 13939 2159 13969 2243
rect 14035 2159 14065 2243
rect 14107 2159 14137 2243
rect 14203 2159 14233 2243
rect 14292 2159 14322 2243
rect 14376 2159 14406 2243
rect 14460 2159 14490 2243
rect 14648 2159 14678 2243
rect 14732 2159 14762 2243
rect 14816 2159 14846 2243
rect 14900 2159 14930 2243
rect 14990 2159 15020 2243
rect 15089 2113 15119 2243
rect 15904 2113 15934 2243
rect 16003 2159 16033 2243
rect 16099 2159 16129 2243
rect 16171 2159 16201 2243
rect 16267 2159 16297 2243
rect 16356 2159 16386 2243
rect 16440 2159 16470 2243
rect 16524 2159 16554 2243
rect 16712 2159 16742 2243
rect 16796 2159 16826 2243
rect 16880 2159 16910 2243
rect 16964 2159 16994 2243
rect 17054 2159 17084 2243
rect 17153 2113 17183 2243
<< scpmoshvt >>
rect 18643 43300 18843 43330
rect 18643 43216 18843 43246
rect 18643 43132 18843 43162
rect 18643 43048 18843 43078
rect 18643 42964 18843 42994
rect 18643 42880 18843 42910
rect 18643 42796 18843 42826
rect 18643 42712 18843 42742
rect 18643 42628 18843 42658
rect 18643 42544 18843 42574
rect 18643 42460 18843 42490
rect 18643 42376 18843 42406
rect 18643 42292 18843 42322
rect 18643 42208 18843 42238
rect 18643 42124 18843 42154
rect 18643 42040 18843 42070
rect 18627 41272 18827 41302
rect 18627 41188 18827 41218
rect 18627 41104 18827 41134
rect 18627 41020 18827 41050
rect 18627 40936 18827 40966
rect 18627 40852 18827 40882
rect 18627 40768 18827 40798
rect 18627 40684 18827 40714
rect 18627 40600 18827 40630
rect 18627 40516 18827 40546
rect 18627 40432 18827 40462
rect 18627 40348 18827 40378
rect 18635 39508 18835 39538
rect 18635 39424 18835 39454
rect 18635 39340 18835 39370
rect 18635 39256 18835 39286
rect 18635 39172 18835 39202
rect 18635 39088 18835 39118
rect 18635 39004 18835 39034
rect 18635 38920 18835 38950
rect 18649 38263 18849 38293
rect 18649 38179 18849 38209
rect 18649 38095 18849 38125
rect 18649 38011 18849 38041
rect 18649 37927 18849 37957
rect 18649 37843 18849 37873
rect 18661 37105 18861 37135
rect 18661 37021 18861 37051
rect 18661 36937 18861 36967
rect 18661 36853 18861 36883
rect 18669 36225 18869 36255
rect 18669 36141 18869 36171
rect 18693 34839 18893 34869
rect 18693 34742 18821 34772
rect 18693 34554 18893 34584
rect 18693 34470 18893 34500
rect 18693 34259 18777 34289
rect 18693 34145 18777 34175
rect 18693 34061 18777 34091
rect 18693 33966 18843 33996
rect 18693 33834 18777 33864
rect 18693 33731 18777 33761
rect 18693 33636 18777 33666
rect 18693 33551 18777 33581
rect 18699 33363 18827 33393
rect 18699 33279 18827 33309
rect 18693 32557 18893 32587
rect 18693 32460 18821 32490
rect 18693 32272 18893 32302
rect 18693 32188 18893 32218
rect 18693 31977 18777 32007
rect 18693 31863 18777 31893
rect 18693 31779 18777 31809
rect 18693 31684 18843 31714
rect 18693 31552 18777 31582
rect 18693 31449 18777 31479
rect 18693 31354 18777 31384
rect 18693 31269 18777 31299
rect 18699 31081 18827 31111
rect 18699 30997 18827 31027
rect 18697 30311 18897 30341
rect 18697 30214 18825 30244
rect 18697 30026 18897 30056
rect 18697 29942 18897 29972
rect 18697 29731 18781 29761
rect 18697 29617 18781 29647
rect 18697 29533 18781 29563
rect 18697 29438 18847 29468
rect 18697 29306 18781 29336
rect 18697 29203 18781 29233
rect 18697 29108 18781 29138
rect 18697 29023 18781 29053
rect 18703 28835 18831 28865
rect 18703 28751 18831 28781
rect 18689 28125 18889 28155
rect 18689 28028 18817 28058
rect 18689 27840 18889 27870
rect 18689 27756 18889 27786
rect 18689 27545 18773 27575
rect 18689 27431 18773 27461
rect 18689 27347 18773 27377
rect 18689 27252 18839 27282
rect 18689 27120 18773 27150
rect 18689 27017 18773 27047
rect 18689 26922 18773 26952
rect 18689 26837 18773 26867
rect 18695 26649 18823 26679
rect 18695 26565 18823 26595
rect 18693 25879 18893 25909
rect 18693 25782 18821 25812
rect 18693 25594 18893 25624
rect 18693 25510 18893 25540
rect 18693 25299 18777 25329
rect 18693 25185 18777 25215
rect 18693 25101 18777 25131
rect 18693 25006 18843 25036
rect 18693 24874 18777 24904
rect 18693 24771 18777 24801
rect 18693 24676 18777 24706
rect 18693 24591 18777 24621
rect 18699 24403 18827 24433
rect 18699 24319 18827 24349
rect 7749 23191 7779 23319
rect 7833 23191 7863 23319
rect 8021 23241 8051 23325
rect 8106 23241 8136 23325
rect 8201 23241 8231 23325
rect 8304 23241 8334 23325
rect 8436 23175 8466 23325
rect 8531 23241 8561 23325
rect 8615 23241 8645 23325
rect 8729 23241 8759 23325
rect 8940 23125 8970 23325
rect 9024 23125 9054 23325
rect 9212 23197 9242 23325
rect 9309 23125 9339 23325
rect 9995 23195 10025 23323
rect 10079 23195 10109 23323
rect 10267 23245 10297 23329
rect 10352 23245 10382 23329
rect 10447 23245 10477 23329
rect 10550 23245 10580 23329
rect 10682 23179 10712 23329
rect 10777 23245 10807 23329
rect 10861 23245 10891 23329
rect 10975 23245 11005 23329
rect 11186 23129 11216 23329
rect 11270 23129 11300 23329
rect 11458 23201 11488 23329
rect 11555 23129 11585 23329
rect 12181 23187 12211 23315
rect 12265 23187 12295 23315
rect 12453 23237 12483 23321
rect 12538 23237 12568 23321
rect 12633 23237 12663 23321
rect 12736 23237 12766 23321
rect 12868 23171 12898 23321
rect 12963 23237 12993 23321
rect 13047 23237 13077 23321
rect 13161 23237 13191 23321
rect 13372 23121 13402 23321
rect 13456 23121 13486 23321
rect 13644 23193 13674 23321
rect 13741 23121 13771 23321
rect 14427 23191 14457 23319
rect 14511 23191 14541 23319
rect 14699 23241 14729 23325
rect 14784 23241 14814 23325
rect 14879 23241 14909 23325
rect 14982 23241 15012 23325
rect 15114 23175 15144 23325
rect 15209 23241 15239 23325
rect 15293 23241 15323 23325
rect 15407 23241 15437 23325
rect 15618 23125 15648 23325
rect 15702 23125 15732 23325
rect 15890 23197 15920 23325
rect 15987 23125 16017 23325
rect 16709 23191 16739 23319
rect 16793 23191 16823 23319
rect 16981 23241 17011 23325
rect 17066 23241 17096 23325
rect 17161 23241 17191 23325
rect 17264 23241 17294 23325
rect 17396 23175 17426 23325
rect 17491 23241 17521 23325
rect 17575 23241 17605 23325
rect 17689 23241 17719 23325
rect 17900 23125 17930 23325
rect 17984 23125 18014 23325
rect 18172 23197 18202 23325
rect 18269 23125 18299 23325
rect 9556 17297 9586 17497
rect 15693 17149 15723 17349
rect 16471 17187 16501 17387
rect 17345 17189 17375 17389
rect 18113 17179 18143 17379
rect 19235 17181 19265 17381
rect 20109 17183 20139 17383
rect 20877 17173 20907 17373
rect 21491 17171 21521 17371
rect 22365 17173 22395 17373
rect 23133 17163 23163 17363
rect 4555 16339 4585 16539
rect 4639 16339 4669 16539
rect 4723 16339 4753 16539
rect 4807 16339 4837 16539
rect 4995 16339 5025 16539
rect 9421 16343 9451 16543
rect 9505 16343 9535 16543
rect 9589 16343 9619 16543
rect 9673 16343 9703 16543
rect 9861 16343 9891 16543
rect 16456 16447 16486 16647
rect 17224 16437 17254 16637
rect 18098 16439 18128 16639
rect 18712 16437 18742 16637
rect 19480 16427 19510 16627
rect 20354 16429 20384 16629
rect 21476 16431 21506 16631
rect 22244 16421 22274 16621
rect 23118 16423 23148 16623
rect 4681 15669 4711 15753
rect 4765 15669 4795 15753
rect 4873 15595 4903 15795
rect 6687 15601 6717 15685
rect 6787 15601 6817 15685
rect 6891 15601 6921 15685
rect 6977 15601 7007 15685
rect 7143 15485 7173 15685
rect 9547 15673 9577 15757
rect 9631 15673 9661 15757
rect 9739 15599 9769 15799
rect 11553 15605 11583 15689
rect 11653 15605 11683 15689
rect 11757 15605 11787 15689
rect 11843 15605 11873 15689
rect 12009 15489 12039 15689
rect 5865 15059 5895 15143
rect 5949 15059 5979 15143
rect 4565 14775 4595 14975
rect 4649 14775 4679 14975
rect 4733 14775 4763 14975
rect 4817 14775 4847 14975
rect 5005 14775 5035 14975
rect 6057 14985 6087 15185
rect 10731 15063 10761 15147
rect 10815 15063 10845 15147
rect 9431 14779 9461 14979
rect 9515 14779 9545 14979
rect 9599 14779 9629 14979
rect 9683 14779 9713 14979
rect 9871 14779 9901 14979
rect 10923 14989 10953 15189
rect 23563 14701 23593 14785
rect 23647 14701 23677 14785
rect 23835 14651 23865 14735
rect 23919 14651 23949 14735
rect 24107 14701 24137 14785
rect 24293 14651 24323 14735
rect 24377 14651 24407 14735
rect 24472 14701 24502 14785
rect 24556 14701 24586 14785
rect 24744 14701 24774 14785
rect 24932 14701 24962 14785
rect 25029 14654 25059 14738
rect 25307 14585 25337 14785
rect 4691 14105 4721 14189
rect 4775 14105 4805 14189
rect 4883 14031 4913 14231
rect 5903 14135 5933 14219
rect 6003 14135 6033 14219
rect 6107 14135 6137 14219
rect 6193 14135 6223 14219
rect 6359 14019 6389 14219
rect 7801 14003 7831 14087
rect 7897 14003 7927 14087
rect 7969 14003 7999 14087
rect 8065 14003 8095 14087
rect 8163 14003 8193 14203
rect 9557 14109 9587 14193
rect 9641 14109 9671 14193
rect 6914 13645 6944 13729
rect 6986 13645 7016 13729
rect 7083 13645 7113 13845
rect 9749 14035 9779 14235
rect 10769 14139 10799 14223
rect 10869 14139 10899 14223
rect 10973 14139 11003 14223
rect 11059 14139 11089 14223
rect 11225 14023 11255 14223
rect 12667 14007 12697 14091
rect 12763 14007 12793 14091
rect 12835 14007 12865 14091
rect 12931 14007 12961 14091
rect 13029 14007 13059 14207
rect 11780 13649 11810 13733
rect 11852 13649 11882 13733
rect 11949 13649 11979 13849
rect 4557 13107 4587 13307
rect 4641 13107 4671 13307
rect 4725 13107 4755 13307
rect 4809 13107 4839 13307
rect 4997 13107 5027 13307
rect 6027 13180 6057 13264
rect 6111 13180 6141 13264
rect 6204 13180 6234 13264
rect 6299 13177 6329 13377
rect 9423 13111 9453 13311
rect 9507 13111 9537 13311
rect 9591 13111 9621 13311
rect 9675 13111 9705 13311
rect 9863 13111 9893 13311
rect 10893 13184 10923 13268
rect 10977 13184 11007 13268
rect 11070 13184 11100 13268
rect 11165 13181 11195 13381
rect 4683 12437 4713 12521
rect 4767 12437 4797 12521
rect 4875 12363 4905 12563
rect 9549 12441 9579 12525
rect 9633 12441 9663 12525
rect 6059 12231 6089 12315
rect 6143 12231 6173 12315
rect 6251 12157 6281 12357
rect 9741 12367 9771 12567
rect 10925 12235 10955 12319
rect 11009 12235 11039 12319
rect 11117 12161 11147 12361
rect 4567 11543 4597 11743
rect 4651 11543 4681 11743
rect 4735 11543 4765 11743
rect 4819 11543 4849 11743
rect 5007 11543 5037 11743
rect 9433 11547 9463 11747
rect 9517 11547 9547 11747
rect 9601 11547 9631 11747
rect 9685 11547 9715 11747
rect 9873 11547 9903 11747
rect 4693 10873 4723 10957
rect 4777 10873 4807 10957
rect 4885 10799 4915 10999
rect 9559 10877 9589 10961
rect 9643 10877 9673 10961
rect 9751 10803 9781 11003
rect 6238 6103 6268 6303
rect 1950 5051 1980 5251
rect 2049 5051 2079 5135
rect 2145 5051 2175 5135
rect 2217 5051 2247 5135
rect 2313 5051 2343 5135
rect 2402 5051 2432 5135
rect 2486 5051 2516 5135
rect 2570 5051 2600 5135
rect 2758 5051 2788 5135
rect 2842 5051 2872 5135
rect 2926 5051 2956 5135
rect 3010 5051 3040 5135
rect 3100 5051 3130 5135
rect 3199 5051 3229 5251
rect 4084 5043 4114 5243
rect 4183 5043 4213 5127
rect 4279 5043 4309 5127
rect 4351 5043 4381 5127
rect 4447 5043 4477 5127
rect 4536 5043 4566 5127
rect 4620 5043 4650 5127
rect 4704 5043 4734 5127
rect 4892 5043 4922 5127
rect 4976 5043 5006 5127
rect 5060 5043 5090 5127
rect 5144 5043 5174 5127
rect 5234 5043 5264 5127
rect 5333 5043 5363 5243
rect 6036 5043 6066 5243
rect 6135 5043 6165 5127
rect 6231 5043 6261 5127
rect 6303 5043 6333 5127
rect 6399 5043 6429 5127
rect 6488 5043 6518 5127
rect 6572 5043 6602 5127
rect 6656 5043 6686 5127
rect 6844 5043 6874 5127
rect 6928 5043 6958 5127
rect 7012 5043 7042 5127
rect 7096 5043 7126 5127
rect 7186 5043 7216 5127
rect 7285 5043 7315 5243
rect 8038 5049 8068 5249
rect 10132 5471 10162 5671
rect 10231 5471 10261 5555
rect 10327 5471 10357 5555
rect 10399 5471 10429 5555
rect 10495 5471 10525 5555
rect 10584 5471 10614 5555
rect 10668 5471 10698 5555
rect 10752 5471 10782 5555
rect 10940 5471 10970 5555
rect 11024 5471 11054 5555
rect 11108 5471 11138 5555
rect 11192 5471 11222 5555
rect 11282 5471 11312 5555
rect 11381 5471 11411 5671
rect 12194 5459 12224 5659
rect 12293 5459 12323 5543
rect 12389 5459 12419 5543
rect 12461 5459 12491 5543
rect 12557 5459 12587 5543
rect 12646 5459 12676 5543
rect 12730 5459 12760 5543
rect 12814 5459 12844 5543
rect 13002 5459 13032 5543
rect 13086 5459 13116 5543
rect 13170 5459 13200 5543
rect 13254 5459 13284 5543
rect 13344 5459 13374 5543
rect 13443 5459 13473 5659
rect 14152 5467 14182 5667
rect 14251 5467 14281 5551
rect 14347 5467 14377 5551
rect 14419 5467 14449 5551
rect 14515 5467 14545 5551
rect 14604 5467 14634 5551
rect 14688 5467 14718 5551
rect 14772 5467 14802 5551
rect 14960 5467 14990 5551
rect 15044 5467 15074 5551
rect 15128 5467 15158 5551
rect 15212 5467 15242 5551
rect 15302 5467 15332 5551
rect 15401 5467 15431 5667
rect 16146 5473 16176 5673
rect 16245 5473 16275 5557
rect 16341 5473 16371 5557
rect 16413 5473 16443 5557
rect 16509 5473 16539 5557
rect 16598 5473 16628 5557
rect 16682 5473 16712 5557
rect 16766 5473 16796 5557
rect 16954 5473 16984 5557
rect 17038 5473 17068 5557
rect 17122 5473 17152 5557
rect 17206 5473 17236 5557
rect 17296 5473 17326 5557
rect 17395 5473 17425 5673
rect 8137 5049 8167 5133
rect 8233 5049 8263 5133
rect 8305 5049 8335 5133
rect 8401 5049 8431 5133
rect 8490 5049 8520 5133
rect 8574 5049 8604 5133
rect 8658 5049 8688 5133
rect 8846 5049 8876 5133
rect 8930 5049 8960 5133
rect 9014 5049 9044 5133
rect 9098 5049 9128 5133
rect 9188 5049 9218 5133
rect 9287 5049 9317 5249
rect 10160 4597 10190 4797
rect 10259 4597 10289 4681
rect 10355 4597 10385 4681
rect 10427 4597 10457 4681
rect 10523 4597 10553 4681
rect 10612 4597 10642 4681
rect 10696 4597 10726 4681
rect 10780 4597 10810 4681
rect 10968 4597 10998 4681
rect 11052 4597 11082 4681
rect 11136 4597 11166 4681
rect 11220 4597 11250 4681
rect 11310 4597 11340 4681
rect 11409 4597 11439 4797
rect 12430 4553 12460 4753
rect 12529 4553 12559 4637
rect 12625 4553 12655 4637
rect 12697 4553 12727 4637
rect 12793 4553 12823 4637
rect 12882 4553 12912 4637
rect 12966 4553 12996 4637
rect 13050 4553 13080 4637
rect 13238 4553 13268 4637
rect 13322 4553 13352 4637
rect 13406 4553 13436 4637
rect 13490 4553 13520 4637
rect 13580 4553 13610 4637
rect 13679 4553 13709 4753
rect 14432 4547 14462 4747
rect 14531 4547 14561 4631
rect 14627 4547 14657 4631
rect 14699 4547 14729 4631
rect 14795 4547 14825 4631
rect 14884 4547 14914 4631
rect 14968 4547 14998 4631
rect 15052 4547 15082 4631
rect 15240 4547 15270 4631
rect 15324 4547 15354 4631
rect 15408 4547 15438 4631
rect 15492 4547 15522 4631
rect 15582 4547 15612 4631
rect 15681 4547 15711 4747
rect 16454 4529 16484 4729
rect 18427 4938 18457 5022
rect 18523 4938 18553 5022
rect 18595 4938 18625 5022
rect 18809 4938 18839 5022
rect 18912 4938 18942 5022
rect 19021 4899 19051 5099
rect 16553 4529 16583 4613
rect 16649 4529 16679 4613
rect 16721 4529 16751 4613
rect 16817 4529 16847 4613
rect 16906 4529 16936 4613
rect 16990 4529 17020 4613
rect 17074 4529 17104 4613
rect 17262 4529 17292 4613
rect 17346 4529 17376 4613
rect 17430 4529 17460 4613
rect 17514 4529 17544 4613
rect 17604 4529 17634 4613
rect 17703 4529 17733 4729
rect 6208 2843 6238 3043
rect 1920 1791 1950 1991
rect 2019 1791 2049 1875
rect 2115 1791 2145 1875
rect 2187 1791 2217 1875
rect 2283 1791 2313 1875
rect 2372 1791 2402 1875
rect 2456 1791 2486 1875
rect 2540 1791 2570 1875
rect 2728 1791 2758 1875
rect 2812 1791 2842 1875
rect 2896 1791 2926 1875
rect 2980 1791 3010 1875
rect 3070 1791 3100 1875
rect 3169 1791 3199 1991
rect 3990 1787 4020 1987
rect 4089 1787 4119 1871
rect 4185 1787 4215 1871
rect 4257 1787 4287 1871
rect 4353 1787 4383 1871
rect 4442 1787 4472 1871
rect 4526 1787 4556 1871
rect 4610 1787 4640 1871
rect 4798 1787 4828 1871
rect 4882 1787 4912 1871
rect 4966 1787 4996 1871
rect 5050 1787 5080 1871
rect 5140 1787 5170 1871
rect 5239 1787 5269 1987
rect 5942 1787 5972 1987
rect 6041 1787 6071 1871
rect 6137 1787 6167 1871
rect 6209 1787 6239 1871
rect 6305 1787 6335 1871
rect 6394 1787 6424 1871
rect 6478 1787 6508 1871
rect 6562 1787 6592 1871
rect 6750 1787 6780 1871
rect 6834 1787 6864 1871
rect 6918 1787 6948 1871
rect 7002 1787 7032 1871
rect 7092 1787 7122 1871
rect 7191 1787 7221 1987
rect 7944 1793 7974 1993
rect 8043 1793 8073 1877
rect 8139 1793 8169 1877
rect 8211 1793 8241 1877
rect 8307 1793 8337 1877
rect 8396 1793 8426 1877
rect 8480 1793 8510 1877
rect 8564 1793 8594 1877
rect 8752 1793 8782 1877
rect 8836 1793 8866 1877
rect 8920 1793 8950 1877
rect 9004 1793 9034 1877
rect 9094 1793 9124 1877
rect 9193 1793 9223 1993
rect 9896 1793 9926 1993
rect 9995 1793 10025 1877
rect 10091 1793 10121 1877
rect 10163 1793 10193 1877
rect 10259 1793 10289 1877
rect 10348 1793 10378 1877
rect 10432 1793 10462 1877
rect 10516 1793 10546 1877
rect 10704 1793 10734 1877
rect 10788 1793 10818 1877
rect 10872 1793 10902 1877
rect 10956 1793 10986 1877
rect 11046 1793 11076 1877
rect 11145 1793 11175 1993
rect 11888 1793 11918 1993
rect 11987 1793 12017 1877
rect 12083 1793 12113 1877
rect 12155 1793 12185 1877
rect 12251 1793 12281 1877
rect 12340 1793 12370 1877
rect 12424 1793 12454 1877
rect 12508 1793 12538 1877
rect 12696 1793 12726 1877
rect 12780 1793 12810 1877
rect 12864 1793 12894 1877
rect 12948 1793 12978 1877
rect 13038 1793 13068 1877
rect 13137 1793 13167 1993
rect 13840 1793 13870 1993
rect 13939 1793 13969 1877
rect 14035 1793 14065 1877
rect 14107 1793 14137 1877
rect 14203 1793 14233 1877
rect 14292 1793 14322 1877
rect 14376 1793 14406 1877
rect 14460 1793 14490 1877
rect 14648 1793 14678 1877
rect 14732 1793 14762 1877
rect 14816 1793 14846 1877
rect 14900 1793 14930 1877
rect 14990 1793 15020 1877
rect 15089 1793 15119 1993
rect 15904 1793 15934 1993
rect 16003 1793 16033 1877
rect 16099 1793 16129 1877
rect 16171 1793 16201 1877
rect 16267 1793 16297 1877
rect 16356 1793 16386 1877
rect 16440 1793 16470 1877
rect 16524 1793 16554 1877
rect 16712 1793 16742 1877
rect 16796 1793 16826 1877
rect 16880 1793 16910 1877
rect 16964 1793 16994 1877
rect 17054 1793 17084 1877
rect 17153 1793 17183 1993
<< ndiff >>
rect 18963 43374 19093 43382
rect 18963 43340 18979 43374
rect 19013 43340 19047 43374
rect 19081 43340 19093 43374
rect 18963 43330 19093 43340
rect 18963 43290 19093 43300
rect 18963 43256 18979 43290
rect 19013 43256 19047 43290
rect 19081 43256 19093 43290
rect 18963 43246 19093 43256
rect 18963 43206 19093 43216
rect 18963 43172 19047 43206
rect 19081 43172 19093 43206
rect 18963 43162 19093 43172
rect 18963 43122 19093 43132
rect 18963 43088 18979 43122
rect 19013 43088 19047 43122
rect 19081 43088 19093 43122
rect 18963 43078 19093 43088
rect 18963 43038 19093 43048
rect 18963 43004 19047 43038
rect 19081 43004 19093 43038
rect 18963 42994 19093 43004
rect 18963 42954 19093 42964
rect 18963 42920 18979 42954
rect 19013 42920 19047 42954
rect 19081 42920 19093 42954
rect 18963 42910 19093 42920
rect 18963 42870 19093 42880
rect 18963 42836 19047 42870
rect 19081 42836 19093 42870
rect 18963 42826 19093 42836
rect 18963 42786 19093 42796
rect 18963 42752 18979 42786
rect 19013 42752 19047 42786
rect 19081 42752 19093 42786
rect 18963 42742 19093 42752
rect 18963 42702 19093 42712
rect 18963 42668 19047 42702
rect 19081 42668 19093 42702
rect 18963 42658 19093 42668
rect 18963 42618 19093 42628
rect 18963 42584 18979 42618
rect 19013 42584 19047 42618
rect 19081 42584 19093 42618
rect 18963 42574 19093 42584
rect 18963 42534 19093 42544
rect 18963 42500 19047 42534
rect 19081 42500 19093 42534
rect 18963 42490 19093 42500
rect 18963 42450 19093 42460
rect 18963 42416 18979 42450
rect 19013 42416 19047 42450
rect 19081 42416 19093 42450
rect 18963 42406 19093 42416
rect 18963 42366 19093 42376
rect 18963 42332 19047 42366
rect 19081 42332 19093 42366
rect 18963 42322 19093 42332
rect 18963 42282 19093 42292
rect 18963 42248 18979 42282
rect 19013 42248 19047 42282
rect 19081 42248 19093 42282
rect 18963 42238 19093 42248
rect 18963 42198 19093 42208
rect 18963 42164 19047 42198
rect 19081 42164 19093 42198
rect 18963 42154 19093 42164
rect 18963 42114 19093 42124
rect 18963 42080 18979 42114
rect 19013 42080 19047 42114
rect 19081 42080 19093 42114
rect 18963 42070 19093 42080
rect 18963 42030 19093 42040
rect 18963 41996 18979 42030
rect 19013 41996 19047 42030
rect 19081 41996 19093 42030
rect 18963 41988 19093 41996
rect 18947 41397 19077 41405
rect 18947 41363 19031 41397
rect 19065 41363 19077 41397
rect 18947 41302 19077 41363
rect 18947 41262 19077 41272
rect 18947 41228 18963 41262
rect 18997 41228 19031 41262
rect 19065 41228 19077 41262
rect 18947 41218 19077 41228
rect 18947 41178 19077 41188
rect 18947 41144 19031 41178
rect 19065 41144 19077 41178
rect 18947 41134 19077 41144
rect 18947 41094 19077 41104
rect 18947 41060 18963 41094
rect 18997 41060 19031 41094
rect 19065 41060 19077 41094
rect 18947 41050 19077 41060
rect 18947 41010 19077 41020
rect 18947 40976 19031 41010
rect 19065 40976 19077 41010
rect 18947 40966 19077 40976
rect 18947 40926 19077 40936
rect 18947 40892 18963 40926
rect 18997 40892 19031 40926
rect 19065 40892 19077 40926
rect 18947 40882 19077 40892
rect 18947 40842 19077 40852
rect 18947 40808 19031 40842
rect 19065 40808 19077 40842
rect 18947 40798 19077 40808
rect 18947 40758 19077 40768
rect 18947 40724 18963 40758
rect 18997 40724 19031 40758
rect 19065 40724 19077 40758
rect 18947 40714 19077 40724
rect 18947 40674 19077 40684
rect 18947 40640 19031 40674
rect 19065 40640 19077 40674
rect 18947 40630 19077 40640
rect 18947 40590 19077 40600
rect 18947 40556 18963 40590
rect 18997 40556 19031 40590
rect 19065 40556 19077 40590
rect 18947 40546 19077 40556
rect 18947 40506 19077 40516
rect 18947 40472 19031 40506
rect 19065 40472 19077 40506
rect 18947 40462 19077 40472
rect 18947 40422 19077 40432
rect 18947 40388 18963 40422
rect 18997 40388 19031 40422
rect 19065 40388 19077 40422
rect 18947 40378 19077 40388
rect 18947 40338 19077 40348
rect 18947 40304 19031 40338
rect 19065 40304 19077 40338
rect 18947 40296 19077 40304
rect 18955 39582 19085 39590
rect 18955 39548 19039 39582
rect 19073 39548 19085 39582
rect 18955 39538 19085 39548
rect 18955 39498 19085 39508
rect 18955 39464 18971 39498
rect 19005 39464 19039 39498
rect 19073 39464 19085 39498
rect 18955 39454 19085 39464
rect 18955 39414 19085 39424
rect 18955 39380 19039 39414
rect 19073 39380 19085 39414
rect 18955 39370 19085 39380
rect 18955 39330 19085 39340
rect 18955 39296 18971 39330
rect 19005 39296 19039 39330
rect 19073 39296 19085 39330
rect 18955 39286 19085 39296
rect 18955 39246 19085 39256
rect 18955 39212 19039 39246
rect 19073 39212 19085 39246
rect 18955 39202 19085 39212
rect 18955 39162 19085 39172
rect 18955 39128 18971 39162
rect 19005 39128 19039 39162
rect 19073 39128 19085 39162
rect 18955 39118 19085 39128
rect 18955 39078 19085 39088
rect 18955 39044 19039 39078
rect 19073 39044 19085 39078
rect 18955 39034 19085 39044
rect 18955 38994 19085 39004
rect 18955 38960 18971 38994
rect 19005 38960 19039 38994
rect 19073 38960 19085 38994
rect 18955 38950 19085 38960
rect 18955 38910 19085 38920
rect 18955 38876 19039 38910
rect 19073 38876 19085 38910
rect 18955 38868 19085 38876
rect 18969 38337 19099 38347
rect 18969 38303 19052 38337
rect 19086 38303 19099 38337
rect 18969 38293 19099 38303
rect 18969 38253 19099 38263
rect 18969 38219 19045 38253
rect 19079 38219 19099 38253
rect 18969 38209 19099 38219
rect 18969 38169 19099 38179
rect 18969 38135 19053 38169
rect 19087 38135 19099 38169
rect 18969 38125 19099 38135
rect 18969 38085 19099 38095
rect 18969 38051 19045 38085
rect 19079 38051 19099 38085
rect 18969 38041 19099 38051
rect 18969 38001 19099 38011
rect 18969 37967 19053 38001
rect 19087 37967 19099 38001
rect 18969 37957 19099 37967
rect 18969 37917 19099 37927
rect 18969 37883 19045 37917
rect 19079 37883 19099 37917
rect 18969 37873 19099 37883
rect 18969 37809 19099 37843
rect 18969 37775 19053 37809
rect 19087 37775 19099 37809
rect 18969 37767 19099 37775
rect 18981 37179 19111 37187
rect 18981 37145 19064 37179
rect 19098 37145 19111 37179
rect 18981 37135 19111 37145
rect 18981 37095 19111 37105
rect 18981 37061 19057 37095
rect 19091 37061 19111 37095
rect 18981 37051 19111 37061
rect 18981 37011 19111 37021
rect 18981 36977 19065 37011
rect 19099 36977 19111 37011
rect 18981 36967 19111 36977
rect 18981 36927 19111 36937
rect 18981 36893 19057 36927
rect 19091 36893 19111 36927
rect 18981 36883 19111 36893
rect 18981 36843 19111 36853
rect 18981 36809 19065 36843
rect 19099 36809 19111 36843
rect 18981 36801 19111 36809
rect 18989 36299 19119 36307
rect 18989 36265 19001 36299
rect 19035 36265 19073 36299
rect 19107 36265 19119 36299
rect 18989 36255 19119 36265
rect 18989 36215 19119 36225
rect 18989 36181 19001 36215
rect 19035 36181 19073 36215
rect 19107 36181 19119 36215
rect 18989 36171 19119 36181
rect 18989 36131 19119 36141
rect 18989 36097 19001 36131
rect 19035 36097 19073 36131
rect 19107 36097 19119 36131
rect 18989 36089 19119 36097
rect 19013 34913 19143 34921
rect 19013 34879 19059 34913
rect 19093 34879 19143 34913
rect 19013 34869 19143 34879
rect 19013 34829 19143 34839
rect 19013 34795 19097 34829
rect 19131 34795 19143 34829
rect 19013 34789 19143 34795
rect 19059 34774 19143 34789
rect 19059 34734 19143 34744
rect 19059 34700 19071 34734
rect 19105 34700 19143 34734
rect 19059 34692 19143 34700
rect 19013 34630 19143 34638
rect 19013 34596 19026 34630
rect 19060 34596 19094 34630
rect 19128 34596 19143 34630
rect 19013 34586 19143 34596
rect 19013 34546 19143 34556
rect 19013 34512 19067 34546
rect 19101 34512 19143 34546
rect 19013 34502 19143 34512
rect 19013 34462 19143 34472
rect 19013 34428 19028 34462
rect 19062 34428 19096 34462
rect 19130 34428 19143 34462
rect 19013 34420 19143 34428
rect 19059 34356 19143 34364
rect 19059 34322 19083 34356
rect 19117 34322 19143 34356
rect 19059 34312 19143 34322
rect 19059 34232 19143 34282
rect 19071 34217 19143 34232
rect 19071 34158 19143 34187
rect 19071 34124 19083 34158
rect 19117 34124 19143 34158
rect 19071 34111 19143 34124
rect 19071 34060 19143 34081
rect 19015 34055 19143 34060
rect 19015 34021 19083 34055
rect 19117 34021 19143 34055
rect 19015 34010 19143 34021
rect 19015 33936 19143 33980
rect 19015 33930 19089 33936
rect 19059 33902 19089 33930
rect 19123 33902 19143 33936
rect 19059 33891 19143 33902
rect 19059 33811 19143 33861
rect 19071 33792 19143 33811
rect 19071 33737 19143 33762
rect 19071 33703 19083 33737
rect 19117 33703 19143 33737
rect 19071 33693 19143 33703
rect 19071 33631 19143 33663
rect 19059 33626 19143 33631
rect 19059 33592 19083 33626
rect 19117 33592 19143 33626
rect 19059 33581 19143 33592
rect 19059 33541 19143 33551
rect 19059 33507 19097 33541
rect 19131 33507 19143 33541
rect 19059 33499 19143 33507
rect 19059 33437 19143 33445
rect 19059 33403 19071 33437
rect 19105 33403 19143 33437
rect 19059 33393 19143 33403
rect 19059 33353 19143 33363
rect 19059 33319 19097 33353
rect 19131 33319 19143 33353
rect 19059 33309 19143 33319
rect 19059 33269 19143 33279
rect 19059 33235 19071 33269
rect 19105 33235 19143 33269
rect 19059 33227 19143 33235
rect 19013 32631 19143 32639
rect 19013 32597 19059 32631
rect 19093 32597 19143 32631
rect 19013 32587 19143 32597
rect 19013 32547 19143 32557
rect 19013 32513 19097 32547
rect 19131 32513 19143 32547
rect 19013 32507 19143 32513
rect 19059 32492 19143 32507
rect 19059 32452 19143 32462
rect 19059 32418 19071 32452
rect 19105 32418 19143 32452
rect 19059 32410 19143 32418
rect 19013 32348 19143 32356
rect 19013 32314 19026 32348
rect 19060 32314 19094 32348
rect 19128 32314 19143 32348
rect 19013 32304 19143 32314
rect 19013 32264 19143 32274
rect 19013 32230 19067 32264
rect 19101 32230 19143 32264
rect 19013 32220 19143 32230
rect 19013 32180 19143 32190
rect 19013 32146 19028 32180
rect 19062 32146 19096 32180
rect 19130 32146 19143 32180
rect 19013 32138 19143 32146
rect 19059 32074 19143 32082
rect 19059 32040 19083 32074
rect 19117 32040 19143 32074
rect 19059 32030 19143 32040
rect 19059 31950 19143 32000
rect 19071 31935 19143 31950
rect 19071 31876 19143 31905
rect 19071 31842 19083 31876
rect 19117 31842 19143 31876
rect 19071 31829 19143 31842
rect 19071 31778 19143 31799
rect 19015 31773 19143 31778
rect 19015 31739 19083 31773
rect 19117 31739 19143 31773
rect 19015 31728 19143 31739
rect 19015 31654 19143 31698
rect 19015 31648 19089 31654
rect 19059 31620 19089 31648
rect 19123 31620 19143 31654
rect 19059 31609 19143 31620
rect 19059 31529 19143 31579
rect 19071 31510 19143 31529
rect 19071 31455 19143 31480
rect 19071 31421 19083 31455
rect 19117 31421 19143 31455
rect 19071 31411 19143 31421
rect 19071 31349 19143 31381
rect 19059 31344 19143 31349
rect 19059 31310 19083 31344
rect 19117 31310 19143 31344
rect 19059 31299 19143 31310
rect 19059 31259 19143 31269
rect 19059 31225 19097 31259
rect 19131 31225 19143 31259
rect 19059 31217 19143 31225
rect 19059 31155 19143 31163
rect 19059 31121 19071 31155
rect 19105 31121 19143 31155
rect 19059 31111 19143 31121
rect 19059 31071 19143 31081
rect 19059 31037 19097 31071
rect 19131 31037 19143 31071
rect 19059 31027 19143 31037
rect 19059 30987 19143 30997
rect 19059 30953 19071 30987
rect 19105 30953 19143 30987
rect 19059 30945 19143 30953
rect 19017 30385 19147 30393
rect 19017 30351 19063 30385
rect 19097 30351 19147 30385
rect 19017 30341 19147 30351
rect 19017 30301 19147 30311
rect 19017 30267 19101 30301
rect 19135 30267 19147 30301
rect 19017 30261 19147 30267
rect 19063 30246 19147 30261
rect 19063 30206 19147 30216
rect 19063 30172 19075 30206
rect 19109 30172 19147 30206
rect 19063 30164 19147 30172
rect 19017 30102 19147 30110
rect 19017 30068 19030 30102
rect 19064 30068 19098 30102
rect 19132 30068 19147 30102
rect 19017 30058 19147 30068
rect 19017 30018 19147 30028
rect 19017 29984 19071 30018
rect 19105 29984 19147 30018
rect 19017 29974 19147 29984
rect 19017 29934 19147 29944
rect 19017 29900 19032 29934
rect 19066 29900 19100 29934
rect 19134 29900 19147 29934
rect 19017 29892 19147 29900
rect 19063 29828 19147 29836
rect 19063 29794 19087 29828
rect 19121 29794 19147 29828
rect 19063 29784 19147 29794
rect 19063 29704 19147 29754
rect 19075 29689 19147 29704
rect 19075 29630 19147 29659
rect 19075 29596 19087 29630
rect 19121 29596 19147 29630
rect 19075 29583 19147 29596
rect 19075 29532 19147 29553
rect 19019 29527 19147 29532
rect 19019 29493 19087 29527
rect 19121 29493 19147 29527
rect 19019 29482 19147 29493
rect 19019 29408 19147 29452
rect 19019 29402 19093 29408
rect 19063 29374 19093 29402
rect 19127 29374 19147 29408
rect 19063 29363 19147 29374
rect 19063 29283 19147 29333
rect 19075 29264 19147 29283
rect 19075 29209 19147 29234
rect 19075 29175 19087 29209
rect 19121 29175 19147 29209
rect 19075 29165 19147 29175
rect 19075 29103 19147 29135
rect 19063 29098 19147 29103
rect 19063 29064 19087 29098
rect 19121 29064 19147 29098
rect 19063 29053 19147 29064
rect 19063 29013 19147 29023
rect 19063 28979 19101 29013
rect 19135 28979 19147 29013
rect 19063 28971 19147 28979
rect 19063 28909 19147 28917
rect 19063 28875 19075 28909
rect 19109 28875 19147 28909
rect 19063 28865 19147 28875
rect 19063 28825 19147 28835
rect 19063 28791 19101 28825
rect 19135 28791 19147 28825
rect 19063 28781 19147 28791
rect 19063 28741 19147 28751
rect 19063 28707 19075 28741
rect 19109 28707 19147 28741
rect 19063 28699 19147 28707
rect 19009 28199 19139 28207
rect 19009 28165 19055 28199
rect 19089 28165 19139 28199
rect 19009 28155 19139 28165
rect 19009 28115 19139 28125
rect 19009 28081 19093 28115
rect 19127 28081 19139 28115
rect 19009 28075 19139 28081
rect 19055 28060 19139 28075
rect 19055 28020 19139 28030
rect 19055 27986 19067 28020
rect 19101 27986 19139 28020
rect 19055 27978 19139 27986
rect 19009 27916 19139 27924
rect 19009 27882 19022 27916
rect 19056 27882 19090 27916
rect 19124 27882 19139 27916
rect 19009 27872 19139 27882
rect 19009 27832 19139 27842
rect 19009 27798 19063 27832
rect 19097 27798 19139 27832
rect 19009 27788 19139 27798
rect 19009 27748 19139 27758
rect 19009 27714 19024 27748
rect 19058 27714 19092 27748
rect 19126 27714 19139 27748
rect 19009 27706 19139 27714
rect 19055 27642 19139 27650
rect 19055 27608 19079 27642
rect 19113 27608 19139 27642
rect 19055 27598 19139 27608
rect 19055 27518 19139 27568
rect 19067 27503 19139 27518
rect 19067 27444 19139 27473
rect 19067 27410 19079 27444
rect 19113 27410 19139 27444
rect 19067 27397 19139 27410
rect 19067 27346 19139 27367
rect 19011 27341 19139 27346
rect 19011 27307 19079 27341
rect 19113 27307 19139 27341
rect 19011 27296 19139 27307
rect 19011 27222 19139 27266
rect 19011 27216 19085 27222
rect 19055 27188 19085 27216
rect 19119 27188 19139 27222
rect 19055 27177 19139 27188
rect 19055 27097 19139 27147
rect 19067 27078 19139 27097
rect 19067 27023 19139 27048
rect 19067 26989 19079 27023
rect 19113 26989 19139 27023
rect 19067 26979 19139 26989
rect 19067 26917 19139 26949
rect 19055 26912 19139 26917
rect 19055 26878 19079 26912
rect 19113 26878 19139 26912
rect 19055 26867 19139 26878
rect 19055 26827 19139 26837
rect 19055 26793 19093 26827
rect 19127 26793 19139 26827
rect 19055 26785 19139 26793
rect 19055 26723 19139 26731
rect 19055 26689 19067 26723
rect 19101 26689 19139 26723
rect 19055 26679 19139 26689
rect 19055 26639 19139 26649
rect 19055 26605 19093 26639
rect 19127 26605 19139 26639
rect 19055 26595 19139 26605
rect 19055 26555 19139 26565
rect 19055 26521 19067 26555
rect 19101 26521 19139 26555
rect 19055 26513 19139 26521
rect 19013 25953 19143 25961
rect 19013 25919 19059 25953
rect 19093 25919 19143 25953
rect 19013 25909 19143 25919
rect 19013 25869 19143 25879
rect 19013 25835 19097 25869
rect 19131 25835 19143 25869
rect 19013 25829 19143 25835
rect 19059 25814 19143 25829
rect 19059 25774 19143 25784
rect 19059 25740 19071 25774
rect 19105 25740 19143 25774
rect 19059 25732 19143 25740
rect 19013 25670 19143 25678
rect 19013 25636 19026 25670
rect 19060 25636 19094 25670
rect 19128 25636 19143 25670
rect 19013 25626 19143 25636
rect 19013 25586 19143 25596
rect 19013 25552 19067 25586
rect 19101 25552 19143 25586
rect 19013 25542 19143 25552
rect 19013 25502 19143 25512
rect 19013 25468 19028 25502
rect 19062 25468 19096 25502
rect 19130 25468 19143 25502
rect 19013 25460 19143 25468
rect 19059 25396 19143 25404
rect 19059 25362 19083 25396
rect 19117 25362 19143 25396
rect 19059 25352 19143 25362
rect 19059 25272 19143 25322
rect 19071 25257 19143 25272
rect 19071 25198 19143 25227
rect 19071 25164 19083 25198
rect 19117 25164 19143 25198
rect 19071 25151 19143 25164
rect 19071 25100 19143 25121
rect 19015 25095 19143 25100
rect 19015 25061 19083 25095
rect 19117 25061 19143 25095
rect 19015 25050 19143 25061
rect 19015 24976 19143 25020
rect 19015 24970 19089 24976
rect 19059 24942 19089 24970
rect 19123 24942 19143 24976
rect 19059 24931 19143 24942
rect 19059 24851 19143 24901
rect 19071 24832 19143 24851
rect 19071 24777 19143 24802
rect 19071 24743 19083 24777
rect 19117 24743 19143 24777
rect 19071 24733 19143 24743
rect 19071 24671 19143 24703
rect 19059 24666 19143 24671
rect 19059 24632 19083 24666
rect 19117 24632 19143 24666
rect 19059 24621 19143 24632
rect 19059 24581 19143 24591
rect 19059 24547 19097 24581
rect 19131 24547 19143 24581
rect 19059 24539 19143 24547
rect 19059 24477 19143 24485
rect 19059 24443 19071 24477
rect 19105 24443 19143 24477
rect 19059 24433 19143 24443
rect 19059 24393 19143 24403
rect 19059 24359 19097 24393
rect 19131 24359 19143 24393
rect 19059 24349 19143 24359
rect 19059 24309 19143 24319
rect 19059 24275 19071 24309
rect 19105 24275 19143 24309
rect 19059 24267 19143 24275
rect 7697 22947 7749 22959
rect 7697 22913 7705 22947
rect 7739 22913 7749 22947
rect 7697 22875 7749 22913
rect 7779 22921 7833 22959
rect 7779 22887 7789 22921
rect 7823 22887 7833 22921
rect 7779 22875 7833 22887
rect 7863 22947 7915 22959
rect 7863 22913 7873 22947
rect 7907 22913 7915 22947
rect 7863 22875 7915 22913
rect 7969 22921 8021 22959
rect 7969 22887 7977 22921
rect 8011 22887 8021 22921
rect 7969 22875 8021 22887
rect 8051 22947 8101 22959
rect 8400 22959 8450 23003
rect 8281 22947 8331 22959
rect 8051 22935 8133 22947
rect 8051 22901 8062 22935
rect 8096 22901 8133 22935
rect 8051 22875 8133 22901
rect 8163 22935 8232 22947
rect 8163 22901 8173 22935
rect 8207 22901 8232 22935
rect 8163 22875 8232 22901
rect 8262 22875 8331 22947
rect 8361 22929 8450 22959
rect 8361 22895 8372 22929
rect 8406 22895 8450 22929
rect 8361 22875 8450 22895
rect 8480 22947 8530 23003
rect 8890 22990 8942 23005
rect 8702 22947 8752 22959
rect 8480 22935 8551 22947
rect 8480 22901 8491 22935
rect 8525 22901 8551 22935
rect 8480 22875 8551 22901
rect 8581 22935 8657 22947
rect 8581 22901 8594 22935
rect 8628 22901 8657 22935
rect 8581 22875 8657 22901
rect 8687 22875 8752 22947
rect 8782 22935 8834 22959
rect 8782 22901 8792 22935
rect 8826 22901 8834 22935
rect 8782 22875 8834 22901
rect 8890 22956 8898 22990
rect 8932 22956 8942 22990
rect 8890 22922 8942 22956
rect 8890 22888 8898 22922
rect 8932 22888 8942 22922
rect 8890 22875 8942 22888
rect 8972 22951 9026 23005
rect 8972 22917 8982 22951
rect 9016 22917 9026 22951
rect 8972 22875 9026 22917
rect 9056 22992 9108 23005
rect 9056 22958 9066 22992
rect 9100 22958 9108 22992
rect 9259 22959 9309 23005
rect 9056 22924 9108 22958
rect 9056 22890 9066 22924
rect 9100 22890 9108 22924
rect 9056 22875 9108 22890
rect 9162 22947 9214 22959
rect 9162 22913 9170 22947
rect 9204 22913 9214 22947
rect 9162 22875 9214 22913
rect 9244 22921 9309 22959
rect 9244 22887 9265 22921
rect 9299 22887 9309 22921
rect 9244 22875 9309 22887
rect 9339 22959 9391 23005
rect 9339 22925 9349 22959
rect 9383 22925 9391 22959
rect 9339 22875 9391 22925
rect 9943 22951 9995 22963
rect 9943 22917 9951 22951
rect 9985 22917 9995 22951
rect 9943 22879 9995 22917
rect 10025 22925 10079 22963
rect 10025 22891 10035 22925
rect 10069 22891 10079 22925
rect 10025 22879 10079 22891
rect 10109 22951 10161 22963
rect 10109 22917 10119 22951
rect 10153 22917 10161 22951
rect 10109 22879 10161 22917
rect 10215 22925 10267 22963
rect 10215 22891 10223 22925
rect 10257 22891 10267 22925
rect 10215 22879 10267 22891
rect 10297 22951 10347 22963
rect 10646 22963 10696 23007
rect 10527 22951 10577 22963
rect 10297 22939 10379 22951
rect 10297 22905 10308 22939
rect 10342 22905 10379 22939
rect 10297 22879 10379 22905
rect 10409 22939 10478 22951
rect 10409 22905 10419 22939
rect 10453 22905 10478 22939
rect 10409 22879 10478 22905
rect 10508 22879 10577 22951
rect 10607 22933 10696 22963
rect 10607 22899 10618 22933
rect 10652 22899 10696 22933
rect 10607 22879 10696 22899
rect 10726 22951 10776 23007
rect 11136 22994 11188 23009
rect 10948 22951 10998 22963
rect 10726 22939 10797 22951
rect 10726 22905 10737 22939
rect 10771 22905 10797 22939
rect 10726 22879 10797 22905
rect 10827 22939 10903 22951
rect 10827 22905 10840 22939
rect 10874 22905 10903 22939
rect 10827 22879 10903 22905
rect 10933 22879 10998 22951
rect 11028 22939 11080 22963
rect 11028 22905 11038 22939
rect 11072 22905 11080 22939
rect 11028 22879 11080 22905
rect 11136 22960 11144 22994
rect 11178 22960 11188 22994
rect 11136 22926 11188 22960
rect 11136 22892 11144 22926
rect 11178 22892 11188 22926
rect 11136 22879 11188 22892
rect 11218 22955 11272 23009
rect 11218 22921 11228 22955
rect 11262 22921 11272 22955
rect 11218 22879 11272 22921
rect 11302 22996 11354 23009
rect 11302 22962 11312 22996
rect 11346 22962 11354 22996
rect 11505 22963 11555 23009
rect 11302 22928 11354 22962
rect 11302 22894 11312 22928
rect 11346 22894 11354 22928
rect 11302 22879 11354 22894
rect 11408 22951 11460 22963
rect 11408 22917 11416 22951
rect 11450 22917 11460 22951
rect 11408 22879 11460 22917
rect 11490 22925 11555 22963
rect 11490 22891 11511 22925
rect 11545 22891 11555 22925
rect 11490 22879 11555 22891
rect 11585 22963 11637 23009
rect 11585 22929 11595 22963
rect 11629 22929 11637 22963
rect 11585 22879 11637 22929
rect 12129 22943 12181 22955
rect 12129 22909 12137 22943
rect 12171 22909 12181 22943
rect 12129 22871 12181 22909
rect 12211 22917 12265 22955
rect 12211 22883 12221 22917
rect 12255 22883 12265 22917
rect 12211 22871 12265 22883
rect 12295 22943 12347 22955
rect 12295 22909 12305 22943
rect 12339 22909 12347 22943
rect 12295 22871 12347 22909
rect 12401 22917 12453 22955
rect 12401 22883 12409 22917
rect 12443 22883 12453 22917
rect 12401 22871 12453 22883
rect 12483 22943 12533 22955
rect 12832 22955 12882 22999
rect 12713 22943 12763 22955
rect 12483 22931 12565 22943
rect 12483 22897 12494 22931
rect 12528 22897 12565 22931
rect 12483 22871 12565 22897
rect 12595 22931 12664 22943
rect 12595 22897 12605 22931
rect 12639 22897 12664 22931
rect 12595 22871 12664 22897
rect 12694 22871 12763 22943
rect 12793 22925 12882 22955
rect 12793 22891 12804 22925
rect 12838 22891 12882 22925
rect 12793 22871 12882 22891
rect 12912 22943 12962 22999
rect 13322 22986 13374 23001
rect 13134 22943 13184 22955
rect 12912 22931 12983 22943
rect 12912 22897 12923 22931
rect 12957 22897 12983 22931
rect 12912 22871 12983 22897
rect 13013 22931 13089 22943
rect 13013 22897 13026 22931
rect 13060 22897 13089 22931
rect 13013 22871 13089 22897
rect 13119 22871 13184 22943
rect 13214 22931 13266 22955
rect 13214 22897 13224 22931
rect 13258 22897 13266 22931
rect 13214 22871 13266 22897
rect 13322 22952 13330 22986
rect 13364 22952 13374 22986
rect 13322 22918 13374 22952
rect 13322 22884 13330 22918
rect 13364 22884 13374 22918
rect 13322 22871 13374 22884
rect 13404 22947 13458 23001
rect 13404 22913 13414 22947
rect 13448 22913 13458 22947
rect 13404 22871 13458 22913
rect 13488 22988 13540 23001
rect 13488 22954 13498 22988
rect 13532 22954 13540 22988
rect 13691 22955 13741 23001
rect 13488 22920 13540 22954
rect 13488 22886 13498 22920
rect 13532 22886 13540 22920
rect 13488 22871 13540 22886
rect 13594 22943 13646 22955
rect 13594 22909 13602 22943
rect 13636 22909 13646 22943
rect 13594 22871 13646 22909
rect 13676 22917 13741 22955
rect 13676 22883 13697 22917
rect 13731 22883 13741 22917
rect 13676 22871 13741 22883
rect 13771 22955 13823 23001
rect 13771 22921 13781 22955
rect 13815 22921 13823 22955
rect 13771 22871 13823 22921
rect 14375 22947 14427 22959
rect 14375 22913 14383 22947
rect 14417 22913 14427 22947
rect 14375 22875 14427 22913
rect 14457 22921 14511 22959
rect 14457 22887 14467 22921
rect 14501 22887 14511 22921
rect 14457 22875 14511 22887
rect 14541 22947 14593 22959
rect 14541 22913 14551 22947
rect 14585 22913 14593 22947
rect 14541 22875 14593 22913
rect 14647 22921 14699 22959
rect 14647 22887 14655 22921
rect 14689 22887 14699 22921
rect 14647 22875 14699 22887
rect 14729 22947 14779 22959
rect 15078 22959 15128 23003
rect 14959 22947 15009 22959
rect 14729 22935 14811 22947
rect 14729 22901 14740 22935
rect 14774 22901 14811 22935
rect 14729 22875 14811 22901
rect 14841 22935 14910 22947
rect 14841 22901 14851 22935
rect 14885 22901 14910 22935
rect 14841 22875 14910 22901
rect 14940 22875 15009 22947
rect 15039 22929 15128 22959
rect 15039 22895 15050 22929
rect 15084 22895 15128 22929
rect 15039 22875 15128 22895
rect 15158 22947 15208 23003
rect 15568 22990 15620 23005
rect 15380 22947 15430 22959
rect 15158 22935 15229 22947
rect 15158 22901 15169 22935
rect 15203 22901 15229 22935
rect 15158 22875 15229 22901
rect 15259 22935 15335 22947
rect 15259 22901 15272 22935
rect 15306 22901 15335 22935
rect 15259 22875 15335 22901
rect 15365 22875 15430 22947
rect 15460 22935 15512 22959
rect 15460 22901 15470 22935
rect 15504 22901 15512 22935
rect 15460 22875 15512 22901
rect 15568 22956 15576 22990
rect 15610 22956 15620 22990
rect 15568 22922 15620 22956
rect 15568 22888 15576 22922
rect 15610 22888 15620 22922
rect 15568 22875 15620 22888
rect 15650 22951 15704 23005
rect 15650 22917 15660 22951
rect 15694 22917 15704 22951
rect 15650 22875 15704 22917
rect 15734 22992 15786 23005
rect 15734 22958 15744 22992
rect 15778 22958 15786 22992
rect 15937 22959 15987 23005
rect 15734 22924 15786 22958
rect 15734 22890 15744 22924
rect 15778 22890 15786 22924
rect 15734 22875 15786 22890
rect 15840 22947 15892 22959
rect 15840 22913 15848 22947
rect 15882 22913 15892 22947
rect 15840 22875 15892 22913
rect 15922 22921 15987 22959
rect 15922 22887 15943 22921
rect 15977 22887 15987 22921
rect 15922 22875 15987 22887
rect 16017 22959 16069 23005
rect 16017 22925 16027 22959
rect 16061 22925 16069 22959
rect 16017 22875 16069 22925
rect 16657 22947 16709 22959
rect 16657 22913 16665 22947
rect 16699 22913 16709 22947
rect 16657 22875 16709 22913
rect 16739 22921 16793 22959
rect 16739 22887 16749 22921
rect 16783 22887 16793 22921
rect 16739 22875 16793 22887
rect 16823 22947 16875 22959
rect 16823 22913 16833 22947
rect 16867 22913 16875 22947
rect 16823 22875 16875 22913
rect 16929 22921 16981 22959
rect 16929 22887 16937 22921
rect 16971 22887 16981 22921
rect 16929 22875 16981 22887
rect 17011 22947 17061 22959
rect 17360 22959 17410 23003
rect 17241 22947 17291 22959
rect 17011 22935 17093 22947
rect 17011 22901 17022 22935
rect 17056 22901 17093 22935
rect 17011 22875 17093 22901
rect 17123 22935 17192 22947
rect 17123 22901 17133 22935
rect 17167 22901 17192 22935
rect 17123 22875 17192 22901
rect 17222 22875 17291 22947
rect 17321 22929 17410 22959
rect 17321 22895 17332 22929
rect 17366 22895 17410 22929
rect 17321 22875 17410 22895
rect 17440 22947 17490 23003
rect 17850 22990 17902 23005
rect 17662 22947 17712 22959
rect 17440 22935 17511 22947
rect 17440 22901 17451 22935
rect 17485 22901 17511 22935
rect 17440 22875 17511 22901
rect 17541 22935 17617 22947
rect 17541 22901 17554 22935
rect 17588 22901 17617 22935
rect 17541 22875 17617 22901
rect 17647 22875 17712 22947
rect 17742 22935 17794 22959
rect 17742 22901 17752 22935
rect 17786 22901 17794 22935
rect 17742 22875 17794 22901
rect 17850 22956 17858 22990
rect 17892 22956 17902 22990
rect 17850 22922 17902 22956
rect 17850 22888 17858 22922
rect 17892 22888 17902 22922
rect 17850 22875 17902 22888
rect 17932 22951 17986 23005
rect 17932 22917 17942 22951
rect 17976 22917 17986 22951
rect 17932 22875 17986 22917
rect 18016 22992 18068 23005
rect 18016 22958 18026 22992
rect 18060 22958 18068 22992
rect 18219 22959 18269 23005
rect 18016 22924 18068 22958
rect 18016 22890 18026 22924
rect 18060 22890 18068 22924
rect 18016 22875 18068 22890
rect 18122 22947 18174 22959
rect 18122 22913 18130 22947
rect 18164 22913 18174 22947
rect 18122 22875 18174 22913
rect 18204 22921 18269 22959
rect 18204 22887 18225 22921
rect 18259 22887 18269 22921
rect 18204 22875 18269 22887
rect 18299 22959 18351 23005
rect 18299 22925 18309 22959
rect 18343 22925 18351 22959
rect 18299 22875 18351 22925
rect 9504 17731 9556 17747
rect 9504 17697 9512 17731
rect 9546 17697 9556 17731
rect 9504 17663 9556 17697
rect 9504 17629 9512 17663
rect 9546 17629 9556 17663
rect 9504 17617 9556 17629
rect 9586 17731 9638 17747
rect 9586 17697 9596 17731
rect 9630 17697 9638 17731
rect 9586 17663 9638 17697
rect 9586 17629 9596 17663
rect 9630 17629 9638 17663
rect 9586 17617 9638 17629
rect 16419 17621 16471 17637
rect 15641 17583 15693 17599
rect 15641 17549 15649 17583
rect 15683 17549 15693 17583
rect 15641 17515 15693 17549
rect 15641 17481 15649 17515
rect 15683 17481 15693 17515
rect 15641 17469 15693 17481
rect 15723 17583 15775 17599
rect 15723 17549 15733 17583
rect 15767 17549 15775 17583
rect 15723 17515 15775 17549
rect 16419 17587 16427 17621
rect 16461 17587 16471 17621
rect 16419 17553 16471 17587
rect 16419 17519 16427 17553
rect 16461 17519 16471 17553
rect 15723 17481 15733 17515
rect 15767 17481 15775 17515
rect 16419 17507 16471 17519
rect 16501 17621 16553 17637
rect 17293 17623 17345 17639
rect 16501 17587 16511 17621
rect 16545 17587 16553 17621
rect 16501 17553 16553 17587
rect 16501 17519 16511 17553
rect 16545 17519 16553 17553
rect 16501 17507 16553 17519
rect 17293 17589 17301 17623
rect 17335 17589 17345 17623
rect 17293 17555 17345 17589
rect 17293 17521 17301 17555
rect 17335 17521 17345 17555
rect 17293 17509 17345 17521
rect 17375 17623 17427 17639
rect 17375 17589 17385 17623
rect 17419 17589 17427 17623
rect 18061 17613 18113 17629
rect 17375 17555 17427 17589
rect 17375 17521 17385 17555
rect 17419 17521 17427 17555
rect 17375 17509 17427 17521
rect 15723 17469 15775 17481
rect 18061 17579 18069 17613
rect 18103 17579 18113 17613
rect 18061 17545 18113 17579
rect 18061 17511 18069 17545
rect 18103 17511 18113 17545
rect 18061 17499 18113 17511
rect 18143 17613 18195 17629
rect 19183 17615 19235 17631
rect 18143 17579 18153 17613
rect 18187 17579 18195 17613
rect 18143 17545 18195 17579
rect 18143 17511 18153 17545
rect 18187 17511 18195 17545
rect 18143 17499 18195 17511
rect 19183 17581 19191 17615
rect 19225 17581 19235 17615
rect 19183 17547 19235 17581
rect 19183 17513 19191 17547
rect 19225 17513 19235 17547
rect 19183 17501 19235 17513
rect 19265 17615 19317 17631
rect 20057 17617 20109 17633
rect 19265 17581 19275 17615
rect 19309 17581 19317 17615
rect 19265 17547 19317 17581
rect 19265 17513 19275 17547
rect 19309 17513 19317 17547
rect 19265 17501 19317 17513
rect 20057 17583 20065 17617
rect 20099 17583 20109 17617
rect 20057 17549 20109 17583
rect 20057 17515 20065 17549
rect 20099 17515 20109 17549
rect 20057 17503 20109 17515
rect 20139 17617 20191 17633
rect 20139 17583 20149 17617
rect 20183 17583 20191 17617
rect 20825 17607 20877 17623
rect 20139 17549 20191 17583
rect 20139 17515 20149 17549
rect 20183 17515 20191 17549
rect 20139 17503 20191 17515
rect 20825 17573 20833 17607
rect 20867 17573 20877 17607
rect 20825 17539 20877 17573
rect 20825 17505 20833 17539
rect 20867 17505 20877 17539
rect 20825 17493 20877 17505
rect 20907 17607 20959 17623
rect 20907 17573 20917 17607
rect 20951 17573 20959 17607
rect 20907 17539 20959 17573
rect 20907 17505 20917 17539
rect 20951 17505 20959 17539
rect 20907 17493 20959 17505
rect 21439 17605 21491 17621
rect 21439 17571 21447 17605
rect 21481 17571 21491 17605
rect 21439 17537 21491 17571
rect 21439 17503 21447 17537
rect 21481 17503 21491 17537
rect 21439 17491 21491 17503
rect 21521 17605 21573 17621
rect 22313 17607 22365 17623
rect 21521 17571 21531 17605
rect 21565 17571 21573 17605
rect 21521 17537 21573 17571
rect 21521 17503 21531 17537
rect 21565 17503 21573 17537
rect 21521 17491 21573 17503
rect 22313 17573 22321 17607
rect 22355 17573 22365 17607
rect 22313 17539 22365 17573
rect 22313 17505 22321 17539
rect 22355 17505 22365 17539
rect 22313 17493 22365 17505
rect 22395 17607 22447 17623
rect 22395 17573 22405 17607
rect 22439 17573 22447 17607
rect 22395 17539 22447 17573
rect 22395 17505 22405 17539
rect 22439 17505 22447 17539
rect 22395 17493 22447 17505
rect 23081 17597 23133 17613
rect 23081 17563 23089 17597
rect 23123 17563 23133 17597
rect 23081 17529 23133 17563
rect 23081 17495 23089 17529
rect 23123 17495 23133 17529
rect 23081 17483 23133 17495
rect 23163 17597 23215 17613
rect 23163 17563 23173 17597
rect 23207 17563 23215 17597
rect 23163 17529 23215 17563
rect 23163 17495 23173 17529
rect 23207 17495 23215 17529
rect 23163 17483 23215 17495
rect 4503 16137 4555 16219
rect 4503 16103 4511 16137
rect 4545 16103 4555 16137
rect 4503 16089 4555 16103
rect 4585 16159 4639 16219
rect 4585 16125 4595 16159
rect 4629 16125 4639 16159
rect 4585 16089 4639 16125
rect 4669 16137 4723 16219
rect 4669 16103 4679 16137
rect 4713 16103 4723 16137
rect 4669 16089 4723 16103
rect 4753 16089 4807 16219
rect 4837 16139 4991 16219
rect 4837 16105 4847 16139
rect 4881 16105 4947 16139
rect 4981 16105 4991 16139
rect 4837 16089 4991 16105
rect 5021 16210 5085 16219
rect 5021 16176 5037 16210
rect 5071 16176 5085 16210
rect 5021 16142 5085 16176
rect 5021 16108 5037 16142
rect 5071 16108 5085 16142
rect 9369 16141 9421 16223
rect 5021 16089 5085 16108
rect 9369 16107 9377 16141
rect 9411 16107 9421 16141
rect 9369 16093 9421 16107
rect 9451 16163 9505 16223
rect 9451 16129 9461 16163
rect 9495 16129 9505 16163
rect 9451 16093 9505 16129
rect 9535 16141 9589 16223
rect 9535 16107 9545 16141
rect 9579 16107 9589 16141
rect 9535 16093 9589 16107
rect 9619 16093 9673 16223
rect 9703 16143 9857 16223
rect 9703 16109 9713 16143
rect 9747 16109 9813 16143
rect 9847 16109 9857 16143
rect 9703 16093 9857 16109
rect 9887 16214 9951 16223
rect 16404 16315 16456 16327
rect 16404 16281 16412 16315
rect 16446 16281 16456 16315
rect 16404 16247 16456 16281
rect 9887 16180 9903 16214
rect 9937 16180 9951 16214
rect 16404 16213 16412 16247
rect 16446 16213 16456 16247
rect 16404 16197 16456 16213
rect 16486 16315 16538 16327
rect 16486 16281 16496 16315
rect 16530 16281 16538 16315
rect 16486 16247 16538 16281
rect 16486 16213 16496 16247
rect 16530 16213 16538 16247
rect 16486 16197 16538 16213
rect 17172 16305 17224 16317
rect 17172 16271 17180 16305
rect 17214 16271 17224 16305
rect 17172 16237 17224 16271
rect 17172 16203 17180 16237
rect 17214 16203 17224 16237
rect 9887 16146 9951 16180
rect 17172 16187 17224 16203
rect 17254 16305 17306 16317
rect 17254 16271 17264 16305
rect 17298 16271 17306 16305
rect 17254 16237 17306 16271
rect 17254 16203 17264 16237
rect 17298 16203 17306 16237
rect 18046 16307 18098 16319
rect 18046 16273 18054 16307
rect 18088 16273 18098 16307
rect 18046 16239 18098 16273
rect 18046 16205 18054 16239
rect 18088 16205 18098 16239
rect 17254 16187 17306 16203
rect 18046 16189 18098 16205
rect 18128 16307 18180 16319
rect 18128 16273 18138 16307
rect 18172 16273 18180 16307
rect 18128 16239 18180 16273
rect 18128 16205 18138 16239
rect 18172 16205 18180 16239
rect 18128 16189 18180 16205
rect 18660 16305 18712 16317
rect 18660 16271 18668 16305
rect 18702 16271 18712 16305
rect 18660 16237 18712 16271
rect 18660 16203 18668 16237
rect 18702 16203 18712 16237
rect 18660 16187 18712 16203
rect 18742 16305 18794 16317
rect 18742 16271 18752 16305
rect 18786 16271 18794 16305
rect 18742 16237 18794 16271
rect 18742 16203 18752 16237
rect 18786 16203 18794 16237
rect 19428 16295 19480 16307
rect 19428 16261 19436 16295
rect 19470 16261 19480 16295
rect 19428 16227 19480 16261
rect 18742 16187 18794 16203
rect 19428 16193 19436 16227
rect 19470 16193 19480 16227
rect 19428 16177 19480 16193
rect 19510 16295 19562 16307
rect 19510 16261 19520 16295
rect 19554 16261 19562 16295
rect 19510 16227 19562 16261
rect 19510 16193 19520 16227
rect 19554 16193 19562 16227
rect 20302 16297 20354 16309
rect 20302 16263 20310 16297
rect 20344 16263 20354 16297
rect 20302 16229 20354 16263
rect 20302 16195 20310 16229
rect 20344 16195 20354 16229
rect 19510 16177 19562 16193
rect 20302 16179 20354 16195
rect 20384 16297 20436 16309
rect 20384 16263 20394 16297
rect 20428 16263 20436 16297
rect 20384 16229 20436 16263
rect 20384 16195 20394 16229
rect 20428 16195 20436 16229
rect 21424 16299 21476 16311
rect 21424 16265 21432 16299
rect 21466 16265 21476 16299
rect 21424 16231 21476 16265
rect 21424 16197 21432 16231
rect 21466 16197 21476 16231
rect 20384 16179 20436 16195
rect 21424 16181 21476 16197
rect 21506 16299 21558 16311
rect 21506 16265 21516 16299
rect 21550 16265 21558 16299
rect 21506 16231 21558 16265
rect 21506 16197 21516 16231
rect 21550 16197 21558 16231
rect 22192 16289 22244 16301
rect 22192 16255 22200 16289
rect 22234 16255 22244 16289
rect 22192 16221 22244 16255
rect 21506 16181 21558 16197
rect 22192 16187 22200 16221
rect 22234 16187 22244 16221
rect 22192 16171 22244 16187
rect 22274 16289 22326 16301
rect 22274 16255 22284 16289
rect 22318 16255 22326 16289
rect 22274 16221 22326 16255
rect 22274 16187 22284 16221
rect 22318 16187 22326 16221
rect 23066 16291 23118 16303
rect 23066 16257 23074 16291
rect 23108 16257 23118 16291
rect 23066 16223 23118 16257
rect 23066 16189 23074 16223
rect 23108 16189 23118 16223
rect 22274 16171 22326 16187
rect 23066 16173 23118 16189
rect 23148 16291 23200 16303
rect 23148 16257 23158 16291
rect 23192 16257 23200 16291
rect 23148 16223 23200 16257
rect 23148 16189 23158 16223
rect 23192 16189 23200 16223
rect 23148 16173 23200 16189
rect 9887 16112 9903 16146
rect 9937 16112 9951 16146
rect 9887 16093 9951 16112
rect 4821 15457 4873 15475
rect 4625 15419 4681 15457
rect 4625 15385 4637 15419
rect 4671 15385 4681 15419
rect 4625 15373 4681 15385
rect 4711 15373 4765 15457
rect 4795 15391 4873 15457
rect 4795 15373 4829 15391
rect 4821 15357 4829 15373
rect 4863 15357 4873 15391
rect 4821 15345 4873 15357
rect 4903 15391 4959 15475
rect 4903 15357 4913 15391
rect 4947 15357 4959 15391
rect 4903 15345 4959 15357
rect 9687 15461 9739 15479
rect 9491 15423 9547 15461
rect 9491 15389 9503 15423
rect 9537 15389 9547 15423
rect 9491 15377 9547 15389
rect 9577 15377 9631 15461
rect 9661 15395 9739 15461
rect 9661 15377 9695 15395
rect 7050 15349 7143 15365
rect 7050 15319 7084 15349
rect 6635 15289 6687 15319
rect 6635 15255 6643 15289
rect 6677 15255 6687 15289
rect 6635 15235 6687 15255
rect 6717 15235 6775 15319
rect 6805 15235 6881 15319
rect 6911 15235 6977 15319
rect 7007 15315 7084 15319
rect 7118 15315 7143 15349
rect 7007 15281 7143 15315
rect 7007 15247 7084 15281
rect 7118 15247 7143 15281
rect 7007 15235 7143 15247
rect 7173 15349 7225 15365
rect 7173 15315 7183 15349
rect 7217 15315 7225 15349
rect 7173 15281 7225 15315
rect 7173 15247 7183 15281
rect 7217 15247 7225 15281
rect 9687 15361 9695 15377
rect 9729 15361 9739 15395
rect 9687 15349 9739 15361
rect 9769 15395 9825 15479
rect 9769 15361 9779 15395
rect 9813 15361 9825 15395
rect 9769 15349 9825 15361
rect 11916 15353 12009 15369
rect 11916 15323 11950 15353
rect 11501 15293 11553 15323
rect 11501 15259 11509 15293
rect 11543 15259 11553 15293
rect 7173 15235 7225 15247
rect 11501 15239 11553 15259
rect 11583 15239 11641 15323
rect 11671 15239 11747 15323
rect 11777 15239 11843 15323
rect 11873 15319 11950 15323
rect 11984 15319 12009 15353
rect 11873 15285 12009 15319
rect 11873 15251 11950 15285
rect 11984 15251 12009 15285
rect 11873 15239 12009 15251
rect 12039 15353 12091 15369
rect 12039 15319 12049 15353
rect 12083 15319 12091 15353
rect 12039 15285 12091 15319
rect 12039 15251 12049 15285
rect 12083 15251 12091 15285
rect 12039 15239 12091 15251
rect 6005 14847 6057 14865
rect 5809 14809 5865 14847
rect 5809 14775 5821 14809
rect 5855 14775 5865 14809
rect 5809 14763 5865 14775
rect 5895 14763 5949 14847
rect 5979 14781 6057 14847
rect 5979 14763 6013 14781
rect 6005 14747 6013 14763
rect 6047 14747 6057 14781
rect 6005 14735 6057 14747
rect 6087 14781 6143 14865
rect 6087 14747 6097 14781
rect 6131 14747 6143 14781
rect 10871 14851 10923 14869
rect 10675 14813 10731 14851
rect 10675 14779 10687 14813
rect 10721 14779 10731 14813
rect 10675 14767 10731 14779
rect 10761 14767 10815 14851
rect 10845 14785 10923 14851
rect 10845 14767 10879 14785
rect 6087 14735 6143 14747
rect 10871 14751 10879 14767
rect 10913 14751 10923 14785
rect 10871 14739 10923 14751
rect 10953 14785 11009 14869
rect 10953 14751 10963 14785
rect 10997 14751 11009 14785
rect 10953 14739 11009 14751
rect 4513 14573 4565 14655
rect 4513 14539 4521 14573
rect 4555 14539 4565 14573
rect 4513 14525 4565 14539
rect 4595 14595 4649 14655
rect 4595 14561 4605 14595
rect 4639 14561 4649 14595
rect 4595 14525 4649 14561
rect 4679 14573 4733 14655
rect 4679 14539 4689 14573
rect 4723 14539 4733 14573
rect 4679 14525 4733 14539
rect 4763 14525 4817 14655
rect 4847 14575 5001 14655
rect 4847 14541 4857 14575
rect 4891 14541 4957 14575
rect 4991 14541 5001 14575
rect 4847 14525 5001 14541
rect 5031 14646 5095 14655
rect 5031 14612 5047 14646
rect 5081 14612 5095 14646
rect 5031 14578 5095 14612
rect 5031 14544 5047 14578
rect 5081 14544 5095 14578
rect 9379 14577 9431 14659
rect 5031 14525 5095 14544
rect 9379 14543 9387 14577
rect 9421 14543 9431 14577
rect 9379 14529 9431 14543
rect 9461 14599 9515 14659
rect 9461 14565 9471 14599
rect 9505 14565 9515 14599
rect 9461 14529 9515 14565
rect 9545 14577 9599 14659
rect 9545 14543 9555 14577
rect 9589 14543 9599 14577
rect 9545 14529 9599 14543
rect 9629 14529 9683 14659
rect 9713 14579 9867 14659
rect 9713 14545 9723 14579
rect 9757 14545 9823 14579
rect 9857 14545 9867 14579
rect 9713 14529 9867 14545
rect 9897 14650 9961 14659
rect 9897 14616 9913 14650
rect 9947 14616 9961 14650
rect 9897 14582 9961 14616
rect 9897 14548 9913 14582
rect 9947 14548 9961 14582
rect 9897 14529 9961 14548
rect 23776 14441 23828 14453
rect 23776 14419 23784 14441
rect 23511 14390 23563 14419
rect 23511 14356 23519 14390
rect 23553 14356 23563 14390
rect 23511 14335 23563 14356
rect 23593 14381 23647 14419
rect 23593 14347 23603 14381
rect 23637 14347 23647 14381
rect 23593 14335 23647 14347
rect 23677 14335 23731 14419
rect 23761 14407 23784 14419
rect 23818 14407 23828 14441
rect 23761 14369 23828 14407
rect 23858 14415 23910 14453
rect 23858 14381 23868 14415
rect 23902 14381 23910 14415
rect 23858 14369 23910 14381
rect 23964 14424 24016 14462
rect 23964 14390 23972 14424
rect 24006 14390 24016 14424
rect 23964 14378 24016 14390
rect 24046 14433 24098 14462
rect 24046 14399 24056 14433
rect 24090 14399 24098 14433
rect 24046 14378 24098 14399
rect 24152 14431 24204 14469
rect 24152 14397 24160 14431
rect 24194 14397 24204 14431
rect 24152 14385 24204 14397
rect 24234 14457 24288 14469
rect 24234 14423 24244 14457
rect 24278 14423 24288 14457
rect 24234 14385 24288 14423
rect 24318 14457 24370 14469
rect 24318 14423 24328 14457
rect 24362 14423 24370 14457
rect 24318 14410 24370 14423
rect 25037 14419 25087 14469
rect 24318 14385 24368 14410
rect 24424 14393 24474 14419
rect 23761 14335 23811 14369
rect 24422 14381 24474 14393
rect 24422 14347 24430 14381
rect 24464 14347 24474 14381
rect 24422 14335 24474 14347
rect 24504 14381 24558 14419
rect 24504 14347 24514 14381
rect 24548 14347 24558 14381
rect 24504 14335 24558 14347
rect 24588 14397 24640 14419
rect 24588 14363 24598 14397
rect 24632 14363 24640 14397
rect 24588 14335 24640 14363
rect 24694 14381 24746 14419
rect 24694 14347 24702 14381
rect 24736 14347 24746 14381
rect 24694 14335 24746 14347
rect 24776 14403 24828 14419
rect 24776 14369 24786 14403
rect 24820 14369 24828 14403
rect 24776 14335 24828 14369
rect 24882 14389 24934 14419
rect 24882 14355 24890 14389
rect 24924 14355 24934 14389
rect 24882 14335 24934 14355
rect 24964 14389 25087 14419
rect 24964 14355 25030 14389
rect 25064 14385 25087 14389
rect 25117 14457 25169 14469
rect 25117 14423 25127 14457
rect 25161 14423 25169 14457
rect 25117 14385 25169 14423
rect 25064 14355 25072 14385
rect 24964 14335 25072 14355
rect 25255 14381 25307 14465
rect 25255 14347 25263 14381
rect 25297 14347 25307 14381
rect 25255 14335 25307 14347
rect 25337 14389 25389 14465
rect 25337 14355 25347 14389
rect 25381 14355 25389 14389
rect 25337 14335 25389 14355
rect 4831 13893 4883 13911
rect 4635 13855 4691 13893
rect 4635 13821 4647 13855
rect 4681 13821 4691 13855
rect 4635 13809 4691 13821
rect 4721 13809 4775 13893
rect 4805 13827 4883 13893
rect 4805 13809 4839 13827
rect 4831 13793 4839 13809
rect 4873 13793 4883 13827
rect 4831 13781 4883 13793
rect 4913 13827 4969 13911
rect 4913 13793 4923 13827
rect 4957 13793 4969 13827
rect 4913 13781 4969 13793
rect 6266 13883 6359 13899
rect 6266 13853 6300 13883
rect 5851 13823 5903 13853
rect 5851 13789 5859 13823
rect 5893 13789 5903 13823
rect 5851 13769 5903 13789
rect 5933 13769 5991 13853
rect 6021 13769 6097 13853
rect 6127 13769 6193 13853
rect 6223 13849 6300 13853
rect 6334 13849 6359 13883
rect 6223 13815 6359 13849
rect 6223 13781 6300 13815
rect 6334 13781 6359 13815
rect 6223 13769 6359 13781
rect 6389 13883 6441 13899
rect 6389 13849 6399 13883
rect 6433 13849 6441 13883
rect 6389 13815 6441 13849
rect 6389 13781 6399 13815
rect 6433 13781 6441 13815
rect 6389 13769 6441 13781
rect 9697 13897 9749 13915
rect 8110 13843 8163 13883
rect 7749 13823 7801 13843
rect 7749 13789 7757 13823
rect 7791 13789 7801 13823
rect 7749 13759 7801 13789
rect 7831 13817 7897 13843
rect 7831 13783 7847 13817
rect 7881 13783 7897 13817
rect 7831 13759 7897 13783
rect 7927 13803 7981 13843
rect 7927 13769 7937 13803
rect 7971 13769 7981 13803
rect 7927 13759 7981 13769
rect 8011 13817 8065 13843
rect 8011 13783 8021 13817
rect 8055 13783 8065 13817
rect 8011 13759 8065 13783
rect 8095 13803 8163 13843
rect 8095 13769 8115 13803
rect 8149 13769 8163 13803
rect 8095 13759 8163 13769
rect 8110 13753 8163 13759
rect 8193 13841 8247 13883
rect 8193 13807 8203 13841
rect 8237 13807 8247 13841
rect 8193 13753 8247 13807
rect 9501 13859 9557 13897
rect 9501 13825 9513 13859
rect 9547 13825 9557 13859
rect 9501 13813 9557 13825
rect 9587 13813 9641 13897
rect 9671 13831 9749 13897
rect 9671 13813 9705 13831
rect 9697 13797 9705 13813
rect 9739 13797 9749 13831
rect 9697 13785 9749 13797
rect 9779 13831 9835 13915
rect 9779 13797 9789 13831
rect 9823 13797 9835 13831
rect 9779 13785 9835 13797
rect 11132 13887 11225 13903
rect 11132 13857 11166 13887
rect 10717 13827 10769 13857
rect 10717 13793 10725 13827
rect 10759 13793 10769 13827
rect 10717 13773 10769 13793
rect 10799 13773 10857 13857
rect 10887 13773 10963 13857
rect 10993 13773 11059 13857
rect 11089 13853 11166 13857
rect 11200 13853 11225 13887
rect 11089 13819 11225 13853
rect 11089 13785 11166 13819
rect 11200 13785 11225 13819
rect 11089 13773 11225 13785
rect 11255 13887 11307 13903
rect 11255 13853 11265 13887
rect 11299 13853 11307 13887
rect 11255 13819 11307 13853
rect 11255 13785 11265 13819
rect 11299 13785 11307 13819
rect 11255 13773 11307 13785
rect 12976 13847 13029 13887
rect 12615 13827 12667 13847
rect 12615 13793 12623 13827
rect 12657 13793 12667 13827
rect 12615 13763 12667 13793
rect 12697 13821 12763 13847
rect 12697 13787 12713 13821
rect 12747 13787 12763 13821
rect 12697 13763 12763 13787
rect 12793 13807 12847 13847
rect 12793 13773 12803 13807
rect 12837 13773 12847 13807
rect 12793 13763 12847 13773
rect 12877 13821 12931 13847
rect 12877 13787 12887 13821
rect 12921 13787 12931 13821
rect 12877 13763 12931 13787
rect 12961 13807 13029 13847
rect 12961 13773 12981 13807
rect 13015 13773 13029 13807
rect 12961 13763 13029 13773
rect 12976 13757 13029 13763
rect 13059 13845 13113 13887
rect 13059 13811 13069 13845
rect 13103 13811 13113 13845
rect 13059 13757 13113 13811
rect 7031 13479 7083 13525
rect 6850 13451 6902 13479
rect 6850 13417 6858 13451
rect 6892 13417 6902 13451
rect 6850 13395 6902 13417
rect 6932 13451 6986 13479
rect 6932 13417 6942 13451
rect 6976 13417 6986 13451
rect 6932 13395 6986 13417
rect 7016 13451 7083 13479
rect 7016 13417 7038 13451
rect 7072 13417 7083 13451
rect 7016 13395 7083 13417
rect 7113 13511 7165 13525
rect 7113 13477 7123 13511
rect 7157 13477 7165 13511
rect 7113 13443 7165 13477
rect 7113 13409 7123 13443
rect 7157 13409 7165 13443
rect 11897 13483 11949 13529
rect 11716 13455 11768 13483
rect 11716 13421 11724 13455
rect 11758 13421 11768 13455
rect 7113 13395 7165 13409
rect 11716 13399 11768 13421
rect 11798 13455 11852 13483
rect 11798 13421 11808 13455
rect 11842 13421 11852 13455
rect 11798 13399 11852 13421
rect 11882 13455 11949 13483
rect 11882 13421 11904 13455
rect 11938 13421 11949 13455
rect 11882 13399 11949 13421
rect 11979 13515 12031 13529
rect 11979 13481 11989 13515
rect 12023 13481 12031 13515
rect 11979 13447 12031 13481
rect 11979 13413 11989 13447
rect 12023 13413 12031 13447
rect 11979 13399 12031 13413
rect 6249 13011 6299 13057
rect 4505 12905 4557 12987
rect 4505 12871 4513 12905
rect 4547 12871 4557 12905
rect 4505 12857 4557 12871
rect 4587 12927 4641 12987
rect 4587 12893 4597 12927
rect 4631 12893 4641 12927
rect 4587 12857 4641 12893
rect 4671 12905 4725 12987
rect 4671 12871 4681 12905
rect 4715 12871 4725 12905
rect 4671 12857 4725 12871
rect 4755 12857 4809 12987
rect 4839 12907 4993 12987
rect 4839 12873 4849 12907
rect 4883 12873 4949 12907
rect 4983 12873 4993 12907
rect 4839 12857 4993 12873
rect 5023 12978 5087 12987
rect 5023 12944 5039 12978
rect 5073 12944 5087 12978
rect 5975 12973 6027 13011
rect 5023 12910 5087 12944
rect 5975 12939 5983 12973
rect 6017 12939 6027 12973
rect 5975 12927 6027 12939
rect 6057 12927 6099 13011
rect 6129 12927 6171 13011
rect 6201 12989 6299 13011
rect 6201 12955 6255 12989
rect 6289 12955 6299 12989
rect 6201 12927 6299 12955
rect 6329 12999 6381 13057
rect 6329 12965 6339 12999
rect 6373 12965 6381 12999
rect 11115 13015 11165 13061
rect 6329 12927 6381 12965
rect 5023 12876 5039 12910
rect 5073 12876 5087 12910
rect 9371 12909 9423 12991
rect 5023 12857 5087 12876
rect 9371 12875 9379 12909
rect 9413 12875 9423 12909
rect 9371 12861 9423 12875
rect 9453 12931 9507 12991
rect 9453 12897 9463 12931
rect 9497 12897 9507 12931
rect 9453 12861 9507 12897
rect 9537 12909 9591 12991
rect 9537 12875 9547 12909
rect 9581 12875 9591 12909
rect 9537 12861 9591 12875
rect 9621 12861 9675 12991
rect 9705 12911 9859 12991
rect 9705 12877 9715 12911
rect 9749 12877 9815 12911
rect 9849 12877 9859 12911
rect 9705 12861 9859 12877
rect 9889 12982 9953 12991
rect 9889 12948 9905 12982
rect 9939 12948 9953 12982
rect 10841 12977 10893 13015
rect 9889 12914 9953 12948
rect 10841 12943 10849 12977
rect 10883 12943 10893 12977
rect 10841 12931 10893 12943
rect 10923 12931 10965 13015
rect 10995 12931 11037 13015
rect 11067 12993 11165 13015
rect 11067 12959 11121 12993
rect 11155 12959 11165 12993
rect 11067 12931 11165 12959
rect 11195 13003 11247 13061
rect 11195 12969 11205 13003
rect 11239 12969 11247 13003
rect 11195 12931 11247 12969
rect 9889 12880 9905 12914
rect 9939 12880 9953 12914
rect 9889 12861 9953 12880
rect 4823 12225 4875 12243
rect 4627 12187 4683 12225
rect 4627 12153 4639 12187
rect 4673 12153 4683 12187
rect 4627 12141 4683 12153
rect 4713 12141 4767 12225
rect 4797 12159 4875 12225
rect 4797 12141 4831 12159
rect 4823 12125 4831 12141
rect 4865 12125 4875 12159
rect 4823 12113 4875 12125
rect 4905 12159 4961 12243
rect 4905 12125 4915 12159
rect 4949 12125 4961 12159
rect 4905 12113 4961 12125
rect 9689 12229 9741 12247
rect 9493 12191 9549 12229
rect 9493 12157 9505 12191
rect 9539 12157 9549 12191
rect 9493 12145 9549 12157
rect 9579 12145 9633 12229
rect 9663 12163 9741 12229
rect 9663 12145 9697 12163
rect 9689 12129 9697 12145
rect 9731 12129 9741 12163
rect 9689 12117 9741 12129
rect 9771 12163 9827 12247
rect 9771 12129 9781 12163
rect 9815 12129 9827 12163
rect 9771 12117 9827 12129
rect 6199 12019 6251 12037
rect 6003 11981 6059 12019
rect 6003 11947 6015 11981
rect 6049 11947 6059 11981
rect 6003 11935 6059 11947
rect 6089 11935 6143 12019
rect 6173 11953 6251 12019
rect 6173 11935 6207 11953
rect 6199 11919 6207 11935
rect 6241 11919 6251 11953
rect 6199 11907 6251 11919
rect 6281 11953 6337 12037
rect 6281 11919 6291 11953
rect 6325 11919 6337 11953
rect 11065 12023 11117 12041
rect 10869 11985 10925 12023
rect 10869 11951 10881 11985
rect 10915 11951 10925 11985
rect 10869 11939 10925 11951
rect 10955 11939 11009 12023
rect 11039 11957 11117 12023
rect 11039 11939 11073 11957
rect 6281 11907 6337 11919
rect 11065 11923 11073 11939
rect 11107 11923 11117 11957
rect 11065 11911 11117 11923
rect 11147 11957 11203 12041
rect 11147 11923 11157 11957
rect 11191 11923 11203 11957
rect 11147 11911 11203 11923
rect 4515 11341 4567 11423
rect 4515 11307 4523 11341
rect 4557 11307 4567 11341
rect 4515 11293 4567 11307
rect 4597 11363 4651 11423
rect 4597 11329 4607 11363
rect 4641 11329 4651 11363
rect 4597 11293 4651 11329
rect 4681 11341 4735 11423
rect 4681 11307 4691 11341
rect 4725 11307 4735 11341
rect 4681 11293 4735 11307
rect 4765 11293 4819 11423
rect 4849 11343 5003 11423
rect 4849 11309 4859 11343
rect 4893 11309 4959 11343
rect 4993 11309 5003 11343
rect 4849 11293 5003 11309
rect 5033 11414 5097 11423
rect 5033 11380 5049 11414
rect 5083 11380 5097 11414
rect 5033 11346 5097 11380
rect 5033 11312 5049 11346
rect 5083 11312 5097 11346
rect 9381 11345 9433 11427
rect 5033 11293 5097 11312
rect 9381 11311 9389 11345
rect 9423 11311 9433 11345
rect 9381 11297 9433 11311
rect 9463 11367 9517 11427
rect 9463 11333 9473 11367
rect 9507 11333 9517 11367
rect 9463 11297 9517 11333
rect 9547 11345 9601 11427
rect 9547 11311 9557 11345
rect 9591 11311 9601 11345
rect 9547 11297 9601 11311
rect 9631 11297 9685 11427
rect 9715 11347 9869 11427
rect 9715 11313 9725 11347
rect 9759 11313 9825 11347
rect 9859 11313 9869 11347
rect 9715 11297 9869 11313
rect 9899 11418 9963 11427
rect 9899 11384 9915 11418
rect 9949 11384 9963 11418
rect 9899 11350 9963 11384
rect 9899 11316 9915 11350
rect 9949 11316 9963 11350
rect 9899 11297 9963 11316
rect 4833 10661 4885 10679
rect 4637 10623 4693 10661
rect 4637 10589 4649 10623
rect 4683 10589 4693 10623
rect 4637 10577 4693 10589
rect 4723 10577 4777 10661
rect 4807 10595 4885 10661
rect 4807 10577 4841 10595
rect 4833 10561 4841 10577
rect 4875 10561 4885 10595
rect 4833 10549 4885 10561
rect 4915 10595 4971 10679
rect 4915 10561 4925 10595
rect 4959 10561 4971 10595
rect 9699 10665 9751 10683
rect 9503 10627 9559 10665
rect 9503 10593 9515 10627
rect 9549 10593 9559 10627
rect 9503 10581 9559 10593
rect 9589 10581 9643 10665
rect 9673 10599 9751 10665
rect 9673 10581 9707 10599
rect 4915 10549 4971 10561
rect 9699 10565 9707 10581
rect 9741 10565 9751 10599
rect 9699 10553 9751 10565
rect 9781 10599 9837 10683
rect 9781 10565 9791 10599
rect 9825 10565 9837 10599
rect 9781 10553 9837 10565
rect 6186 6537 6238 6553
rect 6186 6503 6194 6537
rect 6228 6503 6238 6537
rect 6186 6469 6238 6503
rect 6186 6435 6194 6469
rect 6228 6435 6238 6469
rect 6186 6423 6238 6435
rect 6268 6537 6320 6553
rect 6268 6503 6278 6537
rect 6312 6503 6320 6537
rect 6268 6469 6320 6503
rect 6268 6435 6278 6469
rect 6312 6435 6320 6469
rect 6268 6423 6320 6435
rect 10080 5873 10132 5921
rect 10080 5839 10088 5873
rect 10122 5839 10132 5873
rect 10080 5791 10132 5839
rect 10162 5913 10231 5921
rect 10162 5879 10187 5913
rect 10221 5879 10231 5913
rect 10162 5837 10231 5879
rect 10261 5837 10327 5921
rect 10357 5837 10399 5921
rect 10429 5901 10495 5921
rect 10429 5867 10439 5901
rect 10473 5867 10495 5901
rect 10429 5837 10495 5867
rect 10525 5896 10584 5921
rect 10525 5862 10540 5896
rect 10574 5862 10584 5896
rect 10525 5837 10584 5862
rect 10614 5913 10668 5921
rect 10614 5879 10624 5913
rect 10658 5879 10668 5913
rect 10614 5837 10668 5879
rect 10698 5896 10752 5921
rect 10698 5862 10708 5896
rect 10742 5862 10752 5896
rect 10698 5837 10752 5862
rect 10782 5904 10834 5921
rect 10782 5870 10792 5904
rect 10826 5870 10834 5904
rect 10782 5837 10834 5870
rect 10888 5896 10940 5921
rect 10888 5862 10896 5896
rect 10930 5862 10940 5896
rect 10888 5837 10940 5862
rect 10970 5913 11024 5921
rect 10970 5879 10980 5913
rect 11014 5879 11024 5913
rect 10970 5837 11024 5879
rect 11054 5896 11108 5921
rect 11054 5862 11064 5896
rect 11098 5862 11108 5896
rect 11054 5837 11108 5862
rect 11138 5896 11192 5921
rect 11138 5862 11148 5896
rect 11182 5862 11192 5896
rect 11138 5837 11192 5862
rect 11222 5837 11282 5921
rect 11312 5909 11381 5921
rect 11312 5875 11337 5909
rect 11371 5875 11381 5909
rect 11312 5837 11381 5875
rect 10162 5791 10214 5837
rect 1898 5453 1950 5501
rect 1898 5419 1906 5453
rect 1940 5419 1950 5453
rect 1898 5371 1950 5419
rect 1980 5493 2049 5501
rect 1980 5459 2005 5493
rect 2039 5459 2049 5493
rect 1980 5417 2049 5459
rect 2079 5417 2145 5501
rect 2175 5417 2217 5501
rect 2247 5481 2313 5501
rect 2247 5447 2257 5481
rect 2291 5447 2313 5481
rect 2247 5417 2313 5447
rect 2343 5476 2402 5501
rect 2343 5442 2358 5476
rect 2392 5442 2402 5476
rect 2343 5417 2402 5442
rect 2432 5493 2486 5501
rect 2432 5459 2442 5493
rect 2476 5459 2486 5493
rect 2432 5417 2486 5459
rect 2516 5476 2570 5501
rect 2516 5442 2526 5476
rect 2560 5442 2570 5476
rect 2516 5417 2570 5442
rect 2600 5484 2652 5501
rect 2600 5450 2610 5484
rect 2644 5450 2652 5484
rect 2600 5417 2652 5450
rect 2706 5476 2758 5501
rect 2706 5442 2714 5476
rect 2748 5442 2758 5476
rect 2706 5417 2758 5442
rect 2788 5493 2842 5501
rect 2788 5459 2798 5493
rect 2832 5459 2842 5493
rect 2788 5417 2842 5459
rect 2872 5476 2926 5501
rect 2872 5442 2882 5476
rect 2916 5442 2926 5476
rect 2872 5417 2926 5442
rect 2956 5476 3010 5501
rect 2956 5442 2966 5476
rect 3000 5442 3010 5476
rect 2956 5417 3010 5442
rect 3040 5417 3100 5501
rect 3130 5489 3199 5501
rect 3130 5455 3155 5489
rect 3189 5455 3199 5489
rect 3130 5417 3199 5455
rect 1980 5371 2032 5417
rect 3147 5371 3199 5417
rect 3229 5453 3281 5501
rect 3229 5419 3239 5453
rect 3273 5419 3281 5453
rect 3229 5371 3281 5419
rect 4032 5445 4084 5493
rect 4032 5411 4040 5445
rect 4074 5411 4084 5445
rect 4032 5363 4084 5411
rect 4114 5485 4183 5493
rect 4114 5451 4139 5485
rect 4173 5451 4183 5485
rect 4114 5409 4183 5451
rect 4213 5409 4279 5493
rect 4309 5409 4351 5493
rect 4381 5473 4447 5493
rect 4381 5439 4391 5473
rect 4425 5439 4447 5473
rect 4381 5409 4447 5439
rect 4477 5468 4536 5493
rect 4477 5434 4492 5468
rect 4526 5434 4536 5468
rect 4477 5409 4536 5434
rect 4566 5485 4620 5493
rect 4566 5451 4576 5485
rect 4610 5451 4620 5485
rect 4566 5409 4620 5451
rect 4650 5468 4704 5493
rect 4650 5434 4660 5468
rect 4694 5434 4704 5468
rect 4650 5409 4704 5434
rect 4734 5476 4786 5493
rect 4734 5442 4744 5476
rect 4778 5442 4786 5476
rect 4734 5409 4786 5442
rect 4840 5468 4892 5493
rect 4840 5434 4848 5468
rect 4882 5434 4892 5468
rect 4840 5409 4892 5434
rect 4922 5485 4976 5493
rect 4922 5451 4932 5485
rect 4966 5451 4976 5485
rect 4922 5409 4976 5451
rect 5006 5468 5060 5493
rect 5006 5434 5016 5468
rect 5050 5434 5060 5468
rect 5006 5409 5060 5434
rect 5090 5468 5144 5493
rect 5090 5434 5100 5468
rect 5134 5434 5144 5468
rect 5090 5409 5144 5434
rect 5174 5409 5234 5493
rect 5264 5481 5333 5493
rect 5264 5447 5289 5481
rect 5323 5447 5333 5481
rect 5264 5409 5333 5447
rect 4114 5363 4166 5409
rect 5281 5363 5333 5409
rect 5363 5445 5415 5493
rect 5363 5411 5373 5445
rect 5407 5411 5415 5445
rect 5363 5363 5415 5411
rect 5984 5445 6036 5493
rect 5984 5411 5992 5445
rect 6026 5411 6036 5445
rect 5984 5363 6036 5411
rect 6066 5485 6135 5493
rect 6066 5451 6091 5485
rect 6125 5451 6135 5485
rect 6066 5409 6135 5451
rect 6165 5409 6231 5493
rect 6261 5409 6303 5493
rect 6333 5473 6399 5493
rect 6333 5439 6343 5473
rect 6377 5439 6399 5473
rect 6333 5409 6399 5439
rect 6429 5468 6488 5493
rect 6429 5434 6444 5468
rect 6478 5434 6488 5468
rect 6429 5409 6488 5434
rect 6518 5485 6572 5493
rect 6518 5451 6528 5485
rect 6562 5451 6572 5485
rect 6518 5409 6572 5451
rect 6602 5468 6656 5493
rect 6602 5434 6612 5468
rect 6646 5434 6656 5468
rect 6602 5409 6656 5434
rect 6686 5476 6738 5493
rect 6686 5442 6696 5476
rect 6730 5442 6738 5476
rect 6686 5409 6738 5442
rect 6792 5468 6844 5493
rect 6792 5434 6800 5468
rect 6834 5434 6844 5468
rect 6792 5409 6844 5434
rect 6874 5485 6928 5493
rect 6874 5451 6884 5485
rect 6918 5451 6928 5485
rect 6874 5409 6928 5451
rect 6958 5468 7012 5493
rect 6958 5434 6968 5468
rect 7002 5434 7012 5468
rect 6958 5409 7012 5434
rect 7042 5468 7096 5493
rect 7042 5434 7052 5468
rect 7086 5434 7096 5468
rect 7042 5409 7096 5434
rect 7126 5409 7186 5493
rect 7216 5481 7285 5493
rect 7216 5447 7241 5481
rect 7275 5447 7285 5481
rect 7216 5409 7285 5447
rect 6066 5363 6118 5409
rect 7233 5363 7285 5409
rect 7315 5445 7367 5493
rect 7315 5411 7325 5445
rect 7359 5411 7367 5445
rect 7315 5363 7367 5411
rect 7986 5451 8038 5499
rect 7986 5417 7994 5451
rect 8028 5417 8038 5451
rect 7986 5369 8038 5417
rect 8068 5491 8137 5499
rect 8068 5457 8093 5491
rect 8127 5457 8137 5491
rect 8068 5415 8137 5457
rect 8167 5415 8233 5499
rect 8263 5415 8305 5499
rect 8335 5479 8401 5499
rect 8335 5445 8345 5479
rect 8379 5445 8401 5479
rect 8335 5415 8401 5445
rect 8431 5474 8490 5499
rect 8431 5440 8446 5474
rect 8480 5440 8490 5474
rect 8431 5415 8490 5440
rect 8520 5491 8574 5499
rect 8520 5457 8530 5491
rect 8564 5457 8574 5491
rect 8520 5415 8574 5457
rect 8604 5474 8658 5499
rect 8604 5440 8614 5474
rect 8648 5440 8658 5474
rect 8604 5415 8658 5440
rect 8688 5482 8740 5499
rect 8688 5448 8698 5482
rect 8732 5448 8740 5482
rect 8688 5415 8740 5448
rect 8794 5474 8846 5499
rect 8794 5440 8802 5474
rect 8836 5440 8846 5474
rect 8794 5415 8846 5440
rect 8876 5491 8930 5499
rect 8876 5457 8886 5491
rect 8920 5457 8930 5491
rect 8876 5415 8930 5457
rect 8960 5474 9014 5499
rect 8960 5440 8970 5474
rect 9004 5440 9014 5474
rect 8960 5415 9014 5440
rect 9044 5474 9098 5499
rect 9044 5440 9054 5474
rect 9088 5440 9098 5474
rect 9044 5415 9098 5440
rect 9128 5415 9188 5499
rect 9218 5487 9287 5499
rect 9218 5453 9243 5487
rect 9277 5453 9287 5487
rect 9218 5415 9287 5453
rect 8068 5369 8120 5415
rect 9235 5369 9287 5415
rect 9317 5451 9369 5499
rect 11329 5791 11381 5837
rect 11411 5873 11463 5921
rect 11411 5839 11421 5873
rect 11455 5839 11463 5873
rect 11411 5791 11463 5839
rect 12142 5861 12194 5909
rect 12142 5827 12150 5861
rect 12184 5827 12194 5861
rect 12142 5779 12194 5827
rect 12224 5901 12293 5909
rect 12224 5867 12249 5901
rect 12283 5867 12293 5901
rect 12224 5825 12293 5867
rect 12323 5825 12389 5909
rect 12419 5825 12461 5909
rect 12491 5889 12557 5909
rect 12491 5855 12501 5889
rect 12535 5855 12557 5889
rect 12491 5825 12557 5855
rect 12587 5884 12646 5909
rect 12587 5850 12602 5884
rect 12636 5850 12646 5884
rect 12587 5825 12646 5850
rect 12676 5901 12730 5909
rect 12676 5867 12686 5901
rect 12720 5867 12730 5901
rect 12676 5825 12730 5867
rect 12760 5884 12814 5909
rect 12760 5850 12770 5884
rect 12804 5850 12814 5884
rect 12760 5825 12814 5850
rect 12844 5892 12896 5909
rect 12844 5858 12854 5892
rect 12888 5858 12896 5892
rect 12844 5825 12896 5858
rect 12950 5884 13002 5909
rect 12950 5850 12958 5884
rect 12992 5850 13002 5884
rect 12950 5825 13002 5850
rect 13032 5901 13086 5909
rect 13032 5867 13042 5901
rect 13076 5867 13086 5901
rect 13032 5825 13086 5867
rect 13116 5884 13170 5909
rect 13116 5850 13126 5884
rect 13160 5850 13170 5884
rect 13116 5825 13170 5850
rect 13200 5884 13254 5909
rect 13200 5850 13210 5884
rect 13244 5850 13254 5884
rect 13200 5825 13254 5850
rect 13284 5825 13344 5909
rect 13374 5897 13443 5909
rect 13374 5863 13399 5897
rect 13433 5863 13443 5897
rect 13374 5825 13443 5863
rect 12224 5779 12276 5825
rect 9317 5417 9327 5451
rect 9361 5417 9369 5451
rect 13391 5779 13443 5825
rect 13473 5861 13525 5909
rect 13473 5827 13483 5861
rect 13517 5827 13525 5861
rect 13473 5779 13525 5827
rect 14100 5869 14152 5917
rect 14100 5835 14108 5869
rect 14142 5835 14152 5869
rect 14100 5787 14152 5835
rect 14182 5909 14251 5917
rect 14182 5875 14207 5909
rect 14241 5875 14251 5909
rect 14182 5833 14251 5875
rect 14281 5833 14347 5917
rect 14377 5833 14419 5917
rect 14449 5897 14515 5917
rect 14449 5863 14459 5897
rect 14493 5863 14515 5897
rect 14449 5833 14515 5863
rect 14545 5892 14604 5917
rect 14545 5858 14560 5892
rect 14594 5858 14604 5892
rect 14545 5833 14604 5858
rect 14634 5909 14688 5917
rect 14634 5875 14644 5909
rect 14678 5875 14688 5909
rect 14634 5833 14688 5875
rect 14718 5892 14772 5917
rect 14718 5858 14728 5892
rect 14762 5858 14772 5892
rect 14718 5833 14772 5858
rect 14802 5900 14854 5917
rect 14802 5866 14812 5900
rect 14846 5866 14854 5900
rect 14802 5833 14854 5866
rect 14908 5892 14960 5917
rect 14908 5858 14916 5892
rect 14950 5858 14960 5892
rect 14908 5833 14960 5858
rect 14990 5909 15044 5917
rect 14990 5875 15000 5909
rect 15034 5875 15044 5909
rect 14990 5833 15044 5875
rect 15074 5892 15128 5917
rect 15074 5858 15084 5892
rect 15118 5858 15128 5892
rect 15074 5833 15128 5858
rect 15158 5892 15212 5917
rect 15158 5858 15168 5892
rect 15202 5858 15212 5892
rect 15158 5833 15212 5858
rect 15242 5833 15302 5917
rect 15332 5905 15401 5917
rect 15332 5871 15357 5905
rect 15391 5871 15401 5905
rect 15332 5833 15401 5871
rect 14182 5787 14234 5833
rect 15349 5787 15401 5833
rect 15431 5869 15483 5917
rect 15431 5835 15441 5869
rect 15475 5835 15483 5869
rect 15431 5787 15483 5835
rect 16094 5875 16146 5923
rect 16094 5841 16102 5875
rect 16136 5841 16146 5875
rect 16094 5793 16146 5841
rect 16176 5915 16245 5923
rect 16176 5881 16201 5915
rect 16235 5881 16245 5915
rect 16176 5839 16245 5881
rect 16275 5839 16341 5923
rect 16371 5839 16413 5923
rect 16443 5903 16509 5923
rect 16443 5869 16453 5903
rect 16487 5869 16509 5903
rect 16443 5839 16509 5869
rect 16539 5898 16598 5923
rect 16539 5864 16554 5898
rect 16588 5864 16598 5898
rect 16539 5839 16598 5864
rect 16628 5915 16682 5923
rect 16628 5881 16638 5915
rect 16672 5881 16682 5915
rect 16628 5839 16682 5881
rect 16712 5898 16766 5923
rect 16712 5864 16722 5898
rect 16756 5864 16766 5898
rect 16712 5839 16766 5864
rect 16796 5906 16848 5923
rect 16796 5872 16806 5906
rect 16840 5872 16848 5906
rect 16796 5839 16848 5872
rect 16902 5898 16954 5923
rect 16902 5864 16910 5898
rect 16944 5864 16954 5898
rect 16902 5839 16954 5864
rect 16984 5915 17038 5923
rect 16984 5881 16994 5915
rect 17028 5881 17038 5915
rect 16984 5839 17038 5881
rect 17068 5898 17122 5923
rect 17068 5864 17078 5898
rect 17112 5864 17122 5898
rect 17068 5839 17122 5864
rect 17152 5898 17206 5923
rect 17152 5864 17162 5898
rect 17196 5864 17206 5898
rect 17152 5839 17206 5864
rect 17236 5839 17296 5923
rect 17326 5911 17395 5923
rect 17326 5877 17351 5911
rect 17385 5877 17395 5911
rect 17326 5839 17395 5877
rect 16176 5793 16228 5839
rect 17343 5793 17395 5839
rect 17425 5875 17477 5923
rect 17425 5841 17435 5875
rect 17469 5841 17477 5875
rect 17425 5793 17477 5841
rect 9317 5369 9369 5417
rect 18375 5322 18427 5349
rect 18375 5288 18383 5322
rect 18417 5288 18427 5322
rect 18375 5265 18427 5288
rect 18457 5322 18595 5349
rect 18457 5288 18467 5322
rect 18501 5288 18535 5322
rect 18569 5288 18595 5322
rect 18457 5265 18595 5288
rect 18625 5265 18691 5349
rect 18721 5322 18816 5349
rect 18721 5288 18770 5322
rect 18804 5288 18816 5322
rect 18721 5265 18816 5288
rect 18846 5265 18912 5349
rect 18942 5337 19021 5349
rect 18942 5303 18977 5337
rect 19011 5303 19021 5337
rect 18942 5265 19021 5303
rect 10108 4999 10160 5047
rect 10108 4965 10116 4999
rect 10150 4965 10160 4999
rect 10108 4917 10160 4965
rect 10190 5039 10259 5047
rect 10190 5005 10215 5039
rect 10249 5005 10259 5039
rect 10190 4963 10259 5005
rect 10289 4963 10355 5047
rect 10385 4963 10427 5047
rect 10457 5027 10523 5047
rect 10457 4993 10467 5027
rect 10501 4993 10523 5027
rect 10457 4963 10523 4993
rect 10553 5022 10612 5047
rect 10553 4988 10568 5022
rect 10602 4988 10612 5022
rect 10553 4963 10612 4988
rect 10642 5039 10696 5047
rect 10642 5005 10652 5039
rect 10686 5005 10696 5039
rect 10642 4963 10696 5005
rect 10726 5022 10780 5047
rect 10726 4988 10736 5022
rect 10770 4988 10780 5022
rect 10726 4963 10780 4988
rect 10810 5030 10862 5047
rect 10810 4996 10820 5030
rect 10854 4996 10862 5030
rect 10810 4963 10862 4996
rect 10916 5022 10968 5047
rect 10916 4988 10924 5022
rect 10958 4988 10968 5022
rect 10916 4963 10968 4988
rect 10998 5039 11052 5047
rect 10998 5005 11008 5039
rect 11042 5005 11052 5039
rect 10998 4963 11052 5005
rect 11082 5022 11136 5047
rect 11082 4988 11092 5022
rect 11126 4988 11136 5022
rect 11082 4963 11136 4988
rect 11166 5022 11220 5047
rect 11166 4988 11176 5022
rect 11210 4988 11220 5022
rect 11166 4963 11220 4988
rect 11250 4963 11310 5047
rect 11340 5035 11409 5047
rect 11340 5001 11365 5035
rect 11399 5001 11409 5035
rect 11340 4963 11409 5001
rect 10190 4917 10242 4963
rect 11357 4917 11409 4963
rect 11439 4999 11491 5047
rect 11439 4965 11449 4999
rect 11483 4965 11491 4999
rect 11439 4917 11491 4965
rect 12378 4955 12430 5003
rect 12378 4921 12386 4955
rect 12420 4921 12430 4955
rect 12378 4873 12430 4921
rect 12460 4995 12529 5003
rect 12460 4961 12485 4995
rect 12519 4961 12529 4995
rect 12460 4919 12529 4961
rect 12559 4919 12625 5003
rect 12655 4919 12697 5003
rect 12727 4983 12793 5003
rect 12727 4949 12737 4983
rect 12771 4949 12793 4983
rect 12727 4919 12793 4949
rect 12823 4978 12882 5003
rect 12823 4944 12838 4978
rect 12872 4944 12882 4978
rect 12823 4919 12882 4944
rect 12912 4995 12966 5003
rect 12912 4961 12922 4995
rect 12956 4961 12966 4995
rect 12912 4919 12966 4961
rect 12996 4978 13050 5003
rect 12996 4944 13006 4978
rect 13040 4944 13050 4978
rect 12996 4919 13050 4944
rect 13080 4986 13132 5003
rect 13080 4952 13090 4986
rect 13124 4952 13132 4986
rect 13080 4919 13132 4952
rect 13186 4978 13238 5003
rect 13186 4944 13194 4978
rect 13228 4944 13238 4978
rect 13186 4919 13238 4944
rect 13268 4995 13322 5003
rect 13268 4961 13278 4995
rect 13312 4961 13322 4995
rect 13268 4919 13322 4961
rect 13352 4978 13406 5003
rect 13352 4944 13362 4978
rect 13396 4944 13406 4978
rect 13352 4919 13406 4944
rect 13436 4978 13490 5003
rect 13436 4944 13446 4978
rect 13480 4944 13490 4978
rect 13436 4919 13490 4944
rect 13520 4919 13580 5003
rect 13610 4991 13679 5003
rect 13610 4957 13635 4991
rect 13669 4957 13679 4991
rect 13610 4919 13679 4957
rect 12460 4873 12512 4919
rect 13627 4873 13679 4919
rect 13709 4955 13761 5003
rect 18969 5219 19021 5265
rect 19051 5318 19103 5349
rect 19051 5284 19061 5318
rect 19095 5284 19103 5318
rect 19051 5219 19103 5284
rect 13709 4921 13719 4955
rect 13753 4921 13761 4955
rect 13709 4873 13761 4921
rect 14380 4949 14432 4997
rect 14380 4915 14388 4949
rect 14422 4915 14432 4949
rect 14380 4867 14432 4915
rect 14462 4989 14531 4997
rect 14462 4955 14487 4989
rect 14521 4955 14531 4989
rect 14462 4913 14531 4955
rect 14561 4913 14627 4997
rect 14657 4913 14699 4997
rect 14729 4977 14795 4997
rect 14729 4943 14739 4977
rect 14773 4943 14795 4977
rect 14729 4913 14795 4943
rect 14825 4972 14884 4997
rect 14825 4938 14840 4972
rect 14874 4938 14884 4972
rect 14825 4913 14884 4938
rect 14914 4989 14968 4997
rect 14914 4955 14924 4989
rect 14958 4955 14968 4989
rect 14914 4913 14968 4955
rect 14998 4972 15052 4997
rect 14998 4938 15008 4972
rect 15042 4938 15052 4972
rect 14998 4913 15052 4938
rect 15082 4980 15134 4997
rect 15082 4946 15092 4980
rect 15126 4946 15134 4980
rect 15082 4913 15134 4946
rect 15188 4972 15240 4997
rect 15188 4938 15196 4972
rect 15230 4938 15240 4972
rect 15188 4913 15240 4938
rect 15270 4989 15324 4997
rect 15270 4955 15280 4989
rect 15314 4955 15324 4989
rect 15270 4913 15324 4955
rect 15354 4972 15408 4997
rect 15354 4938 15364 4972
rect 15398 4938 15408 4972
rect 15354 4913 15408 4938
rect 15438 4972 15492 4997
rect 15438 4938 15448 4972
rect 15482 4938 15492 4972
rect 15438 4913 15492 4938
rect 15522 4913 15582 4997
rect 15612 4985 15681 4997
rect 15612 4951 15637 4985
rect 15671 4951 15681 4985
rect 15612 4913 15681 4951
rect 14462 4867 14514 4913
rect 15629 4867 15681 4913
rect 15711 4949 15763 4997
rect 15711 4915 15721 4949
rect 15755 4915 15763 4949
rect 15711 4867 15763 4915
rect 16402 4931 16454 4979
rect 16402 4897 16410 4931
rect 16444 4897 16454 4931
rect 16402 4849 16454 4897
rect 16484 4971 16553 4979
rect 16484 4937 16509 4971
rect 16543 4937 16553 4971
rect 16484 4895 16553 4937
rect 16583 4895 16649 4979
rect 16679 4895 16721 4979
rect 16751 4959 16817 4979
rect 16751 4925 16761 4959
rect 16795 4925 16817 4959
rect 16751 4895 16817 4925
rect 16847 4954 16906 4979
rect 16847 4920 16862 4954
rect 16896 4920 16906 4954
rect 16847 4895 16906 4920
rect 16936 4971 16990 4979
rect 16936 4937 16946 4971
rect 16980 4937 16990 4971
rect 16936 4895 16990 4937
rect 17020 4954 17074 4979
rect 17020 4920 17030 4954
rect 17064 4920 17074 4954
rect 17020 4895 17074 4920
rect 17104 4962 17156 4979
rect 17104 4928 17114 4962
rect 17148 4928 17156 4962
rect 17104 4895 17156 4928
rect 17210 4954 17262 4979
rect 17210 4920 17218 4954
rect 17252 4920 17262 4954
rect 17210 4895 17262 4920
rect 17292 4971 17346 4979
rect 17292 4937 17302 4971
rect 17336 4937 17346 4971
rect 17292 4895 17346 4937
rect 17376 4954 17430 4979
rect 17376 4920 17386 4954
rect 17420 4920 17430 4954
rect 17376 4895 17430 4920
rect 17460 4954 17514 4979
rect 17460 4920 17470 4954
rect 17504 4920 17514 4954
rect 17460 4895 17514 4920
rect 17544 4895 17604 4979
rect 17634 4967 17703 4979
rect 17634 4933 17659 4967
rect 17693 4933 17703 4967
rect 17634 4895 17703 4933
rect 16484 4849 16536 4895
rect 17651 4849 17703 4895
rect 17733 4931 17785 4979
rect 17733 4897 17743 4931
rect 17777 4897 17785 4931
rect 17733 4849 17785 4897
rect 6156 3277 6208 3293
rect 6156 3243 6164 3277
rect 6198 3243 6208 3277
rect 6156 3209 6208 3243
rect 6156 3175 6164 3209
rect 6198 3175 6208 3209
rect 6156 3163 6208 3175
rect 6238 3277 6290 3293
rect 6238 3243 6248 3277
rect 6282 3243 6290 3277
rect 6238 3209 6290 3243
rect 6238 3175 6248 3209
rect 6282 3175 6290 3209
rect 6238 3163 6290 3175
rect 1868 2193 1920 2241
rect 1868 2159 1876 2193
rect 1910 2159 1920 2193
rect 1868 2111 1920 2159
rect 1950 2233 2019 2241
rect 1950 2199 1975 2233
rect 2009 2199 2019 2233
rect 1950 2157 2019 2199
rect 2049 2157 2115 2241
rect 2145 2157 2187 2241
rect 2217 2221 2283 2241
rect 2217 2187 2227 2221
rect 2261 2187 2283 2221
rect 2217 2157 2283 2187
rect 2313 2216 2372 2241
rect 2313 2182 2328 2216
rect 2362 2182 2372 2216
rect 2313 2157 2372 2182
rect 2402 2233 2456 2241
rect 2402 2199 2412 2233
rect 2446 2199 2456 2233
rect 2402 2157 2456 2199
rect 2486 2216 2540 2241
rect 2486 2182 2496 2216
rect 2530 2182 2540 2216
rect 2486 2157 2540 2182
rect 2570 2224 2622 2241
rect 2570 2190 2580 2224
rect 2614 2190 2622 2224
rect 2570 2157 2622 2190
rect 2676 2216 2728 2241
rect 2676 2182 2684 2216
rect 2718 2182 2728 2216
rect 2676 2157 2728 2182
rect 2758 2233 2812 2241
rect 2758 2199 2768 2233
rect 2802 2199 2812 2233
rect 2758 2157 2812 2199
rect 2842 2216 2896 2241
rect 2842 2182 2852 2216
rect 2886 2182 2896 2216
rect 2842 2157 2896 2182
rect 2926 2216 2980 2241
rect 2926 2182 2936 2216
rect 2970 2182 2980 2216
rect 2926 2157 2980 2182
rect 3010 2157 3070 2241
rect 3100 2229 3169 2241
rect 3100 2195 3125 2229
rect 3159 2195 3169 2229
rect 3100 2157 3169 2195
rect 1950 2111 2002 2157
rect 3117 2111 3169 2157
rect 3199 2193 3251 2241
rect 3199 2159 3209 2193
rect 3243 2159 3251 2193
rect 3199 2111 3251 2159
rect 3938 2189 3990 2237
rect 3938 2155 3946 2189
rect 3980 2155 3990 2189
rect 3938 2107 3990 2155
rect 4020 2229 4089 2237
rect 4020 2195 4045 2229
rect 4079 2195 4089 2229
rect 4020 2153 4089 2195
rect 4119 2153 4185 2237
rect 4215 2153 4257 2237
rect 4287 2217 4353 2237
rect 4287 2183 4297 2217
rect 4331 2183 4353 2217
rect 4287 2153 4353 2183
rect 4383 2212 4442 2237
rect 4383 2178 4398 2212
rect 4432 2178 4442 2212
rect 4383 2153 4442 2178
rect 4472 2229 4526 2237
rect 4472 2195 4482 2229
rect 4516 2195 4526 2229
rect 4472 2153 4526 2195
rect 4556 2212 4610 2237
rect 4556 2178 4566 2212
rect 4600 2178 4610 2212
rect 4556 2153 4610 2178
rect 4640 2220 4692 2237
rect 4640 2186 4650 2220
rect 4684 2186 4692 2220
rect 4640 2153 4692 2186
rect 4746 2212 4798 2237
rect 4746 2178 4754 2212
rect 4788 2178 4798 2212
rect 4746 2153 4798 2178
rect 4828 2229 4882 2237
rect 4828 2195 4838 2229
rect 4872 2195 4882 2229
rect 4828 2153 4882 2195
rect 4912 2212 4966 2237
rect 4912 2178 4922 2212
rect 4956 2178 4966 2212
rect 4912 2153 4966 2178
rect 4996 2212 5050 2237
rect 4996 2178 5006 2212
rect 5040 2178 5050 2212
rect 4996 2153 5050 2178
rect 5080 2153 5140 2237
rect 5170 2225 5239 2237
rect 5170 2191 5195 2225
rect 5229 2191 5239 2225
rect 5170 2153 5239 2191
rect 4020 2107 4072 2153
rect 5187 2107 5239 2153
rect 5269 2189 5321 2237
rect 5269 2155 5279 2189
rect 5313 2155 5321 2189
rect 5269 2107 5321 2155
rect 5890 2189 5942 2237
rect 5890 2155 5898 2189
rect 5932 2155 5942 2189
rect 5890 2107 5942 2155
rect 5972 2229 6041 2237
rect 5972 2195 5997 2229
rect 6031 2195 6041 2229
rect 5972 2153 6041 2195
rect 6071 2153 6137 2237
rect 6167 2153 6209 2237
rect 6239 2217 6305 2237
rect 6239 2183 6249 2217
rect 6283 2183 6305 2217
rect 6239 2153 6305 2183
rect 6335 2212 6394 2237
rect 6335 2178 6350 2212
rect 6384 2178 6394 2212
rect 6335 2153 6394 2178
rect 6424 2229 6478 2237
rect 6424 2195 6434 2229
rect 6468 2195 6478 2229
rect 6424 2153 6478 2195
rect 6508 2212 6562 2237
rect 6508 2178 6518 2212
rect 6552 2178 6562 2212
rect 6508 2153 6562 2178
rect 6592 2220 6644 2237
rect 6592 2186 6602 2220
rect 6636 2186 6644 2220
rect 6592 2153 6644 2186
rect 6698 2212 6750 2237
rect 6698 2178 6706 2212
rect 6740 2178 6750 2212
rect 6698 2153 6750 2178
rect 6780 2229 6834 2237
rect 6780 2195 6790 2229
rect 6824 2195 6834 2229
rect 6780 2153 6834 2195
rect 6864 2212 6918 2237
rect 6864 2178 6874 2212
rect 6908 2178 6918 2212
rect 6864 2153 6918 2178
rect 6948 2212 7002 2237
rect 6948 2178 6958 2212
rect 6992 2178 7002 2212
rect 6948 2153 7002 2178
rect 7032 2153 7092 2237
rect 7122 2225 7191 2237
rect 7122 2191 7147 2225
rect 7181 2191 7191 2225
rect 7122 2153 7191 2191
rect 5972 2107 6024 2153
rect 7139 2107 7191 2153
rect 7221 2189 7273 2237
rect 7221 2155 7231 2189
rect 7265 2155 7273 2189
rect 7221 2107 7273 2155
rect 7892 2195 7944 2243
rect 7892 2161 7900 2195
rect 7934 2161 7944 2195
rect 7892 2113 7944 2161
rect 7974 2235 8043 2243
rect 7974 2201 7999 2235
rect 8033 2201 8043 2235
rect 7974 2159 8043 2201
rect 8073 2159 8139 2243
rect 8169 2159 8211 2243
rect 8241 2223 8307 2243
rect 8241 2189 8251 2223
rect 8285 2189 8307 2223
rect 8241 2159 8307 2189
rect 8337 2218 8396 2243
rect 8337 2184 8352 2218
rect 8386 2184 8396 2218
rect 8337 2159 8396 2184
rect 8426 2235 8480 2243
rect 8426 2201 8436 2235
rect 8470 2201 8480 2235
rect 8426 2159 8480 2201
rect 8510 2218 8564 2243
rect 8510 2184 8520 2218
rect 8554 2184 8564 2218
rect 8510 2159 8564 2184
rect 8594 2226 8646 2243
rect 8594 2192 8604 2226
rect 8638 2192 8646 2226
rect 8594 2159 8646 2192
rect 8700 2218 8752 2243
rect 8700 2184 8708 2218
rect 8742 2184 8752 2218
rect 8700 2159 8752 2184
rect 8782 2235 8836 2243
rect 8782 2201 8792 2235
rect 8826 2201 8836 2235
rect 8782 2159 8836 2201
rect 8866 2218 8920 2243
rect 8866 2184 8876 2218
rect 8910 2184 8920 2218
rect 8866 2159 8920 2184
rect 8950 2218 9004 2243
rect 8950 2184 8960 2218
rect 8994 2184 9004 2218
rect 8950 2159 9004 2184
rect 9034 2159 9094 2243
rect 9124 2231 9193 2243
rect 9124 2197 9149 2231
rect 9183 2197 9193 2231
rect 9124 2159 9193 2197
rect 7974 2113 8026 2159
rect 9141 2113 9193 2159
rect 9223 2195 9275 2243
rect 9223 2161 9233 2195
rect 9267 2161 9275 2195
rect 9223 2113 9275 2161
rect 9844 2195 9896 2243
rect 9844 2161 9852 2195
rect 9886 2161 9896 2195
rect 9844 2113 9896 2161
rect 9926 2235 9995 2243
rect 9926 2201 9951 2235
rect 9985 2201 9995 2235
rect 9926 2159 9995 2201
rect 10025 2159 10091 2243
rect 10121 2159 10163 2243
rect 10193 2223 10259 2243
rect 10193 2189 10203 2223
rect 10237 2189 10259 2223
rect 10193 2159 10259 2189
rect 10289 2218 10348 2243
rect 10289 2184 10304 2218
rect 10338 2184 10348 2218
rect 10289 2159 10348 2184
rect 10378 2235 10432 2243
rect 10378 2201 10388 2235
rect 10422 2201 10432 2235
rect 10378 2159 10432 2201
rect 10462 2218 10516 2243
rect 10462 2184 10472 2218
rect 10506 2184 10516 2218
rect 10462 2159 10516 2184
rect 10546 2226 10598 2243
rect 10546 2192 10556 2226
rect 10590 2192 10598 2226
rect 10546 2159 10598 2192
rect 10652 2218 10704 2243
rect 10652 2184 10660 2218
rect 10694 2184 10704 2218
rect 10652 2159 10704 2184
rect 10734 2235 10788 2243
rect 10734 2201 10744 2235
rect 10778 2201 10788 2235
rect 10734 2159 10788 2201
rect 10818 2218 10872 2243
rect 10818 2184 10828 2218
rect 10862 2184 10872 2218
rect 10818 2159 10872 2184
rect 10902 2218 10956 2243
rect 10902 2184 10912 2218
rect 10946 2184 10956 2218
rect 10902 2159 10956 2184
rect 10986 2159 11046 2243
rect 11076 2231 11145 2243
rect 11076 2197 11101 2231
rect 11135 2197 11145 2231
rect 11076 2159 11145 2197
rect 9926 2113 9978 2159
rect 11093 2113 11145 2159
rect 11175 2195 11227 2243
rect 11175 2161 11185 2195
rect 11219 2161 11227 2195
rect 11175 2113 11227 2161
rect 11836 2195 11888 2243
rect 11836 2161 11844 2195
rect 11878 2161 11888 2195
rect 11836 2113 11888 2161
rect 11918 2235 11987 2243
rect 11918 2201 11943 2235
rect 11977 2201 11987 2235
rect 11918 2159 11987 2201
rect 12017 2159 12083 2243
rect 12113 2159 12155 2243
rect 12185 2223 12251 2243
rect 12185 2189 12195 2223
rect 12229 2189 12251 2223
rect 12185 2159 12251 2189
rect 12281 2218 12340 2243
rect 12281 2184 12296 2218
rect 12330 2184 12340 2218
rect 12281 2159 12340 2184
rect 12370 2235 12424 2243
rect 12370 2201 12380 2235
rect 12414 2201 12424 2235
rect 12370 2159 12424 2201
rect 12454 2218 12508 2243
rect 12454 2184 12464 2218
rect 12498 2184 12508 2218
rect 12454 2159 12508 2184
rect 12538 2226 12590 2243
rect 12538 2192 12548 2226
rect 12582 2192 12590 2226
rect 12538 2159 12590 2192
rect 12644 2218 12696 2243
rect 12644 2184 12652 2218
rect 12686 2184 12696 2218
rect 12644 2159 12696 2184
rect 12726 2235 12780 2243
rect 12726 2201 12736 2235
rect 12770 2201 12780 2235
rect 12726 2159 12780 2201
rect 12810 2218 12864 2243
rect 12810 2184 12820 2218
rect 12854 2184 12864 2218
rect 12810 2159 12864 2184
rect 12894 2218 12948 2243
rect 12894 2184 12904 2218
rect 12938 2184 12948 2218
rect 12894 2159 12948 2184
rect 12978 2159 13038 2243
rect 13068 2231 13137 2243
rect 13068 2197 13093 2231
rect 13127 2197 13137 2231
rect 13068 2159 13137 2197
rect 11918 2113 11970 2159
rect 13085 2113 13137 2159
rect 13167 2195 13219 2243
rect 13167 2161 13177 2195
rect 13211 2161 13219 2195
rect 13167 2113 13219 2161
rect 13788 2195 13840 2243
rect 13788 2161 13796 2195
rect 13830 2161 13840 2195
rect 13788 2113 13840 2161
rect 13870 2235 13939 2243
rect 13870 2201 13895 2235
rect 13929 2201 13939 2235
rect 13870 2159 13939 2201
rect 13969 2159 14035 2243
rect 14065 2159 14107 2243
rect 14137 2223 14203 2243
rect 14137 2189 14147 2223
rect 14181 2189 14203 2223
rect 14137 2159 14203 2189
rect 14233 2218 14292 2243
rect 14233 2184 14248 2218
rect 14282 2184 14292 2218
rect 14233 2159 14292 2184
rect 14322 2235 14376 2243
rect 14322 2201 14332 2235
rect 14366 2201 14376 2235
rect 14322 2159 14376 2201
rect 14406 2218 14460 2243
rect 14406 2184 14416 2218
rect 14450 2184 14460 2218
rect 14406 2159 14460 2184
rect 14490 2226 14542 2243
rect 14490 2192 14500 2226
rect 14534 2192 14542 2226
rect 14490 2159 14542 2192
rect 14596 2218 14648 2243
rect 14596 2184 14604 2218
rect 14638 2184 14648 2218
rect 14596 2159 14648 2184
rect 14678 2235 14732 2243
rect 14678 2201 14688 2235
rect 14722 2201 14732 2235
rect 14678 2159 14732 2201
rect 14762 2218 14816 2243
rect 14762 2184 14772 2218
rect 14806 2184 14816 2218
rect 14762 2159 14816 2184
rect 14846 2218 14900 2243
rect 14846 2184 14856 2218
rect 14890 2184 14900 2218
rect 14846 2159 14900 2184
rect 14930 2159 14990 2243
rect 15020 2231 15089 2243
rect 15020 2197 15045 2231
rect 15079 2197 15089 2231
rect 15020 2159 15089 2197
rect 13870 2113 13922 2159
rect 15037 2113 15089 2159
rect 15119 2195 15171 2243
rect 15119 2161 15129 2195
rect 15163 2161 15171 2195
rect 15119 2113 15171 2161
rect 15852 2195 15904 2243
rect 15852 2161 15860 2195
rect 15894 2161 15904 2195
rect 15852 2113 15904 2161
rect 15934 2235 16003 2243
rect 15934 2201 15959 2235
rect 15993 2201 16003 2235
rect 15934 2159 16003 2201
rect 16033 2159 16099 2243
rect 16129 2159 16171 2243
rect 16201 2223 16267 2243
rect 16201 2189 16211 2223
rect 16245 2189 16267 2223
rect 16201 2159 16267 2189
rect 16297 2218 16356 2243
rect 16297 2184 16312 2218
rect 16346 2184 16356 2218
rect 16297 2159 16356 2184
rect 16386 2235 16440 2243
rect 16386 2201 16396 2235
rect 16430 2201 16440 2235
rect 16386 2159 16440 2201
rect 16470 2218 16524 2243
rect 16470 2184 16480 2218
rect 16514 2184 16524 2218
rect 16470 2159 16524 2184
rect 16554 2226 16606 2243
rect 16554 2192 16564 2226
rect 16598 2192 16606 2226
rect 16554 2159 16606 2192
rect 16660 2218 16712 2243
rect 16660 2184 16668 2218
rect 16702 2184 16712 2218
rect 16660 2159 16712 2184
rect 16742 2235 16796 2243
rect 16742 2201 16752 2235
rect 16786 2201 16796 2235
rect 16742 2159 16796 2201
rect 16826 2218 16880 2243
rect 16826 2184 16836 2218
rect 16870 2184 16880 2218
rect 16826 2159 16880 2184
rect 16910 2218 16964 2243
rect 16910 2184 16920 2218
rect 16954 2184 16964 2218
rect 16910 2159 16964 2184
rect 16994 2159 17054 2243
rect 17084 2231 17153 2243
rect 17084 2197 17109 2231
rect 17143 2197 17153 2231
rect 17084 2159 17153 2197
rect 15934 2113 15986 2159
rect 17101 2113 17153 2159
rect 17183 2195 17235 2243
rect 17183 2161 17193 2195
rect 17227 2161 17235 2195
rect 17183 2113 17235 2161
<< pdiff >>
rect 18643 43374 18843 43382
rect 18643 43340 18655 43374
rect 18689 43340 18723 43374
rect 18757 43340 18843 43374
rect 18643 43330 18843 43340
rect 18643 43290 18843 43300
rect 18643 43256 18655 43290
rect 18689 43256 18723 43290
rect 18757 43256 18793 43290
rect 18827 43256 18843 43290
rect 18643 43246 18843 43256
rect 18643 43206 18843 43216
rect 18643 43172 18655 43206
rect 18689 43172 18723 43206
rect 18757 43172 18843 43206
rect 18643 43162 18843 43172
rect 18643 43122 18843 43132
rect 18643 43088 18655 43122
rect 18689 43088 18723 43122
rect 18757 43088 18793 43122
rect 18827 43088 18843 43122
rect 18643 43078 18843 43088
rect 18643 43038 18843 43048
rect 18643 43004 18655 43038
rect 18689 43004 18723 43038
rect 18757 43004 18843 43038
rect 18643 42994 18843 43004
rect 18643 42954 18843 42964
rect 18643 42920 18655 42954
rect 18689 42920 18723 42954
rect 18757 42920 18793 42954
rect 18827 42920 18843 42954
rect 18643 42910 18843 42920
rect 18643 42870 18843 42880
rect 18643 42836 18655 42870
rect 18689 42836 18723 42870
rect 18757 42836 18843 42870
rect 18643 42826 18843 42836
rect 18643 42786 18843 42796
rect 18643 42752 18655 42786
rect 18689 42752 18723 42786
rect 18757 42752 18793 42786
rect 18827 42752 18843 42786
rect 18643 42742 18843 42752
rect 18643 42702 18843 42712
rect 18643 42668 18655 42702
rect 18689 42668 18723 42702
rect 18757 42668 18843 42702
rect 18643 42658 18843 42668
rect 18643 42618 18843 42628
rect 18643 42584 18655 42618
rect 18689 42584 18723 42618
rect 18757 42584 18793 42618
rect 18827 42584 18843 42618
rect 18643 42574 18843 42584
rect 18643 42534 18843 42544
rect 18643 42500 18655 42534
rect 18689 42500 18723 42534
rect 18757 42500 18843 42534
rect 18643 42490 18843 42500
rect 18643 42450 18843 42460
rect 18643 42416 18655 42450
rect 18689 42416 18723 42450
rect 18757 42416 18793 42450
rect 18827 42416 18843 42450
rect 18643 42406 18843 42416
rect 18643 42366 18843 42376
rect 18643 42332 18655 42366
rect 18689 42332 18723 42366
rect 18757 42332 18843 42366
rect 18643 42322 18843 42332
rect 18643 42282 18843 42292
rect 18643 42248 18655 42282
rect 18689 42248 18723 42282
rect 18757 42248 18793 42282
rect 18827 42248 18843 42282
rect 18643 42238 18843 42248
rect 18643 42198 18843 42208
rect 18643 42164 18655 42198
rect 18689 42164 18723 42198
rect 18757 42164 18843 42198
rect 18643 42154 18843 42164
rect 18643 42114 18843 42124
rect 18643 42080 18655 42114
rect 18689 42080 18723 42114
rect 18757 42080 18793 42114
rect 18827 42080 18843 42114
rect 18643 42070 18843 42080
rect 18643 42030 18843 42040
rect 18643 41996 18655 42030
rect 18689 41996 18723 42030
rect 18757 41996 18793 42030
rect 18827 41996 18843 42030
rect 18643 41988 18843 41996
rect 18627 41397 18827 41405
rect 18627 41363 18639 41397
rect 18673 41363 18707 41397
rect 18741 41363 18827 41397
rect 18627 41302 18827 41363
rect 18627 41262 18827 41272
rect 18627 41228 18639 41262
rect 18673 41228 18707 41262
rect 18741 41228 18775 41262
rect 18809 41228 18827 41262
rect 18627 41218 18827 41228
rect 18627 41178 18827 41188
rect 18627 41144 18639 41178
rect 18673 41144 18707 41178
rect 18741 41144 18827 41178
rect 18627 41134 18827 41144
rect 18627 41094 18827 41104
rect 18627 41060 18639 41094
rect 18673 41060 18707 41094
rect 18741 41060 18775 41094
rect 18809 41060 18827 41094
rect 18627 41050 18827 41060
rect 18627 41010 18827 41020
rect 18627 40976 18639 41010
rect 18673 40976 18707 41010
rect 18741 40976 18827 41010
rect 18627 40966 18827 40976
rect 18627 40926 18827 40936
rect 18627 40892 18639 40926
rect 18673 40892 18707 40926
rect 18741 40892 18775 40926
rect 18809 40892 18827 40926
rect 18627 40882 18827 40892
rect 18627 40842 18827 40852
rect 18627 40808 18639 40842
rect 18673 40808 18707 40842
rect 18741 40808 18827 40842
rect 18627 40798 18827 40808
rect 18627 40758 18827 40768
rect 18627 40724 18639 40758
rect 18673 40724 18707 40758
rect 18741 40724 18775 40758
rect 18809 40724 18827 40758
rect 18627 40714 18827 40724
rect 18627 40674 18827 40684
rect 18627 40640 18639 40674
rect 18673 40640 18707 40674
rect 18741 40640 18827 40674
rect 18627 40630 18827 40640
rect 18627 40590 18827 40600
rect 18627 40556 18639 40590
rect 18673 40556 18707 40590
rect 18741 40556 18775 40590
rect 18809 40556 18827 40590
rect 18627 40546 18827 40556
rect 18627 40506 18827 40516
rect 18627 40472 18639 40506
rect 18673 40472 18707 40506
rect 18741 40472 18827 40506
rect 18627 40462 18827 40472
rect 18627 40422 18827 40432
rect 18627 40388 18639 40422
rect 18673 40388 18707 40422
rect 18741 40388 18775 40422
rect 18809 40388 18827 40422
rect 18627 40378 18827 40388
rect 18627 40338 18827 40348
rect 18627 40304 18639 40338
rect 18673 40304 18707 40338
rect 18741 40304 18827 40338
rect 18627 40296 18827 40304
rect 18635 39582 18835 39590
rect 18635 39548 18647 39582
rect 18681 39548 18715 39582
rect 18749 39548 18835 39582
rect 18635 39538 18835 39548
rect 18635 39498 18835 39508
rect 18635 39464 18647 39498
rect 18681 39464 18715 39498
rect 18749 39464 18783 39498
rect 18817 39464 18835 39498
rect 18635 39454 18835 39464
rect 18635 39414 18835 39424
rect 18635 39380 18647 39414
rect 18681 39380 18715 39414
rect 18749 39380 18835 39414
rect 18635 39370 18835 39380
rect 18635 39330 18835 39340
rect 18635 39296 18647 39330
rect 18681 39296 18715 39330
rect 18749 39296 18783 39330
rect 18817 39296 18835 39330
rect 18635 39286 18835 39296
rect 18635 39246 18835 39256
rect 18635 39212 18647 39246
rect 18681 39212 18715 39246
rect 18749 39212 18835 39246
rect 18635 39202 18835 39212
rect 18635 39162 18835 39172
rect 18635 39128 18647 39162
rect 18681 39128 18715 39162
rect 18749 39128 18783 39162
rect 18817 39128 18835 39162
rect 18635 39118 18835 39128
rect 18635 39078 18835 39088
rect 18635 39044 18647 39078
rect 18681 39044 18715 39078
rect 18749 39044 18835 39078
rect 18635 39034 18835 39044
rect 18635 38994 18835 39004
rect 18635 38960 18647 38994
rect 18681 38960 18715 38994
rect 18749 38960 18783 38994
rect 18817 38960 18835 38994
rect 18635 38950 18835 38960
rect 18635 38910 18835 38920
rect 18635 38876 18647 38910
rect 18681 38876 18715 38910
rect 18749 38876 18835 38910
rect 18635 38868 18835 38876
rect 18649 38337 18849 38347
rect 18649 38303 18661 38337
rect 18695 38303 18849 38337
rect 18649 38293 18849 38303
rect 18649 38253 18849 38263
rect 18649 38219 18661 38253
rect 18695 38219 18729 38253
rect 18763 38219 18797 38253
rect 18831 38219 18849 38253
rect 18649 38209 18849 38219
rect 18649 38169 18849 38179
rect 18649 38135 18661 38169
rect 18695 38135 18729 38169
rect 18763 38135 18849 38169
rect 18649 38125 18849 38135
rect 18649 38085 18849 38095
rect 18649 38051 18661 38085
rect 18695 38051 18729 38085
rect 18763 38051 18797 38085
rect 18831 38051 18849 38085
rect 18649 38041 18849 38051
rect 18649 38001 18849 38011
rect 18649 37967 18661 38001
rect 18695 37967 18729 38001
rect 18763 37967 18849 38001
rect 18649 37957 18849 37967
rect 18649 37917 18849 37927
rect 18649 37883 18661 37917
rect 18695 37883 18729 37917
rect 18763 37883 18797 37917
rect 18831 37883 18849 37917
rect 18649 37873 18849 37883
rect 18649 37799 18849 37843
rect 18649 37765 18661 37799
rect 18695 37765 18729 37799
rect 18763 37765 18797 37799
rect 18831 37765 18849 37799
rect 18649 37757 18849 37765
rect 18661 37179 18861 37187
rect 18661 37145 18673 37179
rect 18707 37145 18861 37179
rect 18661 37135 18861 37145
rect 18661 37095 18861 37105
rect 18661 37061 18673 37095
rect 18707 37061 18741 37095
rect 18775 37061 18809 37095
rect 18843 37061 18861 37095
rect 18661 37051 18861 37061
rect 18661 37011 18861 37021
rect 18661 36977 18673 37011
rect 18707 36977 18741 37011
rect 18775 36977 18861 37011
rect 18661 36967 18861 36977
rect 18661 36927 18861 36937
rect 18661 36893 18673 36927
rect 18707 36893 18741 36927
rect 18775 36893 18809 36927
rect 18843 36893 18861 36927
rect 18661 36883 18861 36893
rect 18661 36843 18861 36853
rect 18661 36809 18673 36843
rect 18707 36809 18741 36843
rect 18775 36809 18809 36843
rect 18843 36809 18861 36843
rect 18661 36801 18861 36809
rect 18669 36299 18869 36307
rect 18669 36265 18681 36299
rect 18715 36265 18749 36299
rect 18783 36265 18817 36299
rect 18851 36265 18869 36299
rect 18669 36255 18869 36265
rect 18669 36215 18869 36225
rect 18669 36181 18681 36215
rect 18715 36181 18749 36215
rect 18783 36181 18817 36215
rect 18851 36181 18869 36215
rect 18669 36171 18869 36181
rect 18669 36131 18869 36141
rect 18669 36097 18681 36131
rect 18715 36097 18749 36131
rect 18783 36097 18817 36131
rect 18851 36097 18869 36131
rect 18669 36089 18869 36097
rect 18693 34913 18893 34921
rect 18693 34879 18705 34913
rect 18739 34879 18776 34913
rect 18810 34879 18847 34913
rect 18881 34879 18893 34913
rect 18693 34869 18893 34879
rect 18693 34829 18893 34839
rect 18693 34795 18705 34829
rect 18739 34795 18773 34829
rect 18807 34795 18841 34829
rect 18875 34795 18893 34829
rect 18693 34787 18893 34795
rect 18693 34772 18821 34787
rect 18693 34732 18821 34742
rect 18693 34698 18705 34732
rect 18739 34698 18773 34732
rect 18807 34698 18821 34732
rect 18693 34690 18821 34698
rect 18693 34628 18893 34636
rect 18693 34594 18711 34628
rect 18745 34594 18779 34628
rect 18813 34594 18847 34628
rect 18881 34594 18893 34628
rect 18693 34584 18893 34594
rect 18693 34544 18893 34554
rect 18693 34510 18735 34544
rect 18769 34510 18815 34544
rect 18849 34510 18893 34544
rect 18693 34500 18893 34510
rect 18693 34458 18893 34470
rect 18693 34424 18705 34458
rect 18739 34424 18776 34458
rect 18810 34424 18847 34458
rect 18881 34424 18893 34458
rect 18693 34416 18893 34424
rect 18693 34334 18777 34342
rect 18693 34300 18713 34334
rect 18747 34300 18777 34334
rect 18693 34289 18777 34300
rect 18693 34175 18777 34259
rect 18693 34135 18777 34145
rect 18693 34101 18723 34135
rect 18757 34101 18777 34135
rect 18693 34091 18777 34101
rect 18693 34046 18777 34061
rect 18693 34040 18843 34046
rect 18693 34006 18713 34040
rect 18747 34006 18843 34040
rect 18693 33996 18843 34006
rect 18693 33956 18843 33966
rect 18693 33922 18705 33956
rect 18739 33922 18773 33956
rect 18807 33922 18843 33956
rect 18693 33879 18843 33922
rect 18693 33864 18777 33879
rect 18693 33761 18777 33834
rect 18693 33717 18777 33731
rect 18693 33683 18718 33717
rect 18752 33683 18777 33717
rect 18693 33666 18777 33683
rect 18693 33625 18777 33636
rect 18693 33591 18713 33625
rect 18747 33591 18777 33625
rect 18693 33581 18777 33591
rect 18693 33541 18777 33551
rect 18693 33507 18705 33541
rect 18739 33507 18777 33541
rect 18693 33499 18777 33507
rect 18699 33437 18827 33445
rect 18699 33403 18713 33437
rect 18747 33403 18781 33437
rect 18815 33403 18827 33437
rect 18699 33393 18827 33403
rect 18699 33353 18827 33363
rect 18699 33319 18729 33353
rect 18763 33319 18827 33353
rect 18699 33309 18827 33319
rect 18699 33269 18827 33279
rect 18699 33235 18713 33269
rect 18747 33235 18781 33269
rect 18815 33235 18827 33269
rect 18699 33227 18827 33235
rect 18693 32631 18893 32639
rect 18693 32597 18705 32631
rect 18739 32597 18776 32631
rect 18810 32597 18847 32631
rect 18881 32597 18893 32631
rect 18693 32587 18893 32597
rect 18693 32547 18893 32557
rect 18693 32513 18705 32547
rect 18739 32513 18773 32547
rect 18807 32513 18841 32547
rect 18875 32513 18893 32547
rect 18693 32505 18893 32513
rect 18693 32490 18821 32505
rect 18693 32450 18821 32460
rect 18693 32416 18705 32450
rect 18739 32416 18773 32450
rect 18807 32416 18821 32450
rect 18693 32408 18821 32416
rect 18693 32346 18893 32354
rect 18693 32312 18711 32346
rect 18745 32312 18779 32346
rect 18813 32312 18847 32346
rect 18881 32312 18893 32346
rect 18693 32302 18893 32312
rect 18693 32262 18893 32272
rect 18693 32228 18735 32262
rect 18769 32228 18815 32262
rect 18849 32228 18893 32262
rect 18693 32218 18893 32228
rect 18693 32176 18893 32188
rect 18693 32142 18705 32176
rect 18739 32142 18776 32176
rect 18810 32142 18847 32176
rect 18881 32142 18893 32176
rect 18693 32134 18893 32142
rect 18693 32052 18777 32060
rect 18693 32018 18713 32052
rect 18747 32018 18777 32052
rect 18693 32007 18777 32018
rect 18693 31893 18777 31977
rect 18693 31853 18777 31863
rect 18693 31819 18723 31853
rect 18757 31819 18777 31853
rect 18693 31809 18777 31819
rect 18693 31764 18777 31779
rect 18693 31758 18843 31764
rect 18693 31724 18713 31758
rect 18747 31724 18843 31758
rect 18693 31714 18843 31724
rect 18693 31674 18843 31684
rect 18693 31640 18705 31674
rect 18739 31640 18773 31674
rect 18807 31640 18843 31674
rect 18693 31597 18843 31640
rect 18693 31582 18777 31597
rect 18693 31479 18777 31552
rect 18693 31435 18777 31449
rect 18693 31401 18718 31435
rect 18752 31401 18777 31435
rect 18693 31384 18777 31401
rect 18693 31343 18777 31354
rect 18693 31309 18713 31343
rect 18747 31309 18777 31343
rect 18693 31299 18777 31309
rect 18693 31259 18777 31269
rect 18693 31225 18705 31259
rect 18739 31225 18777 31259
rect 18693 31217 18777 31225
rect 18699 31155 18827 31163
rect 18699 31121 18713 31155
rect 18747 31121 18781 31155
rect 18815 31121 18827 31155
rect 18699 31111 18827 31121
rect 18699 31071 18827 31081
rect 18699 31037 18729 31071
rect 18763 31037 18827 31071
rect 18699 31027 18827 31037
rect 18699 30987 18827 30997
rect 18699 30953 18713 30987
rect 18747 30953 18781 30987
rect 18815 30953 18827 30987
rect 18699 30945 18827 30953
rect 18697 30385 18897 30393
rect 18697 30351 18709 30385
rect 18743 30351 18780 30385
rect 18814 30351 18851 30385
rect 18885 30351 18897 30385
rect 18697 30341 18897 30351
rect 18697 30301 18897 30311
rect 18697 30267 18709 30301
rect 18743 30267 18777 30301
rect 18811 30267 18845 30301
rect 18879 30267 18897 30301
rect 18697 30259 18897 30267
rect 18697 30244 18825 30259
rect 18697 30204 18825 30214
rect 18697 30170 18709 30204
rect 18743 30170 18777 30204
rect 18811 30170 18825 30204
rect 18697 30162 18825 30170
rect 18697 30100 18897 30108
rect 18697 30066 18715 30100
rect 18749 30066 18783 30100
rect 18817 30066 18851 30100
rect 18885 30066 18897 30100
rect 18697 30056 18897 30066
rect 18697 30016 18897 30026
rect 18697 29982 18739 30016
rect 18773 29982 18819 30016
rect 18853 29982 18897 30016
rect 18697 29972 18897 29982
rect 18697 29930 18897 29942
rect 18697 29896 18709 29930
rect 18743 29896 18780 29930
rect 18814 29896 18851 29930
rect 18885 29896 18897 29930
rect 18697 29888 18897 29896
rect 18697 29806 18781 29814
rect 18697 29772 18717 29806
rect 18751 29772 18781 29806
rect 18697 29761 18781 29772
rect 18697 29647 18781 29731
rect 18697 29607 18781 29617
rect 18697 29573 18727 29607
rect 18761 29573 18781 29607
rect 18697 29563 18781 29573
rect 18697 29518 18781 29533
rect 18697 29512 18847 29518
rect 18697 29478 18717 29512
rect 18751 29478 18847 29512
rect 18697 29468 18847 29478
rect 18697 29428 18847 29438
rect 18697 29394 18709 29428
rect 18743 29394 18777 29428
rect 18811 29394 18847 29428
rect 18697 29351 18847 29394
rect 18697 29336 18781 29351
rect 18697 29233 18781 29306
rect 18697 29189 18781 29203
rect 18697 29155 18722 29189
rect 18756 29155 18781 29189
rect 18697 29138 18781 29155
rect 18697 29097 18781 29108
rect 18697 29063 18717 29097
rect 18751 29063 18781 29097
rect 18697 29053 18781 29063
rect 18697 29013 18781 29023
rect 18697 28979 18709 29013
rect 18743 28979 18781 29013
rect 18697 28971 18781 28979
rect 18703 28909 18831 28917
rect 18703 28875 18717 28909
rect 18751 28875 18785 28909
rect 18819 28875 18831 28909
rect 18703 28865 18831 28875
rect 18703 28825 18831 28835
rect 18703 28791 18733 28825
rect 18767 28791 18831 28825
rect 18703 28781 18831 28791
rect 18703 28741 18831 28751
rect 18703 28707 18717 28741
rect 18751 28707 18785 28741
rect 18819 28707 18831 28741
rect 18703 28699 18831 28707
rect 18689 28199 18889 28207
rect 18689 28165 18701 28199
rect 18735 28165 18772 28199
rect 18806 28165 18843 28199
rect 18877 28165 18889 28199
rect 18689 28155 18889 28165
rect 18689 28115 18889 28125
rect 18689 28081 18701 28115
rect 18735 28081 18769 28115
rect 18803 28081 18837 28115
rect 18871 28081 18889 28115
rect 18689 28073 18889 28081
rect 18689 28058 18817 28073
rect 18689 28018 18817 28028
rect 18689 27984 18701 28018
rect 18735 27984 18769 28018
rect 18803 27984 18817 28018
rect 18689 27976 18817 27984
rect 18689 27914 18889 27922
rect 18689 27880 18707 27914
rect 18741 27880 18775 27914
rect 18809 27880 18843 27914
rect 18877 27880 18889 27914
rect 18689 27870 18889 27880
rect 18689 27830 18889 27840
rect 18689 27796 18731 27830
rect 18765 27796 18811 27830
rect 18845 27796 18889 27830
rect 18689 27786 18889 27796
rect 18689 27744 18889 27756
rect 18689 27710 18701 27744
rect 18735 27710 18772 27744
rect 18806 27710 18843 27744
rect 18877 27710 18889 27744
rect 18689 27702 18889 27710
rect 18689 27620 18773 27628
rect 18689 27586 18709 27620
rect 18743 27586 18773 27620
rect 18689 27575 18773 27586
rect 18689 27461 18773 27545
rect 18689 27421 18773 27431
rect 18689 27387 18719 27421
rect 18753 27387 18773 27421
rect 18689 27377 18773 27387
rect 18689 27332 18773 27347
rect 18689 27326 18839 27332
rect 18689 27292 18709 27326
rect 18743 27292 18839 27326
rect 18689 27282 18839 27292
rect 18689 27242 18839 27252
rect 18689 27208 18701 27242
rect 18735 27208 18769 27242
rect 18803 27208 18839 27242
rect 18689 27165 18839 27208
rect 18689 27150 18773 27165
rect 18689 27047 18773 27120
rect 18689 27003 18773 27017
rect 18689 26969 18714 27003
rect 18748 26969 18773 27003
rect 18689 26952 18773 26969
rect 18689 26911 18773 26922
rect 18689 26877 18709 26911
rect 18743 26877 18773 26911
rect 18689 26867 18773 26877
rect 18689 26827 18773 26837
rect 18689 26793 18701 26827
rect 18735 26793 18773 26827
rect 18689 26785 18773 26793
rect 18695 26723 18823 26731
rect 18695 26689 18709 26723
rect 18743 26689 18777 26723
rect 18811 26689 18823 26723
rect 18695 26679 18823 26689
rect 18695 26639 18823 26649
rect 18695 26605 18725 26639
rect 18759 26605 18823 26639
rect 18695 26595 18823 26605
rect 18695 26555 18823 26565
rect 18695 26521 18709 26555
rect 18743 26521 18777 26555
rect 18811 26521 18823 26555
rect 18695 26513 18823 26521
rect 18693 25953 18893 25961
rect 18693 25919 18705 25953
rect 18739 25919 18776 25953
rect 18810 25919 18847 25953
rect 18881 25919 18893 25953
rect 18693 25909 18893 25919
rect 18693 25869 18893 25879
rect 18693 25835 18705 25869
rect 18739 25835 18773 25869
rect 18807 25835 18841 25869
rect 18875 25835 18893 25869
rect 18693 25827 18893 25835
rect 18693 25812 18821 25827
rect 18693 25772 18821 25782
rect 18693 25738 18705 25772
rect 18739 25738 18773 25772
rect 18807 25738 18821 25772
rect 18693 25730 18821 25738
rect 18693 25668 18893 25676
rect 18693 25634 18711 25668
rect 18745 25634 18779 25668
rect 18813 25634 18847 25668
rect 18881 25634 18893 25668
rect 18693 25624 18893 25634
rect 18693 25584 18893 25594
rect 18693 25550 18735 25584
rect 18769 25550 18815 25584
rect 18849 25550 18893 25584
rect 18693 25540 18893 25550
rect 18693 25498 18893 25510
rect 18693 25464 18705 25498
rect 18739 25464 18776 25498
rect 18810 25464 18847 25498
rect 18881 25464 18893 25498
rect 18693 25456 18893 25464
rect 18693 25374 18777 25382
rect 18693 25340 18713 25374
rect 18747 25340 18777 25374
rect 18693 25329 18777 25340
rect 18693 25215 18777 25299
rect 18693 25175 18777 25185
rect 18693 25141 18723 25175
rect 18757 25141 18777 25175
rect 18693 25131 18777 25141
rect 18693 25086 18777 25101
rect 18693 25080 18843 25086
rect 18693 25046 18713 25080
rect 18747 25046 18843 25080
rect 18693 25036 18843 25046
rect 18693 24996 18843 25006
rect 18693 24962 18705 24996
rect 18739 24962 18773 24996
rect 18807 24962 18843 24996
rect 18693 24919 18843 24962
rect 18693 24904 18777 24919
rect 18693 24801 18777 24874
rect 18693 24757 18777 24771
rect 18693 24723 18718 24757
rect 18752 24723 18777 24757
rect 18693 24706 18777 24723
rect 18693 24665 18777 24676
rect 18693 24631 18713 24665
rect 18747 24631 18777 24665
rect 18693 24621 18777 24631
rect 18693 24581 18777 24591
rect 18693 24547 18705 24581
rect 18739 24547 18777 24581
rect 18693 24539 18777 24547
rect 18699 24477 18827 24485
rect 18699 24443 18713 24477
rect 18747 24443 18781 24477
rect 18815 24443 18827 24477
rect 18699 24433 18827 24443
rect 18699 24393 18827 24403
rect 18699 24359 18729 24393
rect 18763 24359 18827 24393
rect 18699 24349 18827 24359
rect 18699 24309 18827 24319
rect 18699 24275 18713 24309
rect 18747 24275 18781 24309
rect 18815 24275 18827 24309
rect 18699 24267 18827 24275
rect 7697 23305 7749 23319
rect 7697 23271 7705 23305
rect 7739 23271 7749 23305
rect 7697 23237 7749 23271
rect 7697 23203 7705 23237
rect 7739 23203 7749 23237
rect 7697 23191 7749 23203
rect 7779 23289 7833 23319
rect 7779 23255 7789 23289
rect 7823 23255 7833 23289
rect 7779 23191 7833 23255
rect 7863 23305 7915 23319
rect 7863 23271 7873 23305
rect 7907 23271 7915 23305
rect 7863 23237 7915 23271
rect 7969 23313 8021 23325
rect 7969 23279 7977 23313
rect 8011 23279 8021 23313
rect 7969 23241 8021 23279
rect 8051 23305 8106 23325
rect 8051 23271 8061 23305
rect 8095 23271 8106 23305
rect 8051 23241 8106 23271
rect 8136 23300 8201 23325
rect 8136 23266 8153 23300
rect 8187 23266 8201 23300
rect 8136 23241 8201 23266
rect 8231 23241 8304 23325
rect 8334 23313 8436 23325
rect 8334 23279 8392 23313
rect 8426 23279 8436 23313
rect 8334 23245 8436 23279
rect 8334 23241 8392 23245
rect 7863 23203 7873 23237
rect 7907 23203 7915 23237
rect 7863 23191 7915 23203
rect 8349 23211 8392 23241
rect 8426 23211 8436 23245
rect 8349 23175 8436 23211
rect 8466 23305 8531 23325
rect 8466 23271 8476 23305
rect 8510 23271 8531 23305
rect 8466 23241 8531 23271
rect 8561 23295 8615 23325
rect 8561 23261 8571 23295
rect 8605 23261 8615 23295
rect 8561 23241 8615 23261
rect 8645 23241 8729 23325
rect 8759 23305 8812 23325
rect 8759 23271 8770 23305
rect 8804 23271 8812 23305
rect 8759 23241 8812 23271
rect 8886 23313 8940 23325
rect 8886 23279 8894 23313
rect 8928 23279 8940 23313
rect 8886 23242 8940 23279
rect 8466 23175 8516 23241
rect 8886 23208 8894 23242
rect 8928 23208 8940 23242
rect 8886 23171 8940 23208
rect 8886 23137 8894 23171
rect 8928 23137 8940 23171
rect 8886 23125 8940 23137
rect 8970 23283 9024 23325
rect 8970 23249 8980 23283
rect 9014 23249 9024 23283
rect 8970 23203 9024 23249
rect 8970 23169 8980 23203
rect 9014 23169 9024 23203
rect 8970 23125 9024 23169
rect 9054 23307 9106 23325
rect 9054 23273 9064 23307
rect 9098 23273 9106 23307
rect 9054 23239 9106 23273
rect 9054 23205 9064 23239
rect 9098 23205 9106 23239
rect 9054 23171 9106 23205
rect 9160 23313 9212 23325
rect 9160 23279 9168 23313
rect 9202 23279 9212 23313
rect 9160 23245 9212 23279
rect 9160 23211 9168 23245
rect 9202 23211 9212 23245
rect 9160 23197 9212 23211
rect 9242 23313 9309 23325
rect 9242 23279 9265 23313
rect 9299 23279 9309 23313
rect 9242 23245 9309 23279
rect 9242 23211 9265 23245
rect 9299 23211 9309 23245
rect 9242 23197 9309 23211
rect 9054 23137 9064 23171
rect 9098 23137 9106 23171
rect 9054 23125 9106 23137
rect 9257 23177 9309 23197
rect 9257 23143 9265 23177
rect 9299 23143 9309 23177
rect 9257 23125 9309 23143
rect 9339 23313 9391 23325
rect 9339 23279 9349 23313
rect 9383 23279 9391 23313
rect 9943 23309 9995 23323
rect 9339 23242 9391 23279
rect 9339 23208 9349 23242
rect 9383 23208 9391 23242
rect 9339 23171 9391 23208
rect 9339 23137 9349 23171
rect 9383 23137 9391 23171
rect 9339 23125 9391 23137
rect 9943 23275 9951 23309
rect 9985 23275 9995 23309
rect 9943 23241 9995 23275
rect 9943 23207 9951 23241
rect 9985 23207 9995 23241
rect 9943 23195 9995 23207
rect 10025 23293 10079 23323
rect 10025 23259 10035 23293
rect 10069 23259 10079 23293
rect 10025 23195 10079 23259
rect 10109 23309 10161 23323
rect 10109 23275 10119 23309
rect 10153 23275 10161 23309
rect 10109 23241 10161 23275
rect 10215 23317 10267 23329
rect 10215 23283 10223 23317
rect 10257 23283 10267 23317
rect 10215 23245 10267 23283
rect 10297 23309 10352 23329
rect 10297 23275 10307 23309
rect 10341 23275 10352 23309
rect 10297 23245 10352 23275
rect 10382 23304 10447 23329
rect 10382 23270 10399 23304
rect 10433 23270 10447 23304
rect 10382 23245 10447 23270
rect 10477 23245 10550 23329
rect 10580 23317 10682 23329
rect 10580 23283 10638 23317
rect 10672 23283 10682 23317
rect 10580 23249 10682 23283
rect 10580 23245 10638 23249
rect 10109 23207 10119 23241
rect 10153 23207 10161 23241
rect 10109 23195 10161 23207
rect 10595 23215 10638 23245
rect 10672 23215 10682 23249
rect 10595 23179 10682 23215
rect 10712 23309 10777 23329
rect 10712 23275 10722 23309
rect 10756 23275 10777 23309
rect 10712 23245 10777 23275
rect 10807 23299 10861 23329
rect 10807 23265 10817 23299
rect 10851 23265 10861 23299
rect 10807 23245 10861 23265
rect 10891 23245 10975 23329
rect 11005 23309 11058 23329
rect 11005 23275 11016 23309
rect 11050 23275 11058 23309
rect 11005 23245 11058 23275
rect 11132 23317 11186 23329
rect 11132 23283 11140 23317
rect 11174 23283 11186 23317
rect 11132 23246 11186 23283
rect 10712 23179 10762 23245
rect 11132 23212 11140 23246
rect 11174 23212 11186 23246
rect 11132 23175 11186 23212
rect 11132 23141 11140 23175
rect 11174 23141 11186 23175
rect 11132 23129 11186 23141
rect 11216 23287 11270 23329
rect 11216 23253 11226 23287
rect 11260 23253 11270 23287
rect 11216 23207 11270 23253
rect 11216 23173 11226 23207
rect 11260 23173 11270 23207
rect 11216 23129 11270 23173
rect 11300 23311 11352 23329
rect 11300 23277 11310 23311
rect 11344 23277 11352 23311
rect 11300 23243 11352 23277
rect 11300 23209 11310 23243
rect 11344 23209 11352 23243
rect 11300 23175 11352 23209
rect 11406 23317 11458 23329
rect 11406 23283 11414 23317
rect 11448 23283 11458 23317
rect 11406 23249 11458 23283
rect 11406 23215 11414 23249
rect 11448 23215 11458 23249
rect 11406 23201 11458 23215
rect 11488 23317 11555 23329
rect 11488 23283 11511 23317
rect 11545 23283 11555 23317
rect 11488 23249 11555 23283
rect 11488 23215 11511 23249
rect 11545 23215 11555 23249
rect 11488 23201 11555 23215
rect 11300 23141 11310 23175
rect 11344 23141 11352 23175
rect 11300 23129 11352 23141
rect 11503 23181 11555 23201
rect 11503 23147 11511 23181
rect 11545 23147 11555 23181
rect 11503 23129 11555 23147
rect 11585 23317 11637 23329
rect 11585 23283 11595 23317
rect 11629 23283 11637 23317
rect 11585 23246 11637 23283
rect 11585 23212 11595 23246
rect 11629 23212 11637 23246
rect 11585 23175 11637 23212
rect 11585 23141 11595 23175
rect 11629 23141 11637 23175
rect 11585 23129 11637 23141
rect 12129 23301 12181 23315
rect 12129 23267 12137 23301
rect 12171 23267 12181 23301
rect 12129 23233 12181 23267
rect 12129 23199 12137 23233
rect 12171 23199 12181 23233
rect 12129 23187 12181 23199
rect 12211 23285 12265 23315
rect 12211 23251 12221 23285
rect 12255 23251 12265 23285
rect 12211 23187 12265 23251
rect 12295 23301 12347 23315
rect 12295 23267 12305 23301
rect 12339 23267 12347 23301
rect 12295 23233 12347 23267
rect 12401 23309 12453 23321
rect 12401 23275 12409 23309
rect 12443 23275 12453 23309
rect 12401 23237 12453 23275
rect 12483 23301 12538 23321
rect 12483 23267 12493 23301
rect 12527 23267 12538 23301
rect 12483 23237 12538 23267
rect 12568 23296 12633 23321
rect 12568 23262 12585 23296
rect 12619 23262 12633 23296
rect 12568 23237 12633 23262
rect 12663 23237 12736 23321
rect 12766 23309 12868 23321
rect 12766 23275 12824 23309
rect 12858 23275 12868 23309
rect 12766 23241 12868 23275
rect 12766 23237 12824 23241
rect 12295 23199 12305 23233
rect 12339 23199 12347 23233
rect 12295 23187 12347 23199
rect 12781 23207 12824 23237
rect 12858 23207 12868 23241
rect 12781 23171 12868 23207
rect 12898 23301 12963 23321
rect 12898 23267 12908 23301
rect 12942 23267 12963 23301
rect 12898 23237 12963 23267
rect 12993 23291 13047 23321
rect 12993 23257 13003 23291
rect 13037 23257 13047 23291
rect 12993 23237 13047 23257
rect 13077 23237 13161 23321
rect 13191 23301 13244 23321
rect 13191 23267 13202 23301
rect 13236 23267 13244 23301
rect 13191 23237 13244 23267
rect 13318 23309 13372 23321
rect 13318 23275 13326 23309
rect 13360 23275 13372 23309
rect 13318 23238 13372 23275
rect 12898 23171 12948 23237
rect 13318 23204 13326 23238
rect 13360 23204 13372 23238
rect 13318 23167 13372 23204
rect 13318 23133 13326 23167
rect 13360 23133 13372 23167
rect 13318 23121 13372 23133
rect 13402 23279 13456 23321
rect 13402 23245 13412 23279
rect 13446 23245 13456 23279
rect 13402 23199 13456 23245
rect 13402 23165 13412 23199
rect 13446 23165 13456 23199
rect 13402 23121 13456 23165
rect 13486 23303 13538 23321
rect 13486 23269 13496 23303
rect 13530 23269 13538 23303
rect 13486 23235 13538 23269
rect 13486 23201 13496 23235
rect 13530 23201 13538 23235
rect 13486 23167 13538 23201
rect 13592 23309 13644 23321
rect 13592 23275 13600 23309
rect 13634 23275 13644 23309
rect 13592 23241 13644 23275
rect 13592 23207 13600 23241
rect 13634 23207 13644 23241
rect 13592 23193 13644 23207
rect 13674 23309 13741 23321
rect 13674 23275 13697 23309
rect 13731 23275 13741 23309
rect 13674 23241 13741 23275
rect 13674 23207 13697 23241
rect 13731 23207 13741 23241
rect 13674 23193 13741 23207
rect 13486 23133 13496 23167
rect 13530 23133 13538 23167
rect 13486 23121 13538 23133
rect 13689 23173 13741 23193
rect 13689 23139 13697 23173
rect 13731 23139 13741 23173
rect 13689 23121 13741 23139
rect 13771 23309 13823 23321
rect 13771 23275 13781 23309
rect 13815 23275 13823 23309
rect 14375 23305 14427 23319
rect 13771 23238 13823 23275
rect 13771 23204 13781 23238
rect 13815 23204 13823 23238
rect 13771 23167 13823 23204
rect 13771 23133 13781 23167
rect 13815 23133 13823 23167
rect 13771 23121 13823 23133
rect 14375 23271 14383 23305
rect 14417 23271 14427 23305
rect 14375 23237 14427 23271
rect 14375 23203 14383 23237
rect 14417 23203 14427 23237
rect 14375 23191 14427 23203
rect 14457 23289 14511 23319
rect 14457 23255 14467 23289
rect 14501 23255 14511 23289
rect 14457 23191 14511 23255
rect 14541 23305 14593 23319
rect 14541 23271 14551 23305
rect 14585 23271 14593 23305
rect 14541 23237 14593 23271
rect 14647 23313 14699 23325
rect 14647 23279 14655 23313
rect 14689 23279 14699 23313
rect 14647 23241 14699 23279
rect 14729 23305 14784 23325
rect 14729 23271 14739 23305
rect 14773 23271 14784 23305
rect 14729 23241 14784 23271
rect 14814 23300 14879 23325
rect 14814 23266 14831 23300
rect 14865 23266 14879 23300
rect 14814 23241 14879 23266
rect 14909 23241 14982 23325
rect 15012 23313 15114 23325
rect 15012 23279 15070 23313
rect 15104 23279 15114 23313
rect 15012 23245 15114 23279
rect 15012 23241 15070 23245
rect 14541 23203 14551 23237
rect 14585 23203 14593 23237
rect 14541 23191 14593 23203
rect 15027 23211 15070 23241
rect 15104 23211 15114 23245
rect 15027 23175 15114 23211
rect 15144 23305 15209 23325
rect 15144 23271 15154 23305
rect 15188 23271 15209 23305
rect 15144 23241 15209 23271
rect 15239 23295 15293 23325
rect 15239 23261 15249 23295
rect 15283 23261 15293 23295
rect 15239 23241 15293 23261
rect 15323 23241 15407 23325
rect 15437 23305 15490 23325
rect 15437 23271 15448 23305
rect 15482 23271 15490 23305
rect 15437 23241 15490 23271
rect 15564 23313 15618 23325
rect 15564 23279 15572 23313
rect 15606 23279 15618 23313
rect 15564 23242 15618 23279
rect 15144 23175 15194 23241
rect 15564 23208 15572 23242
rect 15606 23208 15618 23242
rect 15564 23171 15618 23208
rect 15564 23137 15572 23171
rect 15606 23137 15618 23171
rect 15564 23125 15618 23137
rect 15648 23283 15702 23325
rect 15648 23249 15658 23283
rect 15692 23249 15702 23283
rect 15648 23203 15702 23249
rect 15648 23169 15658 23203
rect 15692 23169 15702 23203
rect 15648 23125 15702 23169
rect 15732 23307 15784 23325
rect 15732 23273 15742 23307
rect 15776 23273 15784 23307
rect 15732 23239 15784 23273
rect 15732 23205 15742 23239
rect 15776 23205 15784 23239
rect 15732 23171 15784 23205
rect 15838 23313 15890 23325
rect 15838 23279 15846 23313
rect 15880 23279 15890 23313
rect 15838 23245 15890 23279
rect 15838 23211 15846 23245
rect 15880 23211 15890 23245
rect 15838 23197 15890 23211
rect 15920 23313 15987 23325
rect 15920 23279 15943 23313
rect 15977 23279 15987 23313
rect 15920 23245 15987 23279
rect 15920 23211 15943 23245
rect 15977 23211 15987 23245
rect 15920 23197 15987 23211
rect 15732 23137 15742 23171
rect 15776 23137 15784 23171
rect 15732 23125 15784 23137
rect 15935 23177 15987 23197
rect 15935 23143 15943 23177
rect 15977 23143 15987 23177
rect 15935 23125 15987 23143
rect 16017 23313 16069 23325
rect 16017 23279 16027 23313
rect 16061 23279 16069 23313
rect 16017 23242 16069 23279
rect 16017 23208 16027 23242
rect 16061 23208 16069 23242
rect 16017 23171 16069 23208
rect 16017 23137 16027 23171
rect 16061 23137 16069 23171
rect 16017 23125 16069 23137
rect 16657 23305 16709 23319
rect 16657 23271 16665 23305
rect 16699 23271 16709 23305
rect 16657 23237 16709 23271
rect 16657 23203 16665 23237
rect 16699 23203 16709 23237
rect 16657 23191 16709 23203
rect 16739 23289 16793 23319
rect 16739 23255 16749 23289
rect 16783 23255 16793 23289
rect 16739 23191 16793 23255
rect 16823 23305 16875 23319
rect 16823 23271 16833 23305
rect 16867 23271 16875 23305
rect 16823 23237 16875 23271
rect 16929 23313 16981 23325
rect 16929 23279 16937 23313
rect 16971 23279 16981 23313
rect 16929 23241 16981 23279
rect 17011 23305 17066 23325
rect 17011 23271 17021 23305
rect 17055 23271 17066 23305
rect 17011 23241 17066 23271
rect 17096 23300 17161 23325
rect 17096 23266 17113 23300
rect 17147 23266 17161 23300
rect 17096 23241 17161 23266
rect 17191 23241 17264 23325
rect 17294 23313 17396 23325
rect 17294 23279 17352 23313
rect 17386 23279 17396 23313
rect 17294 23245 17396 23279
rect 17294 23241 17352 23245
rect 16823 23203 16833 23237
rect 16867 23203 16875 23237
rect 16823 23191 16875 23203
rect 17309 23211 17352 23241
rect 17386 23211 17396 23245
rect 17309 23175 17396 23211
rect 17426 23305 17491 23325
rect 17426 23271 17436 23305
rect 17470 23271 17491 23305
rect 17426 23241 17491 23271
rect 17521 23295 17575 23325
rect 17521 23261 17531 23295
rect 17565 23261 17575 23295
rect 17521 23241 17575 23261
rect 17605 23241 17689 23325
rect 17719 23305 17772 23325
rect 17719 23271 17730 23305
rect 17764 23271 17772 23305
rect 17719 23241 17772 23271
rect 17846 23313 17900 23325
rect 17846 23279 17854 23313
rect 17888 23279 17900 23313
rect 17846 23242 17900 23279
rect 17426 23175 17476 23241
rect 17846 23208 17854 23242
rect 17888 23208 17900 23242
rect 17846 23171 17900 23208
rect 17846 23137 17854 23171
rect 17888 23137 17900 23171
rect 17846 23125 17900 23137
rect 17930 23283 17984 23325
rect 17930 23249 17940 23283
rect 17974 23249 17984 23283
rect 17930 23203 17984 23249
rect 17930 23169 17940 23203
rect 17974 23169 17984 23203
rect 17930 23125 17984 23169
rect 18014 23307 18066 23325
rect 18014 23273 18024 23307
rect 18058 23273 18066 23307
rect 18014 23239 18066 23273
rect 18014 23205 18024 23239
rect 18058 23205 18066 23239
rect 18014 23171 18066 23205
rect 18120 23313 18172 23325
rect 18120 23279 18128 23313
rect 18162 23279 18172 23313
rect 18120 23245 18172 23279
rect 18120 23211 18128 23245
rect 18162 23211 18172 23245
rect 18120 23197 18172 23211
rect 18202 23313 18269 23325
rect 18202 23279 18225 23313
rect 18259 23279 18269 23313
rect 18202 23245 18269 23279
rect 18202 23211 18225 23245
rect 18259 23211 18269 23245
rect 18202 23197 18269 23211
rect 18014 23137 18024 23171
rect 18058 23137 18066 23171
rect 18014 23125 18066 23137
rect 18217 23177 18269 23197
rect 18217 23143 18225 23177
rect 18259 23143 18269 23177
rect 18217 23125 18269 23143
rect 18299 23313 18351 23325
rect 18299 23279 18309 23313
rect 18343 23279 18351 23313
rect 18299 23242 18351 23279
rect 18299 23208 18309 23242
rect 18343 23208 18351 23242
rect 18299 23171 18351 23208
rect 18299 23137 18309 23171
rect 18343 23137 18351 23171
rect 18299 23125 18351 23137
rect 9504 17479 9556 17497
rect 9504 17445 9512 17479
rect 9546 17445 9556 17479
rect 9504 17411 9556 17445
rect 9504 17377 9512 17411
rect 9546 17377 9556 17411
rect 9504 17343 9556 17377
rect 9504 17309 9512 17343
rect 9546 17309 9556 17343
rect 9504 17297 9556 17309
rect 9586 17479 9638 17497
rect 9586 17445 9596 17479
rect 9630 17445 9638 17479
rect 9586 17411 9638 17445
rect 9586 17377 9596 17411
rect 9630 17377 9638 17411
rect 9586 17343 9638 17377
rect 9586 17309 9596 17343
rect 9630 17309 9638 17343
rect 9586 17297 9638 17309
rect 15641 17331 15693 17349
rect 15641 17297 15649 17331
rect 15683 17297 15693 17331
rect 15641 17263 15693 17297
rect 15641 17229 15649 17263
rect 15683 17229 15693 17263
rect 15641 17195 15693 17229
rect 15641 17161 15649 17195
rect 15683 17161 15693 17195
rect 15641 17149 15693 17161
rect 15723 17331 15775 17349
rect 15723 17297 15733 17331
rect 15767 17297 15775 17331
rect 15723 17263 15775 17297
rect 15723 17229 15733 17263
rect 15767 17229 15775 17263
rect 15723 17195 15775 17229
rect 16419 17369 16471 17387
rect 16419 17335 16427 17369
rect 16461 17335 16471 17369
rect 16419 17301 16471 17335
rect 16419 17267 16427 17301
rect 16461 17267 16471 17301
rect 16419 17233 16471 17267
rect 15723 17161 15733 17195
rect 15767 17161 15775 17195
rect 16419 17199 16427 17233
rect 16461 17199 16471 17233
rect 16419 17187 16471 17199
rect 16501 17369 16553 17387
rect 16501 17335 16511 17369
rect 16545 17335 16553 17369
rect 16501 17301 16553 17335
rect 16501 17267 16511 17301
rect 16545 17267 16553 17301
rect 16501 17233 16553 17267
rect 16501 17199 16511 17233
rect 16545 17199 16553 17233
rect 17293 17371 17345 17389
rect 17293 17337 17301 17371
rect 17335 17337 17345 17371
rect 17293 17303 17345 17337
rect 17293 17269 17301 17303
rect 17335 17269 17345 17303
rect 17293 17235 17345 17269
rect 16501 17187 16553 17199
rect 17293 17201 17301 17235
rect 17335 17201 17345 17235
rect 17293 17189 17345 17201
rect 17375 17371 17427 17389
rect 17375 17337 17385 17371
rect 17419 17337 17427 17371
rect 17375 17303 17427 17337
rect 17375 17269 17385 17303
rect 17419 17269 17427 17303
rect 17375 17235 17427 17269
rect 17375 17201 17385 17235
rect 17419 17201 17427 17235
rect 17375 17189 17427 17201
rect 18061 17361 18113 17379
rect 18061 17327 18069 17361
rect 18103 17327 18113 17361
rect 18061 17293 18113 17327
rect 18061 17259 18069 17293
rect 18103 17259 18113 17293
rect 18061 17225 18113 17259
rect 18061 17191 18069 17225
rect 18103 17191 18113 17225
rect 18061 17179 18113 17191
rect 18143 17361 18195 17379
rect 18143 17327 18153 17361
rect 18187 17327 18195 17361
rect 18143 17293 18195 17327
rect 18143 17259 18153 17293
rect 18187 17259 18195 17293
rect 18143 17225 18195 17259
rect 18143 17191 18153 17225
rect 18187 17191 18195 17225
rect 19183 17363 19235 17381
rect 19183 17329 19191 17363
rect 19225 17329 19235 17363
rect 19183 17295 19235 17329
rect 19183 17261 19191 17295
rect 19225 17261 19235 17295
rect 19183 17227 19235 17261
rect 18143 17179 18195 17191
rect 19183 17193 19191 17227
rect 19225 17193 19235 17227
rect 19183 17181 19235 17193
rect 19265 17363 19317 17381
rect 19265 17329 19275 17363
rect 19309 17329 19317 17363
rect 19265 17295 19317 17329
rect 19265 17261 19275 17295
rect 19309 17261 19317 17295
rect 19265 17227 19317 17261
rect 19265 17193 19275 17227
rect 19309 17193 19317 17227
rect 20057 17365 20109 17383
rect 20057 17331 20065 17365
rect 20099 17331 20109 17365
rect 20057 17297 20109 17331
rect 20057 17263 20065 17297
rect 20099 17263 20109 17297
rect 20057 17229 20109 17263
rect 19265 17181 19317 17193
rect 20057 17195 20065 17229
rect 20099 17195 20109 17229
rect 20057 17183 20109 17195
rect 20139 17365 20191 17383
rect 20139 17331 20149 17365
rect 20183 17331 20191 17365
rect 20139 17297 20191 17331
rect 20139 17263 20149 17297
rect 20183 17263 20191 17297
rect 20139 17229 20191 17263
rect 20139 17195 20149 17229
rect 20183 17195 20191 17229
rect 20139 17183 20191 17195
rect 20825 17355 20877 17373
rect 20825 17321 20833 17355
rect 20867 17321 20877 17355
rect 20825 17287 20877 17321
rect 20825 17253 20833 17287
rect 20867 17253 20877 17287
rect 20825 17219 20877 17253
rect 20825 17185 20833 17219
rect 20867 17185 20877 17219
rect 15723 17149 15775 17161
rect 20825 17173 20877 17185
rect 20907 17355 20959 17373
rect 20907 17321 20917 17355
rect 20951 17321 20959 17355
rect 20907 17287 20959 17321
rect 20907 17253 20917 17287
rect 20951 17253 20959 17287
rect 20907 17219 20959 17253
rect 20907 17185 20917 17219
rect 20951 17185 20959 17219
rect 20907 17173 20959 17185
rect 21439 17353 21491 17371
rect 21439 17319 21447 17353
rect 21481 17319 21491 17353
rect 21439 17285 21491 17319
rect 21439 17251 21447 17285
rect 21481 17251 21491 17285
rect 21439 17217 21491 17251
rect 21439 17183 21447 17217
rect 21481 17183 21491 17217
rect 21439 17171 21491 17183
rect 21521 17353 21573 17371
rect 21521 17319 21531 17353
rect 21565 17319 21573 17353
rect 21521 17285 21573 17319
rect 21521 17251 21531 17285
rect 21565 17251 21573 17285
rect 21521 17217 21573 17251
rect 21521 17183 21531 17217
rect 21565 17183 21573 17217
rect 22313 17355 22365 17373
rect 22313 17321 22321 17355
rect 22355 17321 22365 17355
rect 22313 17287 22365 17321
rect 22313 17253 22321 17287
rect 22355 17253 22365 17287
rect 22313 17219 22365 17253
rect 21521 17171 21573 17183
rect 22313 17185 22321 17219
rect 22355 17185 22365 17219
rect 22313 17173 22365 17185
rect 22395 17355 22447 17373
rect 22395 17321 22405 17355
rect 22439 17321 22447 17355
rect 22395 17287 22447 17321
rect 22395 17253 22405 17287
rect 22439 17253 22447 17287
rect 22395 17219 22447 17253
rect 22395 17185 22405 17219
rect 22439 17185 22447 17219
rect 22395 17173 22447 17185
rect 23081 17345 23133 17363
rect 23081 17311 23089 17345
rect 23123 17311 23133 17345
rect 23081 17277 23133 17311
rect 23081 17243 23089 17277
rect 23123 17243 23133 17277
rect 23081 17209 23133 17243
rect 23081 17175 23089 17209
rect 23123 17175 23133 17209
rect 23081 17163 23133 17175
rect 23163 17345 23215 17363
rect 23163 17311 23173 17345
rect 23207 17311 23215 17345
rect 23163 17277 23215 17311
rect 23163 17243 23173 17277
rect 23207 17243 23215 17277
rect 23163 17209 23215 17243
rect 23163 17175 23173 17209
rect 23207 17175 23215 17209
rect 23163 17163 23215 17175
rect 16404 16635 16456 16647
rect 4503 16527 4555 16539
rect 4503 16493 4511 16527
rect 4545 16493 4555 16527
rect 4503 16459 4555 16493
rect 4503 16425 4511 16459
rect 4545 16425 4555 16459
rect 4503 16339 4555 16425
rect 4585 16339 4639 16539
rect 4669 16517 4723 16539
rect 4669 16483 4679 16517
rect 4713 16483 4723 16517
rect 4669 16449 4723 16483
rect 4669 16415 4679 16449
rect 4713 16415 4723 16449
rect 4669 16339 4723 16415
rect 4753 16517 4807 16539
rect 4753 16483 4763 16517
rect 4797 16483 4807 16517
rect 4753 16449 4807 16483
rect 4753 16415 4763 16449
rect 4797 16415 4807 16449
rect 4753 16339 4807 16415
rect 4837 16517 4889 16539
rect 4837 16483 4847 16517
rect 4881 16483 4889 16517
rect 4837 16339 4889 16483
rect 4943 16517 4995 16539
rect 4943 16483 4951 16517
rect 4985 16483 4995 16517
rect 4943 16449 4995 16483
rect 4943 16415 4951 16449
rect 4985 16415 4995 16449
rect 4943 16339 4995 16415
rect 5025 16519 5085 16539
rect 9369 16531 9421 16543
rect 5025 16485 5035 16519
rect 5069 16485 5085 16519
rect 5025 16451 5085 16485
rect 5025 16417 5035 16451
rect 5069 16417 5085 16451
rect 5025 16383 5085 16417
rect 5025 16349 5035 16383
rect 5069 16349 5085 16383
rect 9369 16497 9377 16531
rect 9411 16497 9421 16531
rect 9369 16463 9421 16497
rect 9369 16429 9377 16463
rect 9411 16429 9421 16463
rect 5025 16339 5085 16349
rect 9369 16343 9421 16429
rect 9451 16343 9505 16543
rect 9535 16521 9589 16543
rect 9535 16487 9545 16521
rect 9579 16487 9589 16521
rect 9535 16453 9589 16487
rect 9535 16419 9545 16453
rect 9579 16419 9589 16453
rect 9535 16343 9589 16419
rect 9619 16521 9673 16543
rect 9619 16487 9629 16521
rect 9663 16487 9673 16521
rect 9619 16453 9673 16487
rect 9619 16419 9629 16453
rect 9663 16419 9673 16453
rect 9619 16343 9673 16419
rect 9703 16521 9755 16543
rect 9703 16487 9713 16521
rect 9747 16487 9755 16521
rect 9703 16343 9755 16487
rect 9809 16521 9861 16543
rect 9809 16487 9817 16521
rect 9851 16487 9861 16521
rect 9809 16453 9861 16487
rect 9809 16419 9817 16453
rect 9851 16419 9861 16453
rect 9809 16343 9861 16419
rect 9891 16523 9951 16543
rect 9891 16489 9901 16523
rect 9935 16489 9951 16523
rect 9891 16455 9951 16489
rect 16404 16601 16412 16635
rect 16446 16601 16456 16635
rect 16404 16567 16456 16601
rect 16404 16533 16412 16567
rect 16446 16533 16456 16567
rect 16404 16499 16456 16533
rect 16404 16465 16412 16499
rect 16446 16465 16456 16499
rect 9891 16421 9901 16455
rect 9935 16421 9951 16455
rect 16404 16447 16456 16465
rect 16486 16635 16538 16647
rect 16486 16601 16496 16635
rect 16530 16601 16538 16635
rect 16486 16567 16538 16601
rect 16486 16533 16496 16567
rect 16530 16533 16538 16567
rect 16486 16499 16538 16533
rect 16486 16465 16496 16499
rect 16530 16465 16538 16499
rect 16486 16447 16538 16465
rect 17172 16625 17224 16637
rect 17172 16591 17180 16625
rect 17214 16591 17224 16625
rect 17172 16557 17224 16591
rect 17172 16523 17180 16557
rect 17214 16523 17224 16557
rect 17172 16489 17224 16523
rect 17172 16455 17180 16489
rect 17214 16455 17224 16489
rect 9891 16387 9951 16421
rect 17172 16437 17224 16455
rect 17254 16625 17306 16637
rect 17254 16591 17264 16625
rect 17298 16591 17306 16625
rect 18046 16627 18098 16639
rect 17254 16557 17306 16591
rect 17254 16523 17264 16557
rect 17298 16523 17306 16557
rect 17254 16489 17306 16523
rect 17254 16455 17264 16489
rect 17298 16455 17306 16489
rect 17254 16437 17306 16455
rect 18046 16593 18054 16627
rect 18088 16593 18098 16627
rect 18046 16559 18098 16593
rect 18046 16525 18054 16559
rect 18088 16525 18098 16559
rect 18046 16491 18098 16525
rect 18046 16457 18054 16491
rect 18088 16457 18098 16491
rect 18046 16439 18098 16457
rect 18128 16627 18180 16639
rect 18128 16593 18138 16627
rect 18172 16593 18180 16627
rect 18128 16559 18180 16593
rect 18128 16525 18138 16559
rect 18172 16525 18180 16559
rect 18128 16491 18180 16525
rect 18128 16457 18138 16491
rect 18172 16457 18180 16491
rect 18128 16439 18180 16457
rect 18660 16625 18712 16637
rect 18660 16591 18668 16625
rect 18702 16591 18712 16625
rect 18660 16557 18712 16591
rect 18660 16523 18668 16557
rect 18702 16523 18712 16557
rect 18660 16489 18712 16523
rect 18660 16455 18668 16489
rect 18702 16455 18712 16489
rect 9891 16353 9901 16387
rect 9935 16353 9951 16387
rect 9891 16343 9951 16353
rect 18660 16437 18712 16455
rect 18742 16625 18794 16637
rect 18742 16591 18752 16625
rect 18786 16591 18794 16625
rect 18742 16557 18794 16591
rect 18742 16523 18752 16557
rect 18786 16523 18794 16557
rect 18742 16489 18794 16523
rect 18742 16455 18752 16489
rect 18786 16455 18794 16489
rect 18742 16437 18794 16455
rect 19428 16615 19480 16627
rect 19428 16581 19436 16615
rect 19470 16581 19480 16615
rect 19428 16547 19480 16581
rect 19428 16513 19436 16547
rect 19470 16513 19480 16547
rect 19428 16479 19480 16513
rect 19428 16445 19436 16479
rect 19470 16445 19480 16479
rect 19428 16427 19480 16445
rect 19510 16615 19562 16627
rect 19510 16581 19520 16615
rect 19554 16581 19562 16615
rect 20302 16617 20354 16629
rect 19510 16547 19562 16581
rect 19510 16513 19520 16547
rect 19554 16513 19562 16547
rect 19510 16479 19562 16513
rect 19510 16445 19520 16479
rect 19554 16445 19562 16479
rect 19510 16427 19562 16445
rect 20302 16583 20310 16617
rect 20344 16583 20354 16617
rect 20302 16549 20354 16583
rect 20302 16515 20310 16549
rect 20344 16515 20354 16549
rect 20302 16481 20354 16515
rect 20302 16447 20310 16481
rect 20344 16447 20354 16481
rect 20302 16429 20354 16447
rect 20384 16617 20436 16629
rect 20384 16583 20394 16617
rect 20428 16583 20436 16617
rect 21424 16619 21476 16631
rect 20384 16549 20436 16583
rect 20384 16515 20394 16549
rect 20428 16515 20436 16549
rect 20384 16481 20436 16515
rect 20384 16447 20394 16481
rect 20428 16447 20436 16481
rect 20384 16429 20436 16447
rect 21424 16585 21432 16619
rect 21466 16585 21476 16619
rect 21424 16551 21476 16585
rect 21424 16517 21432 16551
rect 21466 16517 21476 16551
rect 21424 16483 21476 16517
rect 21424 16449 21432 16483
rect 21466 16449 21476 16483
rect 21424 16431 21476 16449
rect 21506 16619 21558 16631
rect 21506 16585 21516 16619
rect 21550 16585 21558 16619
rect 21506 16551 21558 16585
rect 21506 16517 21516 16551
rect 21550 16517 21558 16551
rect 21506 16483 21558 16517
rect 21506 16449 21516 16483
rect 21550 16449 21558 16483
rect 21506 16431 21558 16449
rect 22192 16609 22244 16621
rect 22192 16575 22200 16609
rect 22234 16575 22244 16609
rect 22192 16541 22244 16575
rect 22192 16507 22200 16541
rect 22234 16507 22244 16541
rect 22192 16473 22244 16507
rect 22192 16439 22200 16473
rect 22234 16439 22244 16473
rect 22192 16421 22244 16439
rect 22274 16609 22326 16621
rect 22274 16575 22284 16609
rect 22318 16575 22326 16609
rect 23066 16611 23118 16623
rect 22274 16541 22326 16575
rect 22274 16507 22284 16541
rect 22318 16507 22326 16541
rect 22274 16473 22326 16507
rect 22274 16439 22284 16473
rect 22318 16439 22326 16473
rect 22274 16421 22326 16439
rect 23066 16577 23074 16611
rect 23108 16577 23118 16611
rect 23066 16543 23118 16577
rect 23066 16509 23074 16543
rect 23108 16509 23118 16543
rect 23066 16475 23118 16509
rect 23066 16441 23074 16475
rect 23108 16441 23118 16475
rect 23066 16423 23118 16441
rect 23148 16611 23200 16623
rect 23148 16577 23158 16611
rect 23192 16577 23200 16611
rect 23148 16543 23200 16577
rect 23148 16509 23158 16543
rect 23192 16509 23200 16543
rect 23148 16475 23200 16509
rect 23148 16441 23158 16475
rect 23192 16441 23200 16475
rect 23148 16423 23200 16441
rect 4821 15783 4873 15795
rect 4821 15753 4829 15783
rect 4625 15741 4681 15753
rect 4625 15707 4637 15741
rect 4671 15707 4681 15741
rect 4625 15669 4681 15707
rect 4711 15741 4765 15753
rect 4711 15707 4721 15741
rect 4755 15707 4765 15741
rect 4711 15669 4765 15707
rect 4795 15749 4829 15753
rect 4863 15749 4873 15783
rect 4795 15715 4873 15749
rect 4795 15681 4829 15715
rect 4863 15681 4873 15715
rect 4795 15669 4873 15681
rect 4811 15595 4873 15669
rect 4903 15783 4998 15795
rect 9687 15787 9739 15799
rect 4903 15749 4933 15783
rect 4967 15749 4998 15783
rect 4903 15715 4998 15749
rect 4903 15681 4933 15715
rect 4967 15681 4998 15715
rect 9687 15757 9695 15787
rect 4903 15595 4998 15681
rect 6635 15673 6687 15685
rect 6635 15639 6643 15673
rect 6677 15639 6687 15673
rect 6635 15601 6687 15639
rect 6717 15665 6787 15685
rect 6717 15631 6735 15665
rect 6769 15631 6787 15665
rect 6717 15601 6787 15631
rect 6817 15673 6891 15685
rect 6817 15639 6837 15673
rect 6871 15639 6891 15673
rect 6817 15601 6891 15639
rect 6921 15665 6977 15685
rect 6921 15631 6932 15665
rect 6966 15631 6977 15665
rect 6921 15601 6977 15631
rect 7007 15673 7143 15685
rect 7007 15639 7083 15673
rect 7117 15639 7143 15673
rect 7007 15605 7143 15639
rect 7007 15601 7083 15605
rect 7026 15571 7083 15601
rect 7117 15571 7143 15605
rect 7026 15485 7143 15571
rect 7173 15673 7225 15685
rect 7173 15639 7183 15673
rect 7217 15639 7225 15673
rect 7173 15605 7225 15639
rect 7173 15571 7183 15605
rect 7217 15571 7225 15605
rect 7173 15537 7225 15571
rect 7173 15503 7183 15537
rect 7217 15503 7225 15537
rect 7173 15485 7225 15503
rect 9491 15745 9547 15757
rect 9491 15711 9503 15745
rect 9537 15711 9547 15745
rect 9491 15673 9547 15711
rect 9577 15745 9631 15757
rect 9577 15711 9587 15745
rect 9621 15711 9631 15745
rect 9577 15673 9631 15711
rect 9661 15753 9695 15757
rect 9729 15753 9739 15787
rect 9661 15719 9739 15753
rect 9661 15685 9695 15719
rect 9729 15685 9739 15719
rect 9661 15673 9739 15685
rect 9677 15599 9739 15673
rect 9769 15787 9864 15799
rect 9769 15753 9799 15787
rect 9833 15753 9864 15787
rect 9769 15719 9864 15753
rect 9769 15685 9799 15719
rect 9833 15685 9864 15719
rect 9769 15599 9864 15685
rect 11501 15677 11553 15689
rect 11501 15643 11509 15677
rect 11543 15643 11553 15677
rect 11501 15605 11553 15643
rect 11583 15669 11653 15689
rect 11583 15635 11601 15669
rect 11635 15635 11653 15669
rect 11583 15605 11653 15635
rect 11683 15677 11757 15689
rect 11683 15643 11703 15677
rect 11737 15643 11757 15677
rect 11683 15605 11757 15643
rect 11787 15669 11843 15689
rect 11787 15635 11798 15669
rect 11832 15635 11843 15669
rect 11787 15605 11843 15635
rect 11873 15677 12009 15689
rect 11873 15643 11949 15677
rect 11983 15643 12009 15677
rect 11873 15609 12009 15643
rect 11873 15605 11949 15609
rect 11892 15575 11949 15605
rect 11983 15575 12009 15609
rect 11892 15489 12009 15575
rect 12039 15677 12091 15689
rect 12039 15643 12049 15677
rect 12083 15643 12091 15677
rect 12039 15609 12091 15643
rect 12039 15575 12049 15609
rect 12083 15575 12091 15609
rect 12039 15541 12091 15575
rect 12039 15507 12049 15541
rect 12083 15507 12091 15541
rect 12039 15489 12091 15507
rect 6005 15173 6057 15185
rect 6005 15143 6013 15173
rect 5809 15131 5865 15143
rect 5809 15097 5821 15131
rect 5855 15097 5865 15131
rect 5809 15059 5865 15097
rect 5895 15131 5949 15143
rect 5895 15097 5905 15131
rect 5939 15097 5949 15131
rect 5895 15059 5949 15097
rect 5979 15139 6013 15143
rect 6047 15139 6057 15173
rect 5979 15105 6057 15139
rect 5979 15071 6013 15105
rect 6047 15071 6057 15105
rect 5979 15059 6057 15071
rect 4513 14963 4565 14975
rect 4513 14929 4521 14963
rect 4555 14929 4565 14963
rect 4513 14895 4565 14929
rect 4513 14861 4521 14895
rect 4555 14861 4565 14895
rect 4513 14775 4565 14861
rect 4595 14775 4649 14975
rect 4679 14953 4733 14975
rect 4679 14919 4689 14953
rect 4723 14919 4733 14953
rect 4679 14885 4733 14919
rect 4679 14851 4689 14885
rect 4723 14851 4733 14885
rect 4679 14775 4733 14851
rect 4763 14953 4817 14975
rect 4763 14919 4773 14953
rect 4807 14919 4817 14953
rect 4763 14885 4817 14919
rect 4763 14851 4773 14885
rect 4807 14851 4817 14885
rect 4763 14775 4817 14851
rect 4847 14953 4899 14975
rect 4847 14919 4857 14953
rect 4891 14919 4899 14953
rect 4847 14775 4899 14919
rect 4953 14953 5005 14975
rect 4953 14919 4961 14953
rect 4995 14919 5005 14953
rect 4953 14885 5005 14919
rect 4953 14851 4961 14885
rect 4995 14851 5005 14885
rect 4953 14775 5005 14851
rect 5035 14955 5095 14975
rect 5035 14921 5045 14955
rect 5079 14921 5095 14955
rect 5035 14887 5095 14921
rect 5035 14853 5045 14887
rect 5079 14853 5095 14887
rect 5035 14819 5095 14853
rect 5995 14985 6057 15059
rect 6087 15173 6182 15185
rect 10871 15177 10923 15189
rect 6087 15139 6117 15173
rect 6151 15139 6182 15173
rect 6087 15105 6182 15139
rect 6087 15071 6117 15105
rect 6151 15071 6182 15105
rect 6087 14985 6182 15071
rect 10871 15147 10879 15177
rect 10675 15135 10731 15147
rect 10675 15101 10687 15135
rect 10721 15101 10731 15135
rect 10675 15063 10731 15101
rect 10761 15135 10815 15147
rect 10761 15101 10771 15135
rect 10805 15101 10815 15135
rect 10761 15063 10815 15101
rect 10845 15143 10879 15147
rect 10913 15143 10923 15177
rect 10845 15109 10923 15143
rect 10845 15075 10879 15109
rect 10913 15075 10923 15109
rect 10845 15063 10923 15075
rect 9379 14967 9431 14979
rect 5035 14785 5045 14819
rect 5079 14785 5095 14819
rect 5035 14775 5095 14785
rect 9379 14933 9387 14967
rect 9421 14933 9431 14967
rect 9379 14899 9431 14933
rect 9379 14865 9387 14899
rect 9421 14865 9431 14899
rect 9379 14779 9431 14865
rect 9461 14779 9515 14979
rect 9545 14957 9599 14979
rect 9545 14923 9555 14957
rect 9589 14923 9599 14957
rect 9545 14889 9599 14923
rect 9545 14855 9555 14889
rect 9589 14855 9599 14889
rect 9545 14779 9599 14855
rect 9629 14957 9683 14979
rect 9629 14923 9639 14957
rect 9673 14923 9683 14957
rect 9629 14889 9683 14923
rect 9629 14855 9639 14889
rect 9673 14855 9683 14889
rect 9629 14779 9683 14855
rect 9713 14957 9765 14979
rect 9713 14923 9723 14957
rect 9757 14923 9765 14957
rect 9713 14779 9765 14923
rect 9819 14957 9871 14979
rect 9819 14923 9827 14957
rect 9861 14923 9871 14957
rect 9819 14889 9871 14923
rect 9819 14855 9827 14889
rect 9861 14855 9871 14889
rect 9819 14779 9871 14855
rect 9901 14959 9961 14979
rect 9901 14925 9911 14959
rect 9945 14925 9961 14959
rect 9901 14891 9961 14925
rect 9901 14857 9911 14891
rect 9945 14857 9961 14891
rect 9901 14823 9961 14857
rect 10861 14989 10923 15063
rect 10953 15177 11048 15189
rect 10953 15143 10983 15177
rect 11017 15143 11048 15177
rect 10953 15109 11048 15143
rect 10953 15075 10983 15109
rect 11017 15075 11048 15109
rect 10953 14989 11048 15075
rect 9901 14789 9911 14823
rect 9945 14789 9961 14823
rect 9901 14779 9961 14789
rect 23511 14765 23563 14785
rect 23511 14731 23519 14765
rect 23553 14731 23563 14765
rect 23511 14701 23563 14731
rect 23593 14773 23647 14785
rect 23593 14739 23603 14773
rect 23637 14739 23647 14773
rect 23593 14701 23647 14739
rect 23677 14765 23729 14785
rect 23677 14731 23687 14765
rect 23721 14731 23729 14765
rect 24055 14765 24107 14785
rect 23677 14701 23729 14731
rect 23783 14697 23835 14735
rect 23783 14663 23791 14697
rect 23825 14663 23835 14697
rect 23783 14651 23835 14663
rect 23865 14713 23919 14735
rect 23865 14679 23875 14713
rect 23909 14679 23919 14713
rect 23865 14651 23919 14679
rect 23949 14709 23999 14735
rect 24055 14731 24063 14765
rect 24097 14731 24107 14765
rect 24055 14719 24107 14731
rect 23949 14697 24001 14709
rect 24057 14701 24107 14719
rect 24137 14773 24189 14785
rect 24137 14739 24147 14773
rect 24181 14739 24189 14773
rect 24137 14727 24189 14739
rect 24422 14735 24472 14785
rect 24137 14701 24187 14727
rect 24243 14709 24293 14735
rect 23949 14663 23959 14697
rect 23993 14663 24001 14697
rect 23949 14651 24001 14663
rect 24241 14697 24293 14709
rect 24241 14663 24249 14697
rect 24283 14663 24293 14697
rect 24241 14651 24293 14663
rect 24323 14713 24377 14735
rect 24323 14679 24333 14713
rect 24367 14679 24377 14713
rect 24323 14651 24377 14679
rect 24407 14701 24472 14735
rect 24502 14773 24556 14785
rect 24502 14739 24512 14773
rect 24546 14739 24556 14773
rect 24502 14701 24556 14739
rect 24586 14765 24638 14785
rect 24586 14731 24596 14765
rect 24630 14731 24638 14765
rect 24586 14701 24638 14731
rect 24692 14773 24744 14785
rect 24692 14739 24700 14773
rect 24734 14739 24744 14773
rect 24692 14701 24744 14739
rect 24774 14765 24826 14785
rect 24774 14731 24784 14765
rect 24818 14731 24826 14765
rect 24774 14701 24826 14731
rect 24880 14765 24932 14785
rect 24880 14731 24888 14765
rect 24922 14731 24932 14765
rect 24880 14701 24932 14731
rect 24962 14773 25014 14785
rect 24962 14739 24972 14773
rect 25006 14739 25014 14773
rect 24962 14738 25014 14739
rect 25255 14773 25307 14785
rect 25255 14739 25263 14773
rect 25297 14739 25307 14773
rect 24962 14701 25029 14738
rect 24407 14651 24457 14701
rect 24977 14654 25029 14701
rect 25059 14713 25187 14738
rect 25059 14679 25069 14713
rect 25103 14679 25187 14713
rect 25059 14654 25187 14679
rect 25255 14585 25307 14739
rect 25337 14765 25389 14785
rect 25337 14731 25347 14765
rect 25381 14731 25389 14765
rect 25337 14585 25389 14731
rect 4831 14219 4883 14231
rect 4831 14189 4839 14219
rect 4635 14177 4691 14189
rect 4635 14143 4647 14177
rect 4681 14143 4691 14177
rect 4635 14105 4691 14143
rect 4721 14177 4775 14189
rect 4721 14143 4731 14177
rect 4765 14143 4775 14177
rect 4721 14105 4775 14143
rect 4805 14185 4839 14189
rect 4873 14185 4883 14219
rect 4805 14151 4883 14185
rect 4805 14117 4839 14151
rect 4873 14117 4883 14151
rect 4805 14105 4883 14117
rect 4821 14031 4883 14105
rect 4913 14219 5008 14231
rect 4913 14185 4943 14219
rect 4977 14185 5008 14219
rect 5851 14207 5903 14219
rect 4913 14151 5008 14185
rect 4913 14117 4943 14151
rect 4977 14117 5008 14151
rect 4913 14031 5008 14117
rect 5851 14173 5859 14207
rect 5893 14173 5903 14207
rect 5851 14135 5903 14173
rect 5933 14199 6003 14219
rect 5933 14165 5951 14199
rect 5985 14165 6003 14199
rect 5933 14135 6003 14165
rect 6033 14207 6107 14219
rect 6033 14173 6053 14207
rect 6087 14173 6107 14207
rect 6033 14135 6107 14173
rect 6137 14199 6193 14219
rect 6137 14165 6148 14199
rect 6182 14165 6193 14199
rect 6137 14135 6193 14165
rect 6223 14207 6359 14219
rect 6223 14173 6299 14207
rect 6333 14173 6359 14207
rect 6223 14139 6359 14173
rect 6223 14135 6299 14139
rect 6242 14105 6299 14135
rect 6333 14105 6359 14139
rect 6242 14019 6359 14105
rect 6389 14207 6441 14219
rect 6389 14173 6399 14207
rect 6433 14173 6441 14207
rect 9697 14223 9749 14235
rect 8110 14191 8163 14203
rect 6389 14139 6441 14173
rect 6389 14105 6399 14139
rect 6433 14105 6441 14139
rect 8110 14157 8118 14191
rect 8152 14157 8163 14191
rect 6389 14071 6441 14105
rect 8110 14123 8163 14157
rect 8110 14089 8118 14123
rect 8152 14089 8163 14123
rect 8110 14087 8163 14089
rect 6389 14037 6399 14071
rect 6433 14037 6441 14071
rect 6389 14019 6441 14037
rect 7749 14060 7801 14087
rect 7749 14026 7757 14060
rect 7791 14026 7801 14060
rect 7749 14003 7801 14026
rect 7831 14003 7897 14087
rect 7927 14003 7969 14087
rect 7999 14003 8065 14087
rect 8095 14003 8163 14087
rect 8193 14160 8247 14203
rect 8193 14126 8203 14160
rect 8237 14126 8247 14160
rect 8193 14092 8247 14126
rect 8193 14058 8203 14092
rect 8237 14058 8247 14092
rect 8193 14003 8247 14058
rect 9697 14193 9705 14223
rect 9501 14181 9557 14193
rect 9501 14147 9513 14181
rect 9547 14147 9557 14181
rect 9501 14109 9557 14147
rect 9587 14181 9641 14193
rect 9587 14147 9597 14181
rect 9631 14147 9641 14181
rect 9587 14109 9641 14147
rect 9671 14189 9705 14193
rect 9739 14189 9749 14223
rect 9671 14155 9749 14189
rect 9671 14121 9705 14155
rect 9739 14121 9749 14155
rect 9671 14109 9749 14121
rect 7031 13817 7083 13845
rect 7031 13783 7039 13817
rect 7073 13783 7083 13817
rect 7031 13749 7083 13783
rect 7031 13729 7039 13749
rect 6862 13697 6914 13729
rect 6862 13663 6870 13697
rect 6904 13663 6914 13697
rect 6862 13645 6914 13663
rect 6944 13645 6986 13729
rect 7016 13715 7039 13729
rect 7073 13715 7083 13749
rect 7016 13645 7083 13715
rect 7113 13833 7181 13845
rect 9687 14035 9749 14109
rect 9779 14223 9874 14235
rect 9779 14189 9809 14223
rect 9843 14189 9874 14223
rect 10717 14211 10769 14223
rect 9779 14155 9874 14189
rect 9779 14121 9809 14155
rect 9843 14121 9874 14155
rect 9779 14035 9874 14121
rect 10717 14177 10725 14211
rect 10759 14177 10769 14211
rect 10717 14139 10769 14177
rect 10799 14203 10869 14223
rect 10799 14169 10817 14203
rect 10851 14169 10869 14203
rect 10799 14139 10869 14169
rect 10899 14211 10973 14223
rect 10899 14177 10919 14211
rect 10953 14177 10973 14211
rect 10899 14139 10973 14177
rect 11003 14203 11059 14223
rect 11003 14169 11014 14203
rect 11048 14169 11059 14203
rect 11003 14139 11059 14169
rect 11089 14211 11225 14223
rect 11089 14177 11165 14211
rect 11199 14177 11225 14211
rect 11089 14143 11225 14177
rect 11089 14139 11165 14143
rect 11108 14109 11165 14139
rect 11199 14109 11225 14143
rect 11108 14023 11225 14109
rect 11255 14211 11307 14223
rect 11255 14177 11265 14211
rect 11299 14177 11307 14211
rect 12976 14195 13029 14207
rect 11255 14143 11307 14177
rect 11255 14109 11265 14143
rect 11299 14109 11307 14143
rect 12976 14161 12984 14195
rect 13018 14161 13029 14195
rect 11255 14075 11307 14109
rect 12976 14127 13029 14161
rect 12976 14093 12984 14127
rect 13018 14093 13029 14127
rect 12976 14091 13029 14093
rect 11255 14041 11265 14075
rect 11299 14041 11307 14075
rect 11255 14023 11307 14041
rect 12615 14064 12667 14091
rect 12615 14030 12623 14064
rect 12657 14030 12667 14064
rect 12615 14007 12667 14030
rect 12697 14007 12763 14091
rect 12793 14007 12835 14091
rect 12865 14007 12931 14091
rect 12961 14007 13029 14091
rect 13059 14164 13113 14207
rect 13059 14130 13069 14164
rect 13103 14130 13113 14164
rect 13059 14096 13113 14130
rect 13059 14062 13069 14096
rect 13103 14062 13113 14096
rect 13059 14007 13113 14062
rect 7113 13799 7139 13833
rect 7173 13799 7181 13833
rect 7113 13765 7181 13799
rect 7113 13731 7139 13765
rect 7173 13731 7181 13765
rect 7113 13645 7181 13731
rect 11897 13821 11949 13849
rect 11897 13787 11905 13821
rect 11939 13787 11949 13821
rect 11897 13753 11949 13787
rect 11897 13733 11905 13753
rect 11728 13701 11780 13733
rect 11728 13667 11736 13701
rect 11770 13667 11780 13701
rect 11728 13649 11780 13667
rect 11810 13649 11852 13733
rect 11882 13719 11905 13733
rect 11939 13719 11949 13753
rect 11882 13649 11949 13719
rect 11979 13837 12047 13849
rect 11979 13803 12005 13837
rect 12039 13803 12047 13837
rect 11979 13769 12047 13803
rect 11979 13735 12005 13769
rect 12039 13735 12047 13769
rect 11979 13649 12047 13735
rect 4505 13295 4557 13307
rect 4505 13261 4513 13295
rect 4547 13261 4557 13295
rect 4505 13227 4557 13261
rect 4505 13193 4513 13227
rect 4547 13193 4557 13227
rect 4505 13107 4557 13193
rect 4587 13107 4641 13307
rect 4671 13285 4725 13307
rect 4671 13251 4681 13285
rect 4715 13251 4725 13285
rect 4671 13217 4725 13251
rect 4671 13183 4681 13217
rect 4715 13183 4725 13217
rect 4671 13107 4725 13183
rect 4755 13285 4809 13307
rect 4755 13251 4765 13285
rect 4799 13251 4809 13285
rect 4755 13217 4809 13251
rect 4755 13183 4765 13217
rect 4799 13183 4809 13217
rect 4755 13107 4809 13183
rect 4839 13285 4891 13307
rect 4839 13251 4849 13285
rect 4883 13251 4891 13285
rect 4839 13107 4891 13251
rect 4945 13285 4997 13307
rect 4945 13251 4953 13285
rect 4987 13251 4997 13285
rect 4945 13217 4997 13251
rect 4945 13183 4953 13217
rect 4987 13183 4997 13217
rect 4945 13107 4997 13183
rect 5027 13287 5087 13307
rect 5027 13253 5037 13287
rect 5071 13253 5087 13287
rect 5027 13219 5087 13253
rect 5027 13185 5037 13219
rect 5071 13185 5087 13219
rect 6247 13365 6299 13377
rect 6247 13331 6255 13365
rect 6289 13331 6299 13365
rect 6247 13318 6299 13331
rect 6249 13264 6299 13318
rect 5975 13226 6027 13264
rect 5975 13192 5983 13226
rect 6017 13192 6027 13226
rect 5027 13151 5087 13185
rect 5975 13180 6027 13192
rect 6057 13256 6111 13264
rect 6057 13222 6067 13256
rect 6101 13222 6111 13256
rect 6057 13180 6111 13222
rect 6141 13237 6204 13264
rect 6141 13203 6160 13237
rect 6194 13203 6204 13237
rect 6141 13180 6204 13203
rect 6234 13180 6299 13264
rect 5027 13117 5037 13151
rect 5071 13117 5087 13151
rect 5027 13107 5087 13117
rect 6249 13177 6299 13180
rect 6329 13351 6381 13377
rect 6329 13317 6339 13351
rect 6373 13317 6381 13351
rect 6329 13283 6381 13317
rect 9371 13299 9423 13311
rect 6329 13249 6339 13283
rect 6373 13249 6381 13283
rect 6329 13177 6381 13249
rect 9371 13265 9379 13299
rect 9413 13265 9423 13299
rect 9371 13231 9423 13265
rect 9371 13197 9379 13231
rect 9413 13197 9423 13231
rect 9371 13111 9423 13197
rect 9453 13111 9507 13311
rect 9537 13289 9591 13311
rect 9537 13255 9547 13289
rect 9581 13255 9591 13289
rect 9537 13221 9591 13255
rect 9537 13187 9547 13221
rect 9581 13187 9591 13221
rect 9537 13111 9591 13187
rect 9621 13289 9675 13311
rect 9621 13255 9631 13289
rect 9665 13255 9675 13289
rect 9621 13221 9675 13255
rect 9621 13187 9631 13221
rect 9665 13187 9675 13221
rect 9621 13111 9675 13187
rect 9705 13289 9757 13311
rect 9705 13255 9715 13289
rect 9749 13255 9757 13289
rect 9705 13111 9757 13255
rect 9811 13289 9863 13311
rect 9811 13255 9819 13289
rect 9853 13255 9863 13289
rect 9811 13221 9863 13255
rect 9811 13187 9819 13221
rect 9853 13187 9863 13221
rect 9811 13111 9863 13187
rect 9893 13291 9953 13311
rect 9893 13257 9903 13291
rect 9937 13257 9953 13291
rect 9893 13223 9953 13257
rect 9893 13189 9903 13223
rect 9937 13189 9953 13223
rect 11113 13369 11165 13381
rect 11113 13335 11121 13369
rect 11155 13335 11165 13369
rect 11113 13322 11165 13335
rect 11115 13268 11165 13322
rect 10841 13230 10893 13268
rect 10841 13196 10849 13230
rect 10883 13196 10893 13230
rect 9893 13155 9953 13189
rect 10841 13184 10893 13196
rect 10923 13260 10977 13268
rect 10923 13226 10933 13260
rect 10967 13226 10977 13260
rect 10923 13184 10977 13226
rect 11007 13241 11070 13268
rect 11007 13207 11026 13241
rect 11060 13207 11070 13241
rect 11007 13184 11070 13207
rect 11100 13184 11165 13268
rect 9893 13121 9903 13155
rect 9937 13121 9953 13155
rect 9893 13111 9953 13121
rect 11115 13181 11165 13184
rect 11195 13355 11247 13381
rect 11195 13321 11205 13355
rect 11239 13321 11247 13355
rect 11195 13287 11247 13321
rect 11195 13253 11205 13287
rect 11239 13253 11247 13287
rect 11195 13181 11247 13253
rect 4823 12551 4875 12563
rect 4823 12521 4831 12551
rect 4627 12509 4683 12521
rect 4627 12475 4639 12509
rect 4673 12475 4683 12509
rect 4627 12437 4683 12475
rect 4713 12509 4767 12521
rect 4713 12475 4723 12509
rect 4757 12475 4767 12509
rect 4713 12437 4767 12475
rect 4797 12517 4831 12521
rect 4865 12517 4875 12551
rect 4797 12483 4875 12517
rect 4797 12449 4831 12483
rect 4865 12449 4875 12483
rect 4797 12437 4875 12449
rect 4813 12363 4875 12437
rect 4905 12551 5000 12563
rect 9689 12555 9741 12567
rect 4905 12517 4935 12551
rect 4969 12517 5000 12551
rect 4905 12483 5000 12517
rect 4905 12449 4935 12483
rect 4969 12449 5000 12483
rect 4905 12363 5000 12449
rect 9689 12525 9697 12555
rect 9493 12513 9549 12525
rect 9493 12479 9505 12513
rect 9539 12479 9549 12513
rect 9493 12441 9549 12479
rect 9579 12513 9633 12525
rect 9579 12479 9589 12513
rect 9623 12479 9633 12513
rect 9579 12441 9633 12479
rect 9663 12521 9697 12525
rect 9731 12521 9741 12555
rect 9663 12487 9741 12521
rect 9663 12453 9697 12487
rect 9731 12453 9741 12487
rect 9663 12441 9741 12453
rect 6199 12345 6251 12357
rect 6199 12315 6207 12345
rect 6003 12303 6059 12315
rect 6003 12269 6015 12303
rect 6049 12269 6059 12303
rect 6003 12231 6059 12269
rect 6089 12303 6143 12315
rect 6089 12269 6099 12303
rect 6133 12269 6143 12303
rect 6089 12231 6143 12269
rect 6173 12311 6207 12315
rect 6241 12311 6251 12345
rect 6173 12277 6251 12311
rect 6173 12243 6207 12277
rect 6241 12243 6251 12277
rect 6173 12231 6251 12243
rect 6189 12157 6251 12231
rect 6281 12345 6376 12357
rect 6281 12311 6311 12345
rect 6345 12311 6376 12345
rect 6281 12277 6376 12311
rect 6281 12243 6311 12277
rect 6345 12243 6376 12277
rect 6281 12157 6376 12243
rect 9679 12367 9741 12441
rect 9771 12555 9866 12567
rect 9771 12521 9801 12555
rect 9835 12521 9866 12555
rect 9771 12487 9866 12521
rect 9771 12453 9801 12487
rect 9835 12453 9866 12487
rect 9771 12367 9866 12453
rect 11065 12349 11117 12361
rect 11065 12319 11073 12349
rect 10869 12307 10925 12319
rect 10869 12273 10881 12307
rect 10915 12273 10925 12307
rect 10869 12235 10925 12273
rect 10955 12307 11009 12319
rect 10955 12273 10965 12307
rect 10999 12273 11009 12307
rect 10955 12235 11009 12273
rect 11039 12315 11073 12319
rect 11107 12315 11117 12349
rect 11039 12281 11117 12315
rect 11039 12247 11073 12281
rect 11107 12247 11117 12281
rect 11039 12235 11117 12247
rect 11055 12161 11117 12235
rect 11147 12349 11242 12361
rect 11147 12315 11177 12349
rect 11211 12315 11242 12349
rect 11147 12281 11242 12315
rect 11147 12247 11177 12281
rect 11211 12247 11242 12281
rect 11147 12161 11242 12247
rect 4515 11731 4567 11743
rect 4515 11697 4523 11731
rect 4557 11697 4567 11731
rect 4515 11663 4567 11697
rect 4515 11629 4523 11663
rect 4557 11629 4567 11663
rect 4515 11543 4567 11629
rect 4597 11543 4651 11743
rect 4681 11721 4735 11743
rect 4681 11687 4691 11721
rect 4725 11687 4735 11721
rect 4681 11653 4735 11687
rect 4681 11619 4691 11653
rect 4725 11619 4735 11653
rect 4681 11543 4735 11619
rect 4765 11721 4819 11743
rect 4765 11687 4775 11721
rect 4809 11687 4819 11721
rect 4765 11653 4819 11687
rect 4765 11619 4775 11653
rect 4809 11619 4819 11653
rect 4765 11543 4819 11619
rect 4849 11721 4901 11743
rect 4849 11687 4859 11721
rect 4893 11687 4901 11721
rect 4849 11543 4901 11687
rect 4955 11721 5007 11743
rect 4955 11687 4963 11721
rect 4997 11687 5007 11721
rect 4955 11653 5007 11687
rect 4955 11619 4963 11653
rect 4997 11619 5007 11653
rect 4955 11543 5007 11619
rect 5037 11723 5097 11743
rect 9381 11735 9433 11747
rect 5037 11689 5047 11723
rect 5081 11689 5097 11723
rect 5037 11655 5097 11689
rect 5037 11621 5047 11655
rect 5081 11621 5097 11655
rect 5037 11587 5097 11621
rect 5037 11553 5047 11587
rect 5081 11553 5097 11587
rect 9381 11701 9389 11735
rect 9423 11701 9433 11735
rect 9381 11667 9433 11701
rect 9381 11633 9389 11667
rect 9423 11633 9433 11667
rect 5037 11543 5097 11553
rect 9381 11547 9433 11633
rect 9463 11547 9517 11747
rect 9547 11725 9601 11747
rect 9547 11691 9557 11725
rect 9591 11691 9601 11725
rect 9547 11657 9601 11691
rect 9547 11623 9557 11657
rect 9591 11623 9601 11657
rect 9547 11547 9601 11623
rect 9631 11725 9685 11747
rect 9631 11691 9641 11725
rect 9675 11691 9685 11725
rect 9631 11657 9685 11691
rect 9631 11623 9641 11657
rect 9675 11623 9685 11657
rect 9631 11547 9685 11623
rect 9715 11725 9767 11747
rect 9715 11691 9725 11725
rect 9759 11691 9767 11725
rect 9715 11547 9767 11691
rect 9821 11725 9873 11747
rect 9821 11691 9829 11725
rect 9863 11691 9873 11725
rect 9821 11657 9873 11691
rect 9821 11623 9829 11657
rect 9863 11623 9873 11657
rect 9821 11547 9873 11623
rect 9903 11727 9963 11747
rect 9903 11693 9913 11727
rect 9947 11693 9963 11727
rect 9903 11659 9963 11693
rect 9903 11625 9913 11659
rect 9947 11625 9963 11659
rect 9903 11591 9963 11625
rect 9903 11557 9913 11591
rect 9947 11557 9963 11591
rect 9903 11547 9963 11557
rect 4833 10987 4885 10999
rect 4833 10957 4841 10987
rect 4637 10945 4693 10957
rect 4637 10911 4649 10945
rect 4683 10911 4693 10945
rect 4637 10873 4693 10911
rect 4723 10945 4777 10957
rect 4723 10911 4733 10945
rect 4767 10911 4777 10945
rect 4723 10873 4777 10911
rect 4807 10953 4841 10957
rect 4875 10953 4885 10987
rect 4807 10919 4885 10953
rect 4807 10885 4841 10919
rect 4875 10885 4885 10919
rect 4807 10873 4885 10885
rect 4823 10799 4885 10873
rect 4915 10987 5010 10999
rect 9699 10991 9751 11003
rect 4915 10953 4945 10987
rect 4979 10953 5010 10987
rect 4915 10919 5010 10953
rect 4915 10885 4945 10919
rect 4979 10885 5010 10919
rect 4915 10799 5010 10885
rect 9699 10961 9707 10991
rect 9503 10949 9559 10961
rect 9503 10915 9515 10949
rect 9549 10915 9559 10949
rect 9503 10877 9559 10915
rect 9589 10949 9643 10961
rect 9589 10915 9599 10949
rect 9633 10915 9643 10949
rect 9589 10877 9643 10915
rect 9673 10957 9707 10961
rect 9741 10957 9751 10991
rect 9673 10923 9751 10957
rect 9673 10889 9707 10923
rect 9741 10889 9751 10923
rect 9673 10877 9751 10889
rect 9689 10803 9751 10877
rect 9781 10991 9876 11003
rect 9781 10957 9811 10991
rect 9845 10957 9876 10991
rect 9781 10923 9876 10957
rect 9781 10889 9811 10923
rect 9845 10889 9876 10923
rect 9781 10803 9876 10889
rect 6186 6285 6238 6303
rect 6186 6251 6194 6285
rect 6228 6251 6238 6285
rect 6186 6217 6238 6251
rect 6186 6183 6194 6217
rect 6228 6183 6238 6217
rect 6186 6149 6238 6183
rect 6186 6115 6194 6149
rect 6228 6115 6238 6149
rect 6186 6103 6238 6115
rect 6268 6285 6320 6303
rect 6268 6251 6278 6285
rect 6312 6251 6320 6285
rect 6268 6217 6320 6251
rect 6268 6183 6278 6217
rect 6312 6183 6320 6217
rect 6268 6149 6320 6183
rect 6268 6115 6278 6149
rect 6312 6115 6320 6149
rect 6268 6103 6320 6115
rect 1898 5213 1950 5251
rect 1898 5179 1906 5213
rect 1940 5179 1950 5213
rect 1898 5123 1950 5179
rect 1898 5089 1906 5123
rect 1940 5089 1950 5123
rect 1898 5051 1950 5089
rect 1980 5135 2032 5251
rect 3147 5135 3199 5251
rect 1980 5093 2049 5135
rect 1980 5059 1990 5093
rect 2024 5059 2049 5093
rect 1980 5051 2049 5059
rect 2079 5051 2145 5135
rect 2175 5051 2217 5135
rect 2247 5105 2313 5135
rect 2247 5071 2257 5105
rect 2291 5071 2313 5105
rect 2247 5051 2313 5071
rect 2343 5110 2402 5135
rect 2343 5076 2358 5110
rect 2392 5076 2402 5110
rect 2343 5051 2402 5076
rect 2432 5093 2486 5135
rect 2432 5059 2442 5093
rect 2476 5059 2486 5093
rect 2432 5051 2486 5059
rect 2516 5110 2570 5135
rect 2516 5076 2526 5110
rect 2560 5076 2570 5110
rect 2516 5051 2570 5076
rect 2600 5097 2652 5135
rect 2600 5063 2610 5097
rect 2644 5063 2652 5097
rect 2600 5051 2652 5063
rect 2706 5110 2758 5135
rect 2706 5076 2714 5110
rect 2748 5076 2758 5110
rect 2706 5051 2758 5076
rect 2788 5093 2842 5135
rect 2788 5059 2798 5093
rect 2832 5059 2842 5093
rect 2788 5051 2842 5059
rect 2872 5110 2926 5135
rect 2872 5076 2882 5110
rect 2916 5076 2926 5110
rect 2872 5051 2926 5076
rect 2956 5110 3010 5135
rect 2956 5076 2966 5110
rect 3000 5076 3010 5110
rect 2956 5051 3010 5076
rect 3040 5051 3100 5135
rect 3130 5101 3199 5135
rect 3130 5067 3155 5101
rect 3189 5067 3199 5101
rect 3130 5051 3199 5067
rect 3229 5210 3281 5251
rect 3229 5176 3239 5210
rect 3273 5176 3281 5210
rect 3229 5116 3281 5176
rect 3229 5082 3239 5116
rect 3273 5082 3281 5116
rect 3229 5051 3281 5082
rect 4032 5205 4084 5243
rect 4032 5171 4040 5205
rect 4074 5171 4084 5205
rect 4032 5115 4084 5171
rect 4032 5081 4040 5115
rect 4074 5081 4084 5115
rect 4032 5043 4084 5081
rect 4114 5127 4166 5243
rect 5281 5127 5333 5243
rect 4114 5085 4183 5127
rect 4114 5051 4124 5085
rect 4158 5051 4183 5085
rect 4114 5043 4183 5051
rect 4213 5043 4279 5127
rect 4309 5043 4351 5127
rect 4381 5097 4447 5127
rect 4381 5063 4391 5097
rect 4425 5063 4447 5097
rect 4381 5043 4447 5063
rect 4477 5102 4536 5127
rect 4477 5068 4492 5102
rect 4526 5068 4536 5102
rect 4477 5043 4536 5068
rect 4566 5085 4620 5127
rect 4566 5051 4576 5085
rect 4610 5051 4620 5085
rect 4566 5043 4620 5051
rect 4650 5102 4704 5127
rect 4650 5068 4660 5102
rect 4694 5068 4704 5102
rect 4650 5043 4704 5068
rect 4734 5089 4786 5127
rect 4734 5055 4744 5089
rect 4778 5055 4786 5089
rect 4734 5043 4786 5055
rect 4840 5102 4892 5127
rect 4840 5068 4848 5102
rect 4882 5068 4892 5102
rect 4840 5043 4892 5068
rect 4922 5085 4976 5127
rect 4922 5051 4932 5085
rect 4966 5051 4976 5085
rect 4922 5043 4976 5051
rect 5006 5102 5060 5127
rect 5006 5068 5016 5102
rect 5050 5068 5060 5102
rect 5006 5043 5060 5068
rect 5090 5102 5144 5127
rect 5090 5068 5100 5102
rect 5134 5068 5144 5102
rect 5090 5043 5144 5068
rect 5174 5043 5234 5127
rect 5264 5093 5333 5127
rect 5264 5059 5289 5093
rect 5323 5059 5333 5093
rect 5264 5043 5333 5059
rect 5363 5202 5415 5243
rect 5363 5168 5373 5202
rect 5407 5168 5415 5202
rect 5363 5108 5415 5168
rect 5363 5074 5373 5108
rect 5407 5074 5415 5108
rect 5363 5043 5415 5074
rect 5984 5205 6036 5243
rect 5984 5171 5992 5205
rect 6026 5171 6036 5205
rect 5984 5115 6036 5171
rect 5984 5081 5992 5115
rect 6026 5081 6036 5115
rect 5984 5043 6036 5081
rect 6066 5127 6118 5243
rect 7233 5127 7285 5243
rect 6066 5085 6135 5127
rect 6066 5051 6076 5085
rect 6110 5051 6135 5085
rect 6066 5043 6135 5051
rect 6165 5043 6231 5127
rect 6261 5043 6303 5127
rect 6333 5097 6399 5127
rect 6333 5063 6343 5097
rect 6377 5063 6399 5097
rect 6333 5043 6399 5063
rect 6429 5102 6488 5127
rect 6429 5068 6444 5102
rect 6478 5068 6488 5102
rect 6429 5043 6488 5068
rect 6518 5085 6572 5127
rect 6518 5051 6528 5085
rect 6562 5051 6572 5085
rect 6518 5043 6572 5051
rect 6602 5102 6656 5127
rect 6602 5068 6612 5102
rect 6646 5068 6656 5102
rect 6602 5043 6656 5068
rect 6686 5089 6738 5127
rect 6686 5055 6696 5089
rect 6730 5055 6738 5089
rect 6686 5043 6738 5055
rect 6792 5102 6844 5127
rect 6792 5068 6800 5102
rect 6834 5068 6844 5102
rect 6792 5043 6844 5068
rect 6874 5085 6928 5127
rect 6874 5051 6884 5085
rect 6918 5051 6928 5085
rect 6874 5043 6928 5051
rect 6958 5102 7012 5127
rect 6958 5068 6968 5102
rect 7002 5068 7012 5102
rect 6958 5043 7012 5068
rect 7042 5102 7096 5127
rect 7042 5068 7052 5102
rect 7086 5068 7096 5102
rect 7042 5043 7096 5068
rect 7126 5043 7186 5127
rect 7216 5093 7285 5127
rect 7216 5059 7241 5093
rect 7275 5059 7285 5093
rect 7216 5043 7285 5059
rect 7315 5202 7367 5243
rect 7315 5168 7325 5202
rect 7359 5168 7367 5202
rect 7315 5108 7367 5168
rect 7315 5074 7325 5108
rect 7359 5074 7367 5108
rect 7315 5043 7367 5074
rect 7986 5211 8038 5249
rect 7986 5177 7994 5211
rect 8028 5177 8038 5211
rect 7986 5121 8038 5177
rect 7986 5087 7994 5121
rect 8028 5087 8038 5121
rect 7986 5049 8038 5087
rect 8068 5133 8120 5249
rect 10080 5633 10132 5671
rect 10080 5599 10088 5633
rect 10122 5599 10132 5633
rect 10080 5543 10132 5599
rect 10080 5509 10088 5543
rect 10122 5509 10132 5543
rect 10080 5471 10132 5509
rect 10162 5555 10214 5671
rect 11329 5555 11381 5671
rect 10162 5513 10231 5555
rect 10162 5479 10172 5513
rect 10206 5479 10231 5513
rect 10162 5471 10231 5479
rect 10261 5471 10327 5555
rect 10357 5471 10399 5555
rect 10429 5525 10495 5555
rect 10429 5491 10439 5525
rect 10473 5491 10495 5525
rect 10429 5471 10495 5491
rect 10525 5530 10584 5555
rect 10525 5496 10540 5530
rect 10574 5496 10584 5530
rect 10525 5471 10584 5496
rect 10614 5513 10668 5555
rect 10614 5479 10624 5513
rect 10658 5479 10668 5513
rect 10614 5471 10668 5479
rect 10698 5530 10752 5555
rect 10698 5496 10708 5530
rect 10742 5496 10752 5530
rect 10698 5471 10752 5496
rect 10782 5517 10834 5555
rect 10782 5483 10792 5517
rect 10826 5483 10834 5517
rect 10782 5471 10834 5483
rect 10888 5530 10940 5555
rect 10888 5496 10896 5530
rect 10930 5496 10940 5530
rect 10888 5471 10940 5496
rect 10970 5513 11024 5555
rect 10970 5479 10980 5513
rect 11014 5479 11024 5513
rect 10970 5471 11024 5479
rect 11054 5530 11108 5555
rect 11054 5496 11064 5530
rect 11098 5496 11108 5530
rect 11054 5471 11108 5496
rect 11138 5530 11192 5555
rect 11138 5496 11148 5530
rect 11182 5496 11192 5530
rect 11138 5471 11192 5496
rect 11222 5471 11282 5555
rect 11312 5521 11381 5555
rect 11312 5487 11337 5521
rect 11371 5487 11381 5521
rect 11312 5471 11381 5487
rect 11411 5630 11463 5671
rect 11411 5596 11421 5630
rect 11455 5596 11463 5630
rect 11411 5536 11463 5596
rect 11411 5502 11421 5536
rect 11455 5502 11463 5536
rect 11411 5471 11463 5502
rect 12142 5621 12194 5659
rect 12142 5587 12150 5621
rect 12184 5587 12194 5621
rect 12142 5531 12194 5587
rect 12142 5497 12150 5531
rect 12184 5497 12194 5531
rect 12142 5459 12194 5497
rect 12224 5543 12276 5659
rect 13391 5543 13443 5659
rect 12224 5501 12293 5543
rect 12224 5467 12234 5501
rect 12268 5467 12293 5501
rect 12224 5459 12293 5467
rect 12323 5459 12389 5543
rect 12419 5459 12461 5543
rect 12491 5513 12557 5543
rect 12491 5479 12501 5513
rect 12535 5479 12557 5513
rect 12491 5459 12557 5479
rect 12587 5518 12646 5543
rect 12587 5484 12602 5518
rect 12636 5484 12646 5518
rect 12587 5459 12646 5484
rect 12676 5501 12730 5543
rect 12676 5467 12686 5501
rect 12720 5467 12730 5501
rect 12676 5459 12730 5467
rect 12760 5518 12814 5543
rect 12760 5484 12770 5518
rect 12804 5484 12814 5518
rect 12760 5459 12814 5484
rect 12844 5505 12896 5543
rect 12844 5471 12854 5505
rect 12888 5471 12896 5505
rect 12844 5459 12896 5471
rect 12950 5518 13002 5543
rect 12950 5484 12958 5518
rect 12992 5484 13002 5518
rect 12950 5459 13002 5484
rect 13032 5501 13086 5543
rect 13032 5467 13042 5501
rect 13076 5467 13086 5501
rect 13032 5459 13086 5467
rect 13116 5518 13170 5543
rect 13116 5484 13126 5518
rect 13160 5484 13170 5518
rect 13116 5459 13170 5484
rect 13200 5518 13254 5543
rect 13200 5484 13210 5518
rect 13244 5484 13254 5518
rect 13200 5459 13254 5484
rect 13284 5459 13344 5543
rect 13374 5509 13443 5543
rect 13374 5475 13399 5509
rect 13433 5475 13443 5509
rect 13374 5459 13443 5475
rect 13473 5618 13525 5659
rect 13473 5584 13483 5618
rect 13517 5584 13525 5618
rect 13473 5524 13525 5584
rect 13473 5490 13483 5524
rect 13517 5490 13525 5524
rect 13473 5459 13525 5490
rect 14100 5629 14152 5667
rect 14100 5595 14108 5629
rect 14142 5595 14152 5629
rect 14100 5539 14152 5595
rect 14100 5505 14108 5539
rect 14142 5505 14152 5539
rect 14100 5467 14152 5505
rect 14182 5551 14234 5667
rect 15349 5551 15401 5667
rect 14182 5509 14251 5551
rect 14182 5475 14192 5509
rect 14226 5475 14251 5509
rect 14182 5467 14251 5475
rect 14281 5467 14347 5551
rect 14377 5467 14419 5551
rect 14449 5521 14515 5551
rect 14449 5487 14459 5521
rect 14493 5487 14515 5521
rect 14449 5467 14515 5487
rect 14545 5526 14604 5551
rect 14545 5492 14560 5526
rect 14594 5492 14604 5526
rect 14545 5467 14604 5492
rect 14634 5509 14688 5551
rect 14634 5475 14644 5509
rect 14678 5475 14688 5509
rect 14634 5467 14688 5475
rect 14718 5526 14772 5551
rect 14718 5492 14728 5526
rect 14762 5492 14772 5526
rect 14718 5467 14772 5492
rect 14802 5513 14854 5551
rect 14802 5479 14812 5513
rect 14846 5479 14854 5513
rect 14802 5467 14854 5479
rect 14908 5526 14960 5551
rect 14908 5492 14916 5526
rect 14950 5492 14960 5526
rect 14908 5467 14960 5492
rect 14990 5509 15044 5551
rect 14990 5475 15000 5509
rect 15034 5475 15044 5509
rect 14990 5467 15044 5475
rect 15074 5526 15128 5551
rect 15074 5492 15084 5526
rect 15118 5492 15128 5526
rect 15074 5467 15128 5492
rect 15158 5526 15212 5551
rect 15158 5492 15168 5526
rect 15202 5492 15212 5526
rect 15158 5467 15212 5492
rect 15242 5467 15302 5551
rect 15332 5517 15401 5551
rect 15332 5483 15357 5517
rect 15391 5483 15401 5517
rect 15332 5467 15401 5483
rect 15431 5626 15483 5667
rect 15431 5592 15441 5626
rect 15475 5592 15483 5626
rect 15431 5532 15483 5592
rect 15431 5498 15441 5532
rect 15475 5498 15483 5532
rect 15431 5467 15483 5498
rect 16094 5635 16146 5673
rect 16094 5601 16102 5635
rect 16136 5601 16146 5635
rect 16094 5545 16146 5601
rect 16094 5511 16102 5545
rect 16136 5511 16146 5545
rect 16094 5473 16146 5511
rect 16176 5557 16228 5673
rect 17343 5557 17395 5673
rect 16176 5515 16245 5557
rect 16176 5481 16186 5515
rect 16220 5481 16245 5515
rect 16176 5473 16245 5481
rect 16275 5473 16341 5557
rect 16371 5473 16413 5557
rect 16443 5527 16509 5557
rect 16443 5493 16453 5527
rect 16487 5493 16509 5527
rect 16443 5473 16509 5493
rect 16539 5532 16598 5557
rect 16539 5498 16554 5532
rect 16588 5498 16598 5532
rect 16539 5473 16598 5498
rect 16628 5515 16682 5557
rect 16628 5481 16638 5515
rect 16672 5481 16682 5515
rect 16628 5473 16682 5481
rect 16712 5532 16766 5557
rect 16712 5498 16722 5532
rect 16756 5498 16766 5532
rect 16712 5473 16766 5498
rect 16796 5519 16848 5557
rect 16796 5485 16806 5519
rect 16840 5485 16848 5519
rect 16796 5473 16848 5485
rect 16902 5532 16954 5557
rect 16902 5498 16910 5532
rect 16944 5498 16954 5532
rect 16902 5473 16954 5498
rect 16984 5515 17038 5557
rect 16984 5481 16994 5515
rect 17028 5481 17038 5515
rect 16984 5473 17038 5481
rect 17068 5532 17122 5557
rect 17068 5498 17078 5532
rect 17112 5498 17122 5532
rect 17068 5473 17122 5498
rect 17152 5532 17206 5557
rect 17152 5498 17162 5532
rect 17196 5498 17206 5532
rect 17152 5473 17206 5498
rect 17236 5473 17296 5557
rect 17326 5523 17395 5557
rect 17326 5489 17351 5523
rect 17385 5489 17395 5523
rect 17326 5473 17395 5489
rect 17425 5632 17477 5673
rect 17425 5598 17435 5632
rect 17469 5598 17477 5632
rect 17425 5538 17477 5598
rect 17425 5504 17435 5538
rect 17469 5504 17477 5538
rect 17425 5473 17477 5504
rect 9235 5133 9287 5249
rect 8068 5091 8137 5133
rect 8068 5057 8078 5091
rect 8112 5057 8137 5091
rect 8068 5049 8137 5057
rect 8167 5049 8233 5133
rect 8263 5049 8305 5133
rect 8335 5103 8401 5133
rect 8335 5069 8345 5103
rect 8379 5069 8401 5103
rect 8335 5049 8401 5069
rect 8431 5108 8490 5133
rect 8431 5074 8446 5108
rect 8480 5074 8490 5108
rect 8431 5049 8490 5074
rect 8520 5091 8574 5133
rect 8520 5057 8530 5091
rect 8564 5057 8574 5091
rect 8520 5049 8574 5057
rect 8604 5108 8658 5133
rect 8604 5074 8614 5108
rect 8648 5074 8658 5108
rect 8604 5049 8658 5074
rect 8688 5095 8740 5133
rect 8688 5061 8698 5095
rect 8732 5061 8740 5095
rect 8688 5049 8740 5061
rect 8794 5108 8846 5133
rect 8794 5074 8802 5108
rect 8836 5074 8846 5108
rect 8794 5049 8846 5074
rect 8876 5091 8930 5133
rect 8876 5057 8886 5091
rect 8920 5057 8930 5091
rect 8876 5049 8930 5057
rect 8960 5108 9014 5133
rect 8960 5074 8970 5108
rect 9004 5074 9014 5108
rect 8960 5049 9014 5074
rect 9044 5108 9098 5133
rect 9044 5074 9054 5108
rect 9088 5074 9098 5108
rect 9044 5049 9098 5074
rect 9128 5049 9188 5133
rect 9218 5099 9287 5133
rect 9218 5065 9243 5099
rect 9277 5065 9287 5099
rect 9218 5049 9287 5065
rect 9317 5208 9369 5249
rect 9317 5174 9327 5208
rect 9361 5174 9369 5208
rect 9317 5114 9369 5174
rect 9317 5080 9327 5114
rect 9361 5080 9369 5114
rect 9317 5049 9369 5080
rect 10108 4759 10160 4797
rect 10108 4725 10116 4759
rect 10150 4725 10160 4759
rect 10108 4669 10160 4725
rect 10108 4635 10116 4669
rect 10150 4635 10160 4669
rect 10108 4597 10160 4635
rect 10190 4681 10242 4797
rect 11357 4681 11409 4797
rect 10190 4639 10259 4681
rect 10190 4605 10200 4639
rect 10234 4605 10259 4639
rect 10190 4597 10259 4605
rect 10289 4597 10355 4681
rect 10385 4597 10427 4681
rect 10457 4651 10523 4681
rect 10457 4617 10467 4651
rect 10501 4617 10523 4651
rect 10457 4597 10523 4617
rect 10553 4656 10612 4681
rect 10553 4622 10568 4656
rect 10602 4622 10612 4656
rect 10553 4597 10612 4622
rect 10642 4639 10696 4681
rect 10642 4605 10652 4639
rect 10686 4605 10696 4639
rect 10642 4597 10696 4605
rect 10726 4656 10780 4681
rect 10726 4622 10736 4656
rect 10770 4622 10780 4656
rect 10726 4597 10780 4622
rect 10810 4643 10862 4681
rect 10810 4609 10820 4643
rect 10854 4609 10862 4643
rect 10810 4597 10862 4609
rect 10916 4656 10968 4681
rect 10916 4622 10924 4656
rect 10958 4622 10968 4656
rect 10916 4597 10968 4622
rect 10998 4639 11052 4681
rect 10998 4605 11008 4639
rect 11042 4605 11052 4639
rect 10998 4597 11052 4605
rect 11082 4656 11136 4681
rect 11082 4622 11092 4656
rect 11126 4622 11136 4656
rect 11082 4597 11136 4622
rect 11166 4656 11220 4681
rect 11166 4622 11176 4656
rect 11210 4622 11220 4656
rect 11166 4597 11220 4622
rect 11250 4597 11310 4681
rect 11340 4647 11409 4681
rect 11340 4613 11365 4647
rect 11399 4613 11409 4647
rect 11340 4597 11409 4613
rect 11439 4756 11491 4797
rect 11439 4722 11449 4756
rect 11483 4722 11491 4756
rect 11439 4662 11491 4722
rect 11439 4628 11449 4662
rect 11483 4628 11491 4662
rect 11439 4597 11491 4628
rect 12378 4715 12430 4753
rect 12378 4681 12386 4715
rect 12420 4681 12430 4715
rect 12378 4625 12430 4681
rect 12378 4591 12386 4625
rect 12420 4591 12430 4625
rect 12378 4553 12430 4591
rect 12460 4637 12512 4753
rect 18969 5081 19021 5099
rect 18969 5047 18977 5081
rect 19011 5047 19021 5081
rect 18969 5022 19021 5047
rect 18371 5005 18427 5022
rect 13627 4637 13679 4753
rect 12460 4595 12529 4637
rect 12460 4561 12470 4595
rect 12504 4561 12529 4595
rect 12460 4553 12529 4561
rect 12559 4553 12625 4637
rect 12655 4553 12697 4637
rect 12727 4607 12793 4637
rect 12727 4573 12737 4607
rect 12771 4573 12793 4607
rect 12727 4553 12793 4573
rect 12823 4612 12882 4637
rect 12823 4578 12838 4612
rect 12872 4578 12882 4612
rect 12823 4553 12882 4578
rect 12912 4595 12966 4637
rect 12912 4561 12922 4595
rect 12956 4561 12966 4595
rect 12912 4553 12966 4561
rect 12996 4612 13050 4637
rect 12996 4578 13006 4612
rect 13040 4578 13050 4612
rect 12996 4553 13050 4578
rect 13080 4599 13132 4637
rect 13080 4565 13090 4599
rect 13124 4565 13132 4599
rect 13080 4553 13132 4565
rect 13186 4612 13238 4637
rect 13186 4578 13194 4612
rect 13228 4578 13238 4612
rect 13186 4553 13238 4578
rect 13268 4595 13322 4637
rect 13268 4561 13278 4595
rect 13312 4561 13322 4595
rect 13268 4553 13322 4561
rect 13352 4612 13406 4637
rect 13352 4578 13362 4612
rect 13396 4578 13406 4612
rect 13352 4553 13406 4578
rect 13436 4612 13490 4637
rect 13436 4578 13446 4612
rect 13480 4578 13490 4612
rect 13436 4553 13490 4578
rect 13520 4553 13580 4637
rect 13610 4603 13679 4637
rect 13610 4569 13635 4603
rect 13669 4569 13679 4603
rect 13610 4553 13679 4569
rect 13709 4712 13761 4753
rect 13709 4678 13719 4712
rect 13753 4678 13761 4712
rect 13709 4618 13761 4678
rect 13709 4584 13719 4618
rect 13753 4584 13761 4618
rect 13709 4553 13761 4584
rect 14380 4709 14432 4747
rect 14380 4675 14388 4709
rect 14422 4675 14432 4709
rect 14380 4619 14432 4675
rect 14380 4585 14388 4619
rect 14422 4585 14432 4619
rect 14380 4547 14432 4585
rect 14462 4631 14514 4747
rect 15629 4631 15681 4747
rect 14462 4589 14531 4631
rect 14462 4555 14472 4589
rect 14506 4555 14531 4589
rect 14462 4547 14531 4555
rect 14561 4547 14627 4631
rect 14657 4547 14699 4631
rect 14729 4601 14795 4631
rect 14729 4567 14739 4601
rect 14773 4567 14795 4601
rect 14729 4547 14795 4567
rect 14825 4606 14884 4631
rect 14825 4572 14840 4606
rect 14874 4572 14884 4606
rect 14825 4547 14884 4572
rect 14914 4589 14968 4631
rect 14914 4555 14924 4589
rect 14958 4555 14968 4589
rect 14914 4547 14968 4555
rect 14998 4606 15052 4631
rect 14998 4572 15008 4606
rect 15042 4572 15052 4606
rect 14998 4547 15052 4572
rect 15082 4593 15134 4631
rect 15082 4559 15092 4593
rect 15126 4559 15134 4593
rect 15082 4547 15134 4559
rect 15188 4606 15240 4631
rect 15188 4572 15196 4606
rect 15230 4572 15240 4606
rect 15188 4547 15240 4572
rect 15270 4589 15324 4631
rect 15270 4555 15280 4589
rect 15314 4555 15324 4589
rect 15270 4547 15324 4555
rect 15354 4606 15408 4631
rect 15354 4572 15364 4606
rect 15398 4572 15408 4606
rect 15354 4547 15408 4572
rect 15438 4606 15492 4631
rect 15438 4572 15448 4606
rect 15482 4572 15492 4606
rect 15438 4547 15492 4572
rect 15522 4547 15582 4631
rect 15612 4597 15681 4631
rect 15612 4563 15637 4597
rect 15671 4563 15681 4597
rect 15612 4547 15681 4563
rect 15711 4706 15763 4747
rect 15711 4672 15721 4706
rect 15755 4672 15763 4706
rect 15711 4612 15763 4672
rect 15711 4578 15721 4612
rect 15755 4578 15763 4612
rect 15711 4547 15763 4578
rect 16402 4691 16454 4729
rect 16402 4657 16410 4691
rect 16444 4657 16454 4691
rect 16402 4601 16454 4657
rect 16402 4567 16410 4601
rect 16444 4567 16454 4601
rect 16402 4529 16454 4567
rect 16484 4613 16536 4729
rect 18371 4971 18383 5005
rect 18417 4971 18427 5005
rect 18371 4938 18427 4971
rect 18457 5005 18523 5022
rect 18457 4971 18469 5005
rect 18503 4971 18523 5005
rect 18457 4938 18523 4971
rect 18553 4938 18595 5022
rect 18625 5005 18809 5022
rect 18625 4971 18666 5005
rect 18700 4971 18741 5005
rect 18775 4971 18809 5005
rect 18625 4938 18809 4971
rect 18839 4938 18912 5022
rect 18942 5013 19021 5022
rect 18942 4979 18977 5013
rect 19011 4979 19021 5013
rect 18942 4945 19021 4979
rect 18942 4938 18977 4945
rect 18969 4911 18977 4938
rect 19011 4911 19021 4945
rect 18969 4899 19021 4911
rect 19051 5081 19103 5099
rect 19051 5047 19061 5081
rect 19095 5047 19103 5081
rect 19051 5013 19103 5047
rect 19051 4979 19061 5013
rect 19095 4979 19103 5013
rect 19051 4945 19103 4979
rect 19051 4911 19061 4945
rect 19095 4911 19103 4945
rect 19051 4899 19103 4911
rect 17651 4613 17703 4729
rect 16484 4571 16553 4613
rect 16484 4537 16494 4571
rect 16528 4537 16553 4571
rect 16484 4529 16553 4537
rect 16583 4529 16649 4613
rect 16679 4529 16721 4613
rect 16751 4583 16817 4613
rect 16751 4549 16761 4583
rect 16795 4549 16817 4583
rect 16751 4529 16817 4549
rect 16847 4588 16906 4613
rect 16847 4554 16862 4588
rect 16896 4554 16906 4588
rect 16847 4529 16906 4554
rect 16936 4571 16990 4613
rect 16936 4537 16946 4571
rect 16980 4537 16990 4571
rect 16936 4529 16990 4537
rect 17020 4588 17074 4613
rect 17020 4554 17030 4588
rect 17064 4554 17074 4588
rect 17020 4529 17074 4554
rect 17104 4575 17156 4613
rect 17104 4541 17114 4575
rect 17148 4541 17156 4575
rect 17104 4529 17156 4541
rect 17210 4588 17262 4613
rect 17210 4554 17218 4588
rect 17252 4554 17262 4588
rect 17210 4529 17262 4554
rect 17292 4571 17346 4613
rect 17292 4537 17302 4571
rect 17336 4537 17346 4571
rect 17292 4529 17346 4537
rect 17376 4588 17430 4613
rect 17376 4554 17386 4588
rect 17420 4554 17430 4588
rect 17376 4529 17430 4554
rect 17460 4588 17514 4613
rect 17460 4554 17470 4588
rect 17504 4554 17514 4588
rect 17460 4529 17514 4554
rect 17544 4529 17604 4613
rect 17634 4579 17703 4613
rect 17634 4545 17659 4579
rect 17693 4545 17703 4579
rect 17634 4529 17703 4545
rect 17733 4688 17785 4729
rect 17733 4654 17743 4688
rect 17777 4654 17785 4688
rect 17733 4594 17785 4654
rect 17733 4560 17743 4594
rect 17777 4560 17785 4594
rect 17733 4529 17785 4560
rect 6156 3025 6208 3043
rect 6156 2991 6164 3025
rect 6198 2991 6208 3025
rect 6156 2957 6208 2991
rect 6156 2923 6164 2957
rect 6198 2923 6208 2957
rect 6156 2889 6208 2923
rect 6156 2855 6164 2889
rect 6198 2855 6208 2889
rect 6156 2843 6208 2855
rect 6238 3025 6290 3043
rect 6238 2991 6248 3025
rect 6282 2991 6290 3025
rect 6238 2957 6290 2991
rect 6238 2923 6248 2957
rect 6282 2923 6290 2957
rect 6238 2889 6290 2923
rect 6238 2855 6248 2889
rect 6282 2855 6290 2889
rect 6238 2843 6290 2855
rect 1868 1953 1920 1991
rect 1868 1919 1876 1953
rect 1910 1919 1920 1953
rect 1868 1863 1920 1919
rect 1868 1829 1876 1863
rect 1910 1829 1920 1863
rect 1868 1791 1920 1829
rect 1950 1875 2002 1991
rect 3117 1875 3169 1991
rect 1950 1833 2019 1875
rect 1950 1799 1960 1833
rect 1994 1799 2019 1833
rect 1950 1791 2019 1799
rect 2049 1791 2115 1875
rect 2145 1791 2187 1875
rect 2217 1845 2283 1875
rect 2217 1811 2227 1845
rect 2261 1811 2283 1845
rect 2217 1791 2283 1811
rect 2313 1850 2372 1875
rect 2313 1816 2328 1850
rect 2362 1816 2372 1850
rect 2313 1791 2372 1816
rect 2402 1833 2456 1875
rect 2402 1799 2412 1833
rect 2446 1799 2456 1833
rect 2402 1791 2456 1799
rect 2486 1850 2540 1875
rect 2486 1816 2496 1850
rect 2530 1816 2540 1850
rect 2486 1791 2540 1816
rect 2570 1837 2622 1875
rect 2570 1803 2580 1837
rect 2614 1803 2622 1837
rect 2570 1791 2622 1803
rect 2676 1850 2728 1875
rect 2676 1816 2684 1850
rect 2718 1816 2728 1850
rect 2676 1791 2728 1816
rect 2758 1833 2812 1875
rect 2758 1799 2768 1833
rect 2802 1799 2812 1833
rect 2758 1791 2812 1799
rect 2842 1850 2896 1875
rect 2842 1816 2852 1850
rect 2886 1816 2896 1850
rect 2842 1791 2896 1816
rect 2926 1850 2980 1875
rect 2926 1816 2936 1850
rect 2970 1816 2980 1850
rect 2926 1791 2980 1816
rect 3010 1791 3070 1875
rect 3100 1841 3169 1875
rect 3100 1807 3125 1841
rect 3159 1807 3169 1841
rect 3100 1791 3169 1807
rect 3199 1950 3251 1991
rect 3199 1916 3209 1950
rect 3243 1916 3251 1950
rect 3199 1856 3251 1916
rect 3199 1822 3209 1856
rect 3243 1822 3251 1856
rect 3199 1791 3251 1822
rect 3938 1949 3990 1987
rect 3938 1915 3946 1949
rect 3980 1915 3990 1949
rect 3938 1859 3990 1915
rect 3938 1825 3946 1859
rect 3980 1825 3990 1859
rect 3938 1787 3990 1825
rect 4020 1871 4072 1987
rect 5187 1871 5239 1987
rect 4020 1829 4089 1871
rect 4020 1795 4030 1829
rect 4064 1795 4089 1829
rect 4020 1787 4089 1795
rect 4119 1787 4185 1871
rect 4215 1787 4257 1871
rect 4287 1841 4353 1871
rect 4287 1807 4297 1841
rect 4331 1807 4353 1841
rect 4287 1787 4353 1807
rect 4383 1846 4442 1871
rect 4383 1812 4398 1846
rect 4432 1812 4442 1846
rect 4383 1787 4442 1812
rect 4472 1829 4526 1871
rect 4472 1795 4482 1829
rect 4516 1795 4526 1829
rect 4472 1787 4526 1795
rect 4556 1846 4610 1871
rect 4556 1812 4566 1846
rect 4600 1812 4610 1846
rect 4556 1787 4610 1812
rect 4640 1833 4692 1871
rect 4640 1799 4650 1833
rect 4684 1799 4692 1833
rect 4640 1787 4692 1799
rect 4746 1846 4798 1871
rect 4746 1812 4754 1846
rect 4788 1812 4798 1846
rect 4746 1787 4798 1812
rect 4828 1829 4882 1871
rect 4828 1795 4838 1829
rect 4872 1795 4882 1829
rect 4828 1787 4882 1795
rect 4912 1846 4966 1871
rect 4912 1812 4922 1846
rect 4956 1812 4966 1846
rect 4912 1787 4966 1812
rect 4996 1846 5050 1871
rect 4996 1812 5006 1846
rect 5040 1812 5050 1846
rect 4996 1787 5050 1812
rect 5080 1787 5140 1871
rect 5170 1837 5239 1871
rect 5170 1803 5195 1837
rect 5229 1803 5239 1837
rect 5170 1787 5239 1803
rect 5269 1946 5321 1987
rect 5269 1912 5279 1946
rect 5313 1912 5321 1946
rect 5269 1852 5321 1912
rect 5269 1818 5279 1852
rect 5313 1818 5321 1852
rect 5269 1787 5321 1818
rect 5890 1949 5942 1987
rect 5890 1915 5898 1949
rect 5932 1915 5942 1949
rect 5890 1859 5942 1915
rect 5890 1825 5898 1859
rect 5932 1825 5942 1859
rect 5890 1787 5942 1825
rect 5972 1871 6024 1987
rect 7139 1871 7191 1987
rect 5972 1829 6041 1871
rect 5972 1795 5982 1829
rect 6016 1795 6041 1829
rect 5972 1787 6041 1795
rect 6071 1787 6137 1871
rect 6167 1787 6209 1871
rect 6239 1841 6305 1871
rect 6239 1807 6249 1841
rect 6283 1807 6305 1841
rect 6239 1787 6305 1807
rect 6335 1846 6394 1871
rect 6335 1812 6350 1846
rect 6384 1812 6394 1846
rect 6335 1787 6394 1812
rect 6424 1829 6478 1871
rect 6424 1795 6434 1829
rect 6468 1795 6478 1829
rect 6424 1787 6478 1795
rect 6508 1846 6562 1871
rect 6508 1812 6518 1846
rect 6552 1812 6562 1846
rect 6508 1787 6562 1812
rect 6592 1833 6644 1871
rect 6592 1799 6602 1833
rect 6636 1799 6644 1833
rect 6592 1787 6644 1799
rect 6698 1846 6750 1871
rect 6698 1812 6706 1846
rect 6740 1812 6750 1846
rect 6698 1787 6750 1812
rect 6780 1829 6834 1871
rect 6780 1795 6790 1829
rect 6824 1795 6834 1829
rect 6780 1787 6834 1795
rect 6864 1846 6918 1871
rect 6864 1812 6874 1846
rect 6908 1812 6918 1846
rect 6864 1787 6918 1812
rect 6948 1846 7002 1871
rect 6948 1812 6958 1846
rect 6992 1812 7002 1846
rect 6948 1787 7002 1812
rect 7032 1787 7092 1871
rect 7122 1837 7191 1871
rect 7122 1803 7147 1837
rect 7181 1803 7191 1837
rect 7122 1787 7191 1803
rect 7221 1946 7273 1987
rect 7221 1912 7231 1946
rect 7265 1912 7273 1946
rect 7221 1852 7273 1912
rect 7221 1818 7231 1852
rect 7265 1818 7273 1852
rect 7221 1787 7273 1818
rect 7892 1955 7944 1993
rect 7892 1921 7900 1955
rect 7934 1921 7944 1955
rect 7892 1865 7944 1921
rect 7892 1831 7900 1865
rect 7934 1831 7944 1865
rect 7892 1793 7944 1831
rect 7974 1877 8026 1993
rect 9141 1877 9193 1993
rect 7974 1835 8043 1877
rect 7974 1801 7984 1835
rect 8018 1801 8043 1835
rect 7974 1793 8043 1801
rect 8073 1793 8139 1877
rect 8169 1793 8211 1877
rect 8241 1847 8307 1877
rect 8241 1813 8251 1847
rect 8285 1813 8307 1847
rect 8241 1793 8307 1813
rect 8337 1852 8396 1877
rect 8337 1818 8352 1852
rect 8386 1818 8396 1852
rect 8337 1793 8396 1818
rect 8426 1835 8480 1877
rect 8426 1801 8436 1835
rect 8470 1801 8480 1835
rect 8426 1793 8480 1801
rect 8510 1852 8564 1877
rect 8510 1818 8520 1852
rect 8554 1818 8564 1852
rect 8510 1793 8564 1818
rect 8594 1839 8646 1877
rect 8594 1805 8604 1839
rect 8638 1805 8646 1839
rect 8594 1793 8646 1805
rect 8700 1852 8752 1877
rect 8700 1818 8708 1852
rect 8742 1818 8752 1852
rect 8700 1793 8752 1818
rect 8782 1835 8836 1877
rect 8782 1801 8792 1835
rect 8826 1801 8836 1835
rect 8782 1793 8836 1801
rect 8866 1852 8920 1877
rect 8866 1818 8876 1852
rect 8910 1818 8920 1852
rect 8866 1793 8920 1818
rect 8950 1852 9004 1877
rect 8950 1818 8960 1852
rect 8994 1818 9004 1852
rect 8950 1793 9004 1818
rect 9034 1793 9094 1877
rect 9124 1843 9193 1877
rect 9124 1809 9149 1843
rect 9183 1809 9193 1843
rect 9124 1793 9193 1809
rect 9223 1952 9275 1993
rect 9223 1918 9233 1952
rect 9267 1918 9275 1952
rect 9223 1858 9275 1918
rect 9223 1824 9233 1858
rect 9267 1824 9275 1858
rect 9223 1793 9275 1824
rect 9844 1955 9896 1993
rect 9844 1921 9852 1955
rect 9886 1921 9896 1955
rect 9844 1865 9896 1921
rect 9844 1831 9852 1865
rect 9886 1831 9896 1865
rect 9844 1793 9896 1831
rect 9926 1877 9978 1993
rect 11093 1877 11145 1993
rect 9926 1835 9995 1877
rect 9926 1801 9936 1835
rect 9970 1801 9995 1835
rect 9926 1793 9995 1801
rect 10025 1793 10091 1877
rect 10121 1793 10163 1877
rect 10193 1847 10259 1877
rect 10193 1813 10203 1847
rect 10237 1813 10259 1847
rect 10193 1793 10259 1813
rect 10289 1852 10348 1877
rect 10289 1818 10304 1852
rect 10338 1818 10348 1852
rect 10289 1793 10348 1818
rect 10378 1835 10432 1877
rect 10378 1801 10388 1835
rect 10422 1801 10432 1835
rect 10378 1793 10432 1801
rect 10462 1852 10516 1877
rect 10462 1818 10472 1852
rect 10506 1818 10516 1852
rect 10462 1793 10516 1818
rect 10546 1839 10598 1877
rect 10546 1805 10556 1839
rect 10590 1805 10598 1839
rect 10546 1793 10598 1805
rect 10652 1852 10704 1877
rect 10652 1818 10660 1852
rect 10694 1818 10704 1852
rect 10652 1793 10704 1818
rect 10734 1835 10788 1877
rect 10734 1801 10744 1835
rect 10778 1801 10788 1835
rect 10734 1793 10788 1801
rect 10818 1852 10872 1877
rect 10818 1818 10828 1852
rect 10862 1818 10872 1852
rect 10818 1793 10872 1818
rect 10902 1852 10956 1877
rect 10902 1818 10912 1852
rect 10946 1818 10956 1852
rect 10902 1793 10956 1818
rect 10986 1793 11046 1877
rect 11076 1843 11145 1877
rect 11076 1809 11101 1843
rect 11135 1809 11145 1843
rect 11076 1793 11145 1809
rect 11175 1952 11227 1993
rect 11175 1918 11185 1952
rect 11219 1918 11227 1952
rect 11175 1858 11227 1918
rect 11175 1824 11185 1858
rect 11219 1824 11227 1858
rect 11175 1793 11227 1824
rect 11836 1955 11888 1993
rect 11836 1921 11844 1955
rect 11878 1921 11888 1955
rect 11836 1865 11888 1921
rect 11836 1831 11844 1865
rect 11878 1831 11888 1865
rect 11836 1793 11888 1831
rect 11918 1877 11970 1993
rect 13085 1877 13137 1993
rect 11918 1835 11987 1877
rect 11918 1801 11928 1835
rect 11962 1801 11987 1835
rect 11918 1793 11987 1801
rect 12017 1793 12083 1877
rect 12113 1793 12155 1877
rect 12185 1847 12251 1877
rect 12185 1813 12195 1847
rect 12229 1813 12251 1847
rect 12185 1793 12251 1813
rect 12281 1852 12340 1877
rect 12281 1818 12296 1852
rect 12330 1818 12340 1852
rect 12281 1793 12340 1818
rect 12370 1835 12424 1877
rect 12370 1801 12380 1835
rect 12414 1801 12424 1835
rect 12370 1793 12424 1801
rect 12454 1852 12508 1877
rect 12454 1818 12464 1852
rect 12498 1818 12508 1852
rect 12454 1793 12508 1818
rect 12538 1839 12590 1877
rect 12538 1805 12548 1839
rect 12582 1805 12590 1839
rect 12538 1793 12590 1805
rect 12644 1852 12696 1877
rect 12644 1818 12652 1852
rect 12686 1818 12696 1852
rect 12644 1793 12696 1818
rect 12726 1835 12780 1877
rect 12726 1801 12736 1835
rect 12770 1801 12780 1835
rect 12726 1793 12780 1801
rect 12810 1852 12864 1877
rect 12810 1818 12820 1852
rect 12854 1818 12864 1852
rect 12810 1793 12864 1818
rect 12894 1852 12948 1877
rect 12894 1818 12904 1852
rect 12938 1818 12948 1852
rect 12894 1793 12948 1818
rect 12978 1793 13038 1877
rect 13068 1843 13137 1877
rect 13068 1809 13093 1843
rect 13127 1809 13137 1843
rect 13068 1793 13137 1809
rect 13167 1952 13219 1993
rect 13167 1918 13177 1952
rect 13211 1918 13219 1952
rect 13167 1858 13219 1918
rect 13167 1824 13177 1858
rect 13211 1824 13219 1858
rect 13167 1793 13219 1824
rect 13788 1955 13840 1993
rect 13788 1921 13796 1955
rect 13830 1921 13840 1955
rect 13788 1865 13840 1921
rect 13788 1831 13796 1865
rect 13830 1831 13840 1865
rect 13788 1793 13840 1831
rect 13870 1877 13922 1993
rect 15037 1877 15089 1993
rect 13870 1835 13939 1877
rect 13870 1801 13880 1835
rect 13914 1801 13939 1835
rect 13870 1793 13939 1801
rect 13969 1793 14035 1877
rect 14065 1793 14107 1877
rect 14137 1847 14203 1877
rect 14137 1813 14147 1847
rect 14181 1813 14203 1847
rect 14137 1793 14203 1813
rect 14233 1852 14292 1877
rect 14233 1818 14248 1852
rect 14282 1818 14292 1852
rect 14233 1793 14292 1818
rect 14322 1835 14376 1877
rect 14322 1801 14332 1835
rect 14366 1801 14376 1835
rect 14322 1793 14376 1801
rect 14406 1852 14460 1877
rect 14406 1818 14416 1852
rect 14450 1818 14460 1852
rect 14406 1793 14460 1818
rect 14490 1839 14542 1877
rect 14490 1805 14500 1839
rect 14534 1805 14542 1839
rect 14490 1793 14542 1805
rect 14596 1852 14648 1877
rect 14596 1818 14604 1852
rect 14638 1818 14648 1852
rect 14596 1793 14648 1818
rect 14678 1835 14732 1877
rect 14678 1801 14688 1835
rect 14722 1801 14732 1835
rect 14678 1793 14732 1801
rect 14762 1852 14816 1877
rect 14762 1818 14772 1852
rect 14806 1818 14816 1852
rect 14762 1793 14816 1818
rect 14846 1852 14900 1877
rect 14846 1818 14856 1852
rect 14890 1818 14900 1852
rect 14846 1793 14900 1818
rect 14930 1793 14990 1877
rect 15020 1843 15089 1877
rect 15020 1809 15045 1843
rect 15079 1809 15089 1843
rect 15020 1793 15089 1809
rect 15119 1952 15171 1993
rect 15119 1918 15129 1952
rect 15163 1918 15171 1952
rect 15119 1858 15171 1918
rect 15119 1824 15129 1858
rect 15163 1824 15171 1858
rect 15119 1793 15171 1824
rect 15852 1955 15904 1993
rect 15852 1921 15860 1955
rect 15894 1921 15904 1955
rect 15852 1865 15904 1921
rect 15852 1831 15860 1865
rect 15894 1831 15904 1865
rect 15852 1793 15904 1831
rect 15934 1877 15986 1993
rect 17101 1877 17153 1993
rect 15934 1835 16003 1877
rect 15934 1801 15944 1835
rect 15978 1801 16003 1835
rect 15934 1793 16003 1801
rect 16033 1793 16099 1877
rect 16129 1793 16171 1877
rect 16201 1847 16267 1877
rect 16201 1813 16211 1847
rect 16245 1813 16267 1847
rect 16201 1793 16267 1813
rect 16297 1852 16356 1877
rect 16297 1818 16312 1852
rect 16346 1818 16356 1852
rect 16297 1793 16356 1818
rect 16386 1835 16440 1877
rect 16386 1801 16396 1835
rect 16430 1801 16440 1835
rect 16386 1793 16440 1801
rect 16470 1852 16524 1877
rect 16470 1818 16480 1852
rect 16514 1818 16524 1852
rect 16470 1793 16524 1818
rect 16554 1839 16606 1877
rect 16554 1805 16564 1839
rect 16598 1805 16606 1839
rect 16554 1793 16606 1805
rect 16660 1852 16712 1877
rect 16660 1818 16668 1852
rect 16702 1818 16712 1852
rect 16660 1793 16712 1818
rect 16742 1835 16796 1877
rect 16742 1801 16752 1835
rect 16786 1801 16796 1835
rect 16742 1793 16796 1801
rect 16826 1852 16880 1877
rect 16826 1818 16836 1852
rect 16870 1818 16880 1852
rect 16826 1793 16880 1818
rect 16910 1852 16964 1877
rect 16910 1818 16920 1852
rect 16954 1818 16964 1852
rect 16910 1793 16964 1818
rect 16994 1793 17054 1877
rect 17084 1843 17153 1877
rect 17084 1809 17109 1843
rect 17143 1809 17153 1843
rect 17084 1793 17153 1809
rect 17183 1952 17235 1993
rect 17183 1918 17193 1952
rect 17227 1918 17235 1952
rect 17183 1858 17235 1918
rect 17183 1824 17193 1858
rect 17227 1824 17235 1858
rect 17183 1793 17235 1824
<< ndiffc >>
rect 18979 43340 19013 43374
rect 19047 43340 19081 43374
rect 18979 43256 19013 43290
rect 19047 43256 19081 43290
rect 19047 43172 19081 43206
rect 18979 43088 19013 43122
rect 19047 43088 19081 43122
rect 19047 43004 19081 43038
rect 18979 42920 19013 42954
rect 19047 42920 19081 42954
rect 19047 42836 19081 42870
rect 18979 42752 19013 42786
rect 19047 42752 19081 42786
rect 19047 42668 19081 42702
rect 18979 42584 19013 42618
rect 19047 42584 19081 42618
rect 19047 42500 19081 42534
rect 18979 42416 19013 42450
rect 19047 42416 19081 42450
rect 19047 42332 19081 42366
rect 18979 42248 19013 42282
rect 19047 42248 19081 42282
rect 19047 42164 19081 42198
rect 18979 42080 19013 42114
rect 19047 42080 19081 42114
rect 18979 41996 19013 42030
rect 19047 41996 19081 42030
rect 19031 41363 19065 41397
rect 18963 41228 18997 41262
rect 19031 41228 19065 41262
rect 19031 41144 19065 41178
rect 18963 41060 18997 41094
rect 19031 41060 19065 41094
rect 19031 40976 19065 41010
rect 18963 40892 18997 40926
rect 19031 40892 19065 40926
rect 19031 40808 19065 40842
rect 18963 40724 18997 40758
rect 19031 40724 19065 40758
rect 19031 40640 19065 40674
rect 18963 40556 18997 40590
rect 19031 40556 19065 40590
rect 19031 40472 19065 40506
rect 18963 40388 18997 40422
rect 19031 40388 19065 40422
rect 19031 40304 19065 40338
rect 19039 39548 19073 39582
rect 18971 39464 19005 39498
rect 19039 39464 19073 39498
rect 19039 39380 19073 39414
rect 18971 39296 19005 39330
rect 19039 39296 19073 39330
rect 19039 39212 19073 39246
rect 18971 39128 19005 39162
rect 19039 39128 19073 39162
rect 19039 39044 19073 39078
rect 18971 38960 19005 38994
rect 19039 38960 19073 38994
rect 19039 38876 19073 38910
rect 19052 38303 19086 38337
rect 19045 38219 19079 38253
rect 19053 38135 19087 38169
rect 19045 38051 19079 38085
rect 19053 37967 19087 38001
rect 19045 37883 19079 37917
rect 19053 37775 19087 37809
rect 19064 37145 19098 37179
rect 19057 37061 19091 37095
rect 19065 36977 19099 37011
rect 19057 36893 19091 36927
rect 19065 36809 19099 36843
rect 19001 36265 19035 36299
rect 19073 36265 19107 36299
rect 19001 36181 19035 36215
rect 19073 36181 19107 36215
rect 19001 36097 19035 36131
rect 19073 36097 19107 36131
rect 19059 34879 19093 34913
rect 19097 34795 19131 34829
rect 19071 34700 19105 34734
rect 19026 34596 19060 34630
rect 19094 34596 19128 34630
rect 19067 34512 19101 34546
rect 19028 34428 19062 34462
rect 19096 34428 19130 34462
rect 19083 34322 19117 34356
rect 19083 34124 19117 34158
rect 19083 34021 19117 34055
rect 19089 33902 19123 33936
rect 19083 33703 19117 33737
rect 19083 33592 19117 33626
rect 19097 33507 19131 33541
rect 19071 33403 19105 33437
rect 19097 33319 19131 33353
rect 19071 33235 19105 33269
rect 19059 32597 19093 32631
rect 19097 32513 19131 32547
rect 19071 32418 19105 32452
rect 19026 32314 19060 32348
rect 19094 32314 19128 32348
rect 19067 32230 19101 32264
rect 19028 32146 19062 32180
rect 19096 32146 19130 32180
rect 19083 32040 19117 32074
rect 19083 31842 19117 31876
rect 19083 31739 19117 31773
rect 19089 31620 19123 31654
rect 19083 31421 19117 31455
rect 19083 31310 19117 31344
rect 19097 31225 19131 31259
rect 19071 31121 19105 31155
rect 19097 31037 19131 31071
rect 19071 30953 19105 30987
rect 19063 30351 19097 30385
rect 19101 30267 19135 30301
rect 19075 30172 19109 30206
rect 19030 30068 19064 30102
rect 19098 30068 19132 30102
rect 19071 29984 19105 30018
rect 19032 29900 19066 29934
rect 19100 29900 19134 29934
rect 19087 29794 19121 29828
rect 19087 29596 19121 29630
rect 19087 29493 19121 29527
rect 19093 29374 19127 29408
rect 19087 29175 19121 29209
rect 19087 29064 19121 29098
rect 19101 28979 19135 29013
rect 19075 28875 19109 28909
rect 19101 28791 19135 28825
rect 19075 28707 19109 28741
rect 19055 28165 19089 28199
rect 19093 28081 19127 28115
rect 19067 27986 19101 28020
rect 19022 27882 19056 27916
rect 19090 27882 19124 27916
rect 19063 27798 19097 27832
rect 19024 27714 19058 27748
rect 19092 27714 19126 27748
rect 19079 27608 19113 27642
rect 19079 27410 19113 27444
rect 19079 27307 19113 27341
rect 19085 27188 19119 27222
rect 19079 26989 19113 27023
rect 19079 26878 19113 26912
rect 19093 26793 19127 26827
rect 19067 26689 19101 26723
rect 19093 26605 19127 26639
rect 19067 26521 19101 26555
rect 19059 25919 19093 25953
rect 19097 25835 19131 25869
rect 19071 25740 19105 25774
rect 19026 25636 19060 25670
rect 19094 25636 19128 25670
rect 19067 25552 19101 25586
rect 19028 25468 19062 25502
rect 19096 25468 19130 25502
rect 19083 25362 19117 25396
rect 19083 25164 19117 25198
rect 19083 25061 19117 25095
rect 19089 24942 19123 24976
rect 19083 24743 19117 24777
rect 19083 24632 19117 24666
rect 19097 24547 19131 24581
rect 19071 24443 19105 24477
rect 19097 24359 19131 24393
rect 19071 24275 19105 24309
rect 7705 22913 7739 22947
rect 7789 22887 7823 22921
rect 7873 22913 7907 22947
rect 7977 22887 8011 22921
rect 8062 22901 8096 22935
rect 8173 22901 8207 22935
rect 8372 22895 8406 22929
rect 8491 22901 8525 22935
rect 8594 22901 8628 22935
rect 8792 22901 8826 22935
rect 8898 22956 8932 22990
rect 8898 22888 8932 22922
rect 8982 22917 9016 22951
rect 9066 22958 9100 22992
rect 9066 22890 9100 22924
rect 9170 22913 9204 22947
rect 9265 22887 9299 22921
rect 9349 22925 9383 22959
rect 9951 22917 9985 22951
rect 10035 22891 10069 22925
rect 10119 22917 10153 22951
rect 10223 22891 10257 22925
rect 10308 22905 10342 22939
rect 10419 22905 10453 22939
rect 10618 22899 10652 22933
rect 10737 22905 10771 22939
rect 10840 22905 10874 22939
rect 11038 22905 11072 22939
rect 11144 22960 11178 22994
rect 11144 22892 11178 22926
rect 11228 22921 11262 22955
rect 11312 22962 11346 22996
rect 11312 22894 11346 22928
rect 11416 22917 11450 22951
rect 11511 22891 11545 22925
rect 11595 22929 11629 22963
rect 12137 22909 12171 22943
rect 12221 22883 12255 22917
rect 12305 22909 12339 22943
rect 12409 22883 12443 22917
rect 12494 22897 12528 22931
rect 12605 22897 12639 22931
rect 12804 22891 12838 22925
rect 12923 22897 12957 22931
rect 13026 22897 13060 22931
rect 13224 22897 13258 22931
rect 13330 22952 13364 22986
rect 13330 22884 13364 22918
rect 13414 22913 13448 22947
rect 13498 22954 13532 22988
rect 13498 22886 13532 22920
rect 13602 22909 13636 22943
rect 13697 22883 13731 22917
rect 13781 22921 13815 22955
rect 14383 22913 14417 22947
rect 14467 22887 14501 22921
rect 14551 22913 14585 22947
rect 14655 22887 14689 22921
rect 14740 22901 14774 22935
rect 14851 22901 14885 22935
rect 15050 22895 15084 22929
rect 15169 22901 15203 22935
rect 15272 22901 15306 22935
rect 15470 22901 15504 22935
rect 15576 22956 15610 22990
rect 15576 22888 15610 22922
rect 15660 22917 15694 22951
rect 15744 22958 15778 22992
rect 15744 22890 15778 22924
rect 15848 22913 15882 22947
rect 15943 22887 15977 22921
rect 16027 22925 16061 22959
rect 16665 22913 16699 22947
rect 16749 22887 16783 22921
rect 16833 22913 16867 22947
rect 16937 22887 16971 22921
rect 17022 22901 17056 22935
rect 17133 22901 17167 22935
rect 17332 22895 17366 22929
rect 17451 22901 17485 22935
rect 17554 22901 17588 22935
rect 17752 22901 17786 22935
rect 17858 22956 17892 22990
rect 17858 22888 17892 22922
rect 17942 22917 17976 22951
rect 18026 22958 18060 22992
rect 18026 22890 18060 22924
rect 18130 22913 18164 22947
rect 18225 22887 18259 22921
rect 18309 22925 18343 22959
rect 9512 17697 9546 17731
rect 9512 17629 9546 17663
rect 9596 17697 9630 17731
rect 9596 17629 9630 17663
rect 15649 17549 15683 17583
rect 15649 17481 15683 17515
rect 15733 17549 15767 17583
rect 16427 17587 16461 17621
rect 16427 17519 16461 17553
rect 15733 17481 15767 17515
rect 16511 17587 16545 17621
rect 16511 17519 16545 17553
rect 17301 17589 17335 17623
rect 17301 17521 17335 17555
rect 17385 17589 17419 17623
rect 17385 17521 17419 17555
rect 18069 17579 18103 17613
rect 18069 17511 18103 17545
rect 18153 17579 18187 17613
rect 18153 17511 18187 17545
rect 19191 17581 19225 17615
rect 19191 17513 19225 17547
rect 19275 17581 19309 17615
rect 19275 17513 19309 17547
rect 20065 17583 20099 17617
rect 20065 17515 20099 17549
rect 20149 17583 20183 17617
rect 20149 17515 20183 17549
rect 20833 17573 20867 17607
rect 20833 17505 20867 17539
rect 20917 17573 20951 17607
rect 20917 17505 20951 17539
rect 21447 17571 21481 17605
rect 21447 17503 21481 17537
rect 21531 17571 21565 17605
rect 21531 17503 21565 17537
rect 22321 17573 22355 17607
rect 22321 17505 22355 17539
rect 22405 17573 22439 17607
rect 22405 17505 22439 17539
rect 23089 17563 23123 17597
rect 23089 17495 23123 17529
rect 23173 17563 23207 17597
rect 23173 17495 23207 17529
rect 4511 16103 4545 16137
rect 4595 16125 4629 16159
rect 4679 16103 4713 16137
rect 4847 16105 4881 16139
rect 4947 16105 4981 16139
rect 5037 16176 5071 16210
rect 5037 16108 5071 16142
rect 9377 16107 9411 16141
rect 9461 16129 9495 16163
rect 9545 16107 9579 16141
rect 9713 16109 9747 16143
rect 9813 16109 9847 16143
rect 16412 16281 16446 16315
rect 9903 16180 9937 16214
rect 16412 16213 16446 16247
rect 16496 16281 16530 16315
rect 16496 16213 16530 16247
rect 17180 16271 17214 16305
rect 17180 16203 17214 16237
rect 17264 16271 17298 16305
rect 17264 16203 17298 16237
rect 18054 16273 18088 16307
rect 18054 16205 18088 16239
rect 18138 16273 18172 16307
rect 18138 16205 18172 16239
rect 18668 16271 18702 16305
rect 18668 16203 18702 16237
rect 18752 16271 18786 16305
rect 18752 16203 18786 16237
rect 19436 16261 19470 16295
rect 19436 16193 19470 16227
rect 19520 16261 19554 16295
rect 19520 16193 19554 16227
rect 20310 16263 20344 16297
rect 20310 16195 20344 16229
rect 20394 16263 20428 16297
rect 20394 16195 20428 16229
rect 21432 16265 21466 16299
rect 21432 16197 21466 16231
rect 21516 16265 21550 16299
rect 21516 16197 21550 16231
rect 22200 16255 22234 16289
rect 22200 16187 22234 16221
rect 22284 16255 22318 16289
rect 22284 16187 22318 16221
rect 23074 16257 23108 16291
rect 23074 16189 23108 16223
rect 23158 16257 23192 16291
rect 23158 16189 23192 16223
rect 9903 16112 9937 16146
rect 4637 15385 4671 15419
rect 4829 15357 4863 15391
rect 4913 15357 4947 15391
rect 9503 15389 9537 15423
rect 6643 15255 6677 15289
rect 7084 15315 7118 15349
rect 7084 15247 7118 15281
rect 7183 15315 7217 15349
rect 7183 15247 7217 15281
rect 9695 15361 9729 15395
rect 9779 15361 9813 15395
rect 11509 15259 11543 15293
rect 11950 15319 11984 15353
rect 11950 15251 11984 15285
rect 12049 15319 12083 15353
rect 12049 15251 12083 15285
rect 5821 14775 5855 14809
rect 6013 14747 6047 14781
rect 6097 14747 6131 14781
rect 10687 14779 10721 14813
rect 10879 14751 10913 14785
rect 10963 14751 10997 14785
rect 4521 14539 4555 14573
rect 4605 14561 4639 14595
rect 4689 14539 4723 14573
rect 4857 14541 4891 14575
rect 4957 14541 4991 14575
rect 5047 14612 5081 14646
rect 5047 14544 5081 14578
rect 9387 14543 9421 14577
rect 9471 14565 9505 14599
rect 9555 14543 9589 14577
rect 9723 14545 9757 14579
rect 9823 14545 9857 14579
rect 9913 14616 9947 14650
rect 9913 14548 9947 14582
rect 23519 14356 23553 14390
rect 23603 14347 23637 14381
rect 23784 14407 23818 14441
rect 23868 14381 23902 14415
rect 23972 14390 24006 14424
rect 24056 14399 24090 14433
rect 24160 14397 24194 14431
rect 24244 14423 24278 14457
rect 24328 14423 24362 14457
rect 24430 14347 24464 14381
rect 24514 14347 24548 14381
rect 24598 14363 24632 14397
rect 24702 14347 24736 14381
rect 24786 14369 24820 14403
rect 24890 14355 24924 14389
rect 25030 14355 25064 14389
rect 25127 14423 25161 14457
rect 25263 14347 25297 14381
rect 25347 14355 25381 14389
rect 4647 13821 4681 13855
rect 4839 13793 4873 13827
rect 4923 13793 4957 13827
rect 5859 13789 5893 13823
rect 6300 13849 6334 13883
rect 6300 13781 6334 13815
rect 6399 13849 6433 13883
rect 6399 13781 6433 13815
rect 7757 13789 7791 13823
rect 7847 13783 7881 13817
rect 7937 13769 7971 13803
rect 8021 13783 8055 13817
rect 8115 13769 8149 13803
rect 8203 13807 8237 13841
rect 9513 13825 9547 13859
rect 9705 13797 9739 13831
rect 9789 13797 9823 13831
rect 10725 13793 10759 13827
rect 11166 13853 11200 13887
rect 11166 13785 11200 13819
rect 11265 13853 11299 13887
rect 11265 13785 11299 13819
rect 12623 13793 12657 13827
rect 12713 13787 12747 13821
rect 12803 13773 12837 13807
rect 12887 13787 12921 13821
rect 12981 13773 13015 13807
rect 13069 13811 13103 13845
rect 6858 13417 6892 13451
rect 6942 13417 6976 13451
rect 7038 13417 7072 13451
rect 7123 13477 7157 13511
rect 7123 13409 7157 13443
rect 11724 13421 11758 13455
rect 11808 13421 11842 13455
rect 11904 13421 11938 13455
rect 11989 13481 12023 13515
rect 11989 13413 12023 13447
rect 4513 12871 4547 12905
rect 4597 12893 4631 12927
rect 4681 12871 4715 12905
rect 4849 12873 4883 12907
rect 4949 12873 4983 12907
rect 5039 12944 5073 12978
rect 5983 12939 6017 12973
rect 6255 12955 6289 12989
rect 6339 12965 6373 12999
rect 5039 12876 5073 12910
rect 9379 12875 9413 12909
rect 9463 12897 9497 12931
rect 9547 12875 9581 12909
rect 9715 12877 9749 12911
rect 9815 12877 9849 12911
rect 9905 12948 9939 12982
rect 10849 12943 10883 12977
rect 11121 12959 11155 12993
rect 11205 12969 11239 13003
rect 9905 12880 9939 12914
rect 4639 12153 4673 12187
rect 4831 12125 4865 12159
rect 4915 12125 4949 12159
rect 9505 12157 9539 12191
rect 9697 12129 9731 12163
rect 9781 12129 9815 12163
rect 6015 11947 6049 11981
rect 6207 11919 6241 11953
rect 6291 11919 6325 11953
rect 10881 11951 10915 11985
rect 11073 11923 11107 11957
rect 11157 11923 11191 11957
rect 4523 11307 4557 11341
rect 4607 11329 4641 11363
rect 4691 11307 4725 11341
rect 4859 11309 4893 11343
rect 4959 11309 4993 11343
rect 5049 11380 5083 11414
rect 5049 11312 5083 11346
rect 9389 11311 9423 11345
rect 9473 11333 9507 11367
rect 9557 11311 9591 11345
rect 9725 11313 9759 11347
rect 9825 11313 9859 11347
rect 9915 11384 9949 11418
rect 9915 11316 9949 11350
rect 4649 10589 4683 10623
rect 4841 10561 4875 10595
rect 4925 10561 4959 10595
rect 9515 10593 9549 10627
rect 9707 10565 9741 10599
rect 9791 10565 9825 10599
rect 6194 6503 6228 6537
rect 6194 6435 6228 6469
rect 6278 6503 6312 6537
rect 6278 6435 6312 6469
rect 10088 5839 10122 5873
rect 10187 5879 10221 5913
rect 10439 5867 10473 5901
rect 10540 5862 10574 5896
rect 10624 5879 10658 5913
rect 10708 5862 10742 5896
rect 10792 5870 10826 5904
rect 10896 5862 10930 5896
rect 10980 5879 11014 5913
rect 11064 5862 11098 5896
rect 11148 5862 11182 5896
rect 11337 5875 11371 5909
rect 1906 5419 1940 5453
rect 2005 5459 2039 5493
rect 2257 5447 2291 5481
rect 2358 5442 2392 5476
rect 2442 5459 2476 5493
rect 2526 5442 2560 5476
rect 2610 5450 2644 5484
rect 2714 5442 2748 5476
rect 2798 5459 2832 5493
rect 2882 5442 2916 5476
rect 2966 5442 3000 5476
rect 3155 5455 3189 5489
rect 3239 5419 3273 5453
rect 4040 5411 4074 5445
rect 4139 5451 4173 5485
rect 4391 5439 4425 5473
rect 4492 5434 4526 5468
rect 4576 5451 4610 5485
rect 4660 5434 4694 5468
rect 4744 5442 4778 5476
rect 4848 5434 4882 5468
rect 4932 5451 4966 5485
rect 5016 5434 5050 5468
rect 5100 5434 5134 5468
rect 5289 5447 5323 5481
rect 5373 5411 5407 5445
rect 5992 5411 6026 5445
rect 6091 5451 6125 5485
rect 6343 5439 6377 5473
rect 6444 5434 6478 5468
rect 6528 5451 6562 5485
rect 6612 5434 6646 5468
rect 6696 5442 6730 5476
rect 6800 5434 6834 5468
rect 6884 5451 6918 5485
rect 6968 5434 7002 5468
rect 7052 5434 7086 5468
rect 7241 5447 7275 5481
rect 7325 5411 7359 5445
rect 7994 5417 8028 5451
rect 8093 5457 8127 5491
rect 8345 5445 8379 5479
rect 8446 5440 8480 5474
rect 8530 5457 8564 5491
rect 8614 5440 8648 5474
rect 8698 5448 8732 5482
rect 8802 5440 8836 5474
rect 8886 5457 8920 5491
rect 8970 5440 9004 5474
rect 9054 5440 9088 5474
rect 9243 5453 9277 5487
rect 11421 5839 11455 5873
rect 12150 5827 12184 5861
rect 12249 5867 12283 5901
rect 12501 5855 12535 5889
rect 12602 5850 12636 5884
rect 12686 5867 12720 5901
rect 12770 5850 12804 5884
rect 12854 5858 12888 5892
rect 12958 5850 12992 5884
rect 13042 5867 13076 5901
rect 13126 5850 13160 5884
rect 13210 5850 13244 5884
rect 13399 5863 13433 5897
rect 9327 5417 9361 5451
rect 13483 5827 13517 5861
rect 14108 5835 14142 5869
rect 14207 5875 14241 5909
rect 14459 5863 14493 5897
rect 14560 5858 14594 5892
rect 14644 5875 14678 5909
rect 14728 5858 14762 5892
rect 14812 5866 14846 5900
rect 14916 5858 14950 5892
rect 15000 5875 15034 5909
rect 15084 5858 15118 5892
rect 15168 5858 15202 5892
rect 15357 5871 15391 5905
rect 15441 5835 15475 5869
rect 16102 5841 16136 5875
rect 16201 5881 16235 5915
rect 16453 5869 16487 5903
rect 16554 5864 16588 5898
rect 16638 5881 16672 5915
rect 16722 5864 16756 5898
rect 16806 5872 16840 5906
rect 16910 5864 16944 5898
rect 16994 5881 17028 5915
rect 17078 5864 17112 5898
rect 17162 5864 17196 5898
rect 17351 5877 17385 5911
rect 17435 5841 17469 5875
rect 18383 5288 18417 5322
rect 18467 5288 18501 5322
rect 18535 5288 18569 5322
rect 18770 5288 18804 5322
rect 18977 5303 19011 5337
rect 10116 4965 10150 4999
rect 10215 5005 10249 5039
rect 10467 4993 10501 5027
rect 10568 4988 10602 5022
rect 10652 5005 10686 5039
rect 10736 4988 10770 5022
rect 10820 4996 10854 5030
rect 10924 4988 10958 5022
rect 11008 5005 11042 5039
rect 11092 4988 11126 5022
rect 11176 4988 11210 5022
rect 11365 5001 11399 5035
rect 11449 4965 11483 4999
rect 12386 4921 12420 4955
rect 12485 4961 12519 4995
rect 12737 4949 12771 4983
rect 12838 4944 12872 4978
rect 12922 4961 12956 4995
rect 13006 4944 13040 4978
rect 13090 4952 13124 4986
rect 13194 4944 13228 4978
rect 13278 4961 13312 4995
rect 13362 4944 13396 4978
rect 13446 4944 13480 4978
rect 13635 4957 13669 4991
rect 19061 5284 19095 5318
rect 13719 4921 13753 4955
rect 14388 4915 14422 4949
rect 14487 4955 14521 4989
rect 14739 4943 14773 4977
rect 14840 4938 14874 4972
rect 14924 4955 14958 4989
rect 15008 4938 15042 4972
rect 15092 4946 15126 4980
rect 15196 4938 15230 4972
rect 15280 4955 15314 4989
rect 15364 4938 15398 4972
rect 15448 4938 15482 4972
rect 15637 4951 15671 4985
rect 15721 4915 15755 4949
rect 16410 4897 16444 4931
rect 16509 4937 16543 4971
rect 16761 4925 16795 4959
rect 16862 4920 16896 4954
rect 16946 4937 16980 4971
rect 17030 4920 17064 4954
rect 17114 4928 17148 4962
rect 17218 4920 17252 4954
rect 17302 4937 17336 4971
rect 17386 4920 17420 4954
rect 17470 4920 17504 4954
rect 17659 4933 17693 4967
rect 17743 4897 17777 4931
rect 6164 3243 6198 3277
rect 6164 3175 6198 3209
rect 6248 3243 6282 3277
rect 6248 3175 6282 3209
rect 1876 2159 1910 2193
rect 1975 2199 2009 2233
rect 2227 2187 2261 2221
rect 2328 2182 2362 2216
rect 2412 2199 2446 2233
rect 2496 2182 2530 2216
rect 2580 2190 2614 2224
rect 2684 2182 2718 2216
rect 2768 2199 2802 2233
rect 2852 2182 2886 2216
rect 2936 2182 2970 2216
rect 3125 2195 3159 2229
rect 3209 2159 3243 2193
rect 3946 2155 3980 2189
rect 4045 2195 4079 2229
rect 4297 2183 4331 2217
rect 4398 2178 4432 2212
rect 4482 2195 4516 2229
rect 4566 2178 4600 2212
rect 4650 2186 4684 2220
rect 4754 2178 4788 2212
rect 4838 2195 4872 2229
rect 4922 2178 4956 2212
rect 5006 2178 5040 2212
rect 5195 2191 5229 2225
rect 5279 2155 5313 2189
rect 5898 2155 5932 2189
rect 5997 2195 6031 2229
rect 6249 2183 6283 2217
rect 6350 2178 6384 2212
rect 6434 2195 6468 2229
rect 6518 2178 6552 2212
rect 6602 2186 6636 2220
rect 6706 2178 6740 2212
rect 6790 2195 6824 2229
rect 6874 2178 6908 2212
rect 6958 2178 6992 2212
rect 7147 2191 7181 2225
rect 7231 2155 7265 2189
rect 7900 2161 7934 2195
rect 7999 2201 8033 2235
rect 8251 2189 8285 2223
rect 8352 2184 8386 2218
rect 8436 2201 8470 2235
rect 8520 2184 8554 2218
rect 8604 2192 8638 2226
rect 8708 2184 8742 2218
rect 8792 2201 8826 2235
rect 8876 2184 8910 2218
rect 8960 2184 8994 2218
rect 9149 2197 9183 2231
rect 9233 2161 9267 2195
rect 9852 2161 9886 2195
rect 9951 2201 9985 2235
rect 10203 2189 10237 2223
rect 10304 2184 10338 2218
rect 10388 2201 10422 2235
rect 10472 2184 10506 2218
rect 10556 2192 10590 2226
rect 10660 2184 10694 2218
rect 10744 2201 10778 2235
rect 10828 2184 10862 2218
rect 10912 2184 10946 2218
rect 11101 2197 11135 2231
rect 11185 2161 11219 2195
rect 11844 2161 11878 2195
rect 11943 2201 11977 2235
rect 12195 2189 12229 2223
rect 12296 2184 12330 2218
rect 12380 2201 12414 2235
rect 12464 2184 12498 2218
rect 12548 2192 12582 2226
rect 12652 2184 12686 2218
rect 12736 2201 12770 2235
rect 12820 2184 12854 2218
rect 12904 2184 12938 2218
rect 13093 2197 13127 2231
rect 13177 2161 13211 2195
rect 13796 2161 13830 2195
rect 13895 2201 13929 2235
rect 14147 2189 14181 2223
rect 14248 2184 14282 2218
rect 14332 2201 14366 2235
rect 14416 2184 14450 2218
rect 14500 2192 14534 2226
rect 14604 2184 14638 2218
rect 14688 2201 14722 2235
rect 14772 2184 14806 2218
rect 14856 2184 14890 2218
rect 15045 2197 15079 2231
rect 15129 2161 15163 2195
rect 15860 2161 15894 2195
rect 15959 2201 15993 2235
rect 16211 2189 16245 2223
rect 16312 2184 16346 2218
rect 16396 2201 16430 2235
rect 16480 2184 16514 2218
rect 16564 2192 16598 2226
rect 16668 2184 16702 2218
rect 16752 2201 16786 2235
rect 16836 2184 16870 2218
rect 16920 2184 16954 2218
rect 17109 2197 17143 2231
rect 17193 2161 17227 2195
<< pdiffc >>
rect 18655 43340 18689 43374
rect 18723 43340 18757 43374
rect 18655 43256 18689 43290
rect 18723 43256 18757 43290
rect 18793 43256 18827 43290
rect 18655 43172 18689 43206
rect 18723 43172 18757 43206
rect 18655 43088 18689 43122
rect 18723 43088 18757 43122
rect 18793 43088 18827 43122
rect 18655 43004 18689 43038
rect 18723 43004 18757 43038
rect 18655 42920 18689 42954
rect 18723 42920 18757 42954
rect 18793 42920 18827 42954
rect 18655 42836 18689 42870
rect 18723 42836 18757 42870
rect 18655 42752 18689 42786
rect 18723 42752 18757 42786
rect 18793 42752 18827 42786
rect 18655 42668 18689 42702
rect 18723 42668 18757 42702
rect 18655 42584 18689 42618
rect 18723 42584 18757 42618
rect 18793 42584 18827 42618
rect 18655 42500 18689 42534
rect 18723 42500 18757 42534
rect 18655 42416 18689 42450
rect 18723 42416 18757 42450
rect 18793 42416 18827 42450
rect 18655 42332 18689 42366
rect 18723 42332 18757 42366
rect 18655 42248 18689 42282
rect 18723 42248 18757 42282
rect 18793 42248 18827 42282
rect 18655 42164 18689 42198
rect 18723 42164 18757 42198
rect 18655 42080 18689 42114
rect 18723 42080 18757 42114
rect 18793 42080 18827 42114
rect 18655 41996 18689 42030
rect 18723 41996 18757 42030
rect 18793 41996 18827 42030
rect 18639 41363 18673 41397
rect 18707 41363 18741 41397
rect 18639 41228 18673 41262
rect 18707 41228 18741 41262
rect 18775 41228 18809 41262
rect 18639 41144 18673 41178
rect 18707 41144 18741 41178
rect 18639 41060 18673 41094
rect 18707 41060 18741 41094
rect 18775 41060 18809 41094
rect 18639 40976 18673 41010
rect 18707 40976 18741 41010
rect 18639 40892 18673 40926
rect 18707 40892 18741 40926
rect 18775 40892 18809 40926
rect 18639 40808 18673 40842
rect 18707 40808 18741 40842
rect 18639 40724 18673 40758
rect 18707 40724 18741 40758
rect 18775 40724 18809 40758
rect 18639 40640 18673 40674
rect 18707 40640 18741 40674
rect 18639 40556 18673 40590
rect 18707 40556 18741 40590
rect 18775 40556 18809 40590
rect 18639 40472 18673 40506
rect 18707 40472 18741 40506
rect 18639 40388 18673 40422
rect 18707 40388 18741 40422
rect 18775 40388 18809 40422
rect 18639 40304 18673 40338
rect 18707 40304 18741 40338
rect 18647 39548 18681 39582
rect 18715 39548 18749 39582
rect 18647 39464 18681 39498
rect 18715 39464 18749 39498
rect 18783 39464 18817 39498
rect 18647 39380 18681 39414
rect 18715 39380 18749 39414
rect 18647 39296 18681 39330
rect 18715 39296 18749 39330
rect 18783 39296 18817 39330
rect 18647 39212 18681 39246
rect 18715 39212 18749 39246
rect 18647 39128 18681 39162
rect 18715 39128 18749 39162
rect 18783 39128 18817 39162
rect 18647 39044 18681 39078
rect 18715 39044 18749 39078
rect 18647 38960 18681 38994
rect 18715 38960 18749 38994
rect 18783 38960 18817 38994
rect 18647 38876 18681 38910
rect 18715 38876 18749 38910
rect 18661 38303 18695 38337
rect 18661 38219 18695 38253
rect 18729 38219 18763 38253
rect 18797 38219 18831 38253
rect 18661 38135 18695 38169
rect 18729 38135 18763 38169
rect 18661 38051 18695 38085
rect 18729 38051 18763 38085
rect 18797 38051 18831 38085
rect 18661 37967 18695 38001
rect 18729 37967 18763 38001
rect 18661 37883 18695 37917
rect 18729 37883 18763 37917
rect 18797 37883 18831 37917
rect 18661 37765 18695 37799
rect 18729 37765 18763 37799
rect 18797 37765 18831 37799
rect 18673 37145 18707 37179
rect 18673 37061 18707 37095
rect 18741 37061 18775 37095
rect 18809 37061 18843 37095
rect 18673 36977 18707 37011
rect 18741 36977 18775 37011
rect 18673 36893 18707 36927
rect 18741 36893 18775 36927
rect 18809 36893 18843 36927
rect 18673 36809 18707 36843
rect 18741 36809 18775 36843
rect 18809 36809 18843 36843
rect 18681 36265 18715 36299
rect 18749 36265 18783 36299
rect 18817 36265 18851 36299
rect 18681 36181 18715 36215
rect 18749 36181 18783 36215
rect 18817 36181 18851 36215
rect 18681 36097 18715 36131
rect 18749 36097 18783 36131
rect 18817 36097 18851 36131
rect 18705 34879 18739 34913
rect 18776 34879 18810 34913
rect 18847 34879 18881 34913
rect 18705 34795 18739 34829
rect 18773 34795 18807 34829
rect 18841 34795 18875 34829
rect 18705 34698 18739 34732
rect 18773 34698 18807 34732
rect 18711 34594 18745 34628
rect 18779 34594 18813 34628
rect 18847 34594 18881 34628
rect 18735 34510 18769 34544
rect 18815 34510 18849 34544
rect 18705 34424 18739 34458
rect 18776 34424 18810 34458
rect 18847 34424 18881 34458
rect 18713 34300 18747 34334
rect 18723 34101 18757 34135
rect 18713 34006 18747 34040
rect 18705 33922 18739 33956
rect 18773 33922 18807 33956
rect 18718 33683 18752 33717
rect 18713 33591 18747 33625
rect 18705 33507 18739 33541
rect 18713 33403 18747 33437
rect 18781 33403 18815 33437
rect 18729 33319 18763 33353
rect 18713 33235 18747 33269
rect 18781 33235 18815 33269
rect 18705 32597 18739 32631
rect 18776 32597 18810 32631
rect 18847 32597 18881 32631
rect 18705 32513 18739 32547
rect 18773 32513 18807 32547
rect 18841 32513 18875 32547
rect 18705 32416 18739 32450
rect 18773 32416 18807 32450
rect 18711 32312 18745 32346
rect 18779 32312 18813 32346
rect 18847 32312 18881 32346
rect 18735 32228 18769 32262
rect 18815 32228 18849 32262
rect 18705 32142 18739 32176
rect 18776 32142 18810 32176
rect 18847 32142 18881 32176
rect 18713 32018 18747 32052
rect 18723 31819 18757 31853
rect 18713 31724 18747 31758
rect 18705 31640 18739 31674
rect 18773 31640 18807 31674
rect 18718 31401 18752 31435
rect 18713 31309 18747 31343
rect 18705 31225 18739 31259
rect 18713 31121 18747 31155
rect 18781 31121 18815 31155
rect 18729 31037 18763 31071
rect 18713 30953 18747 30987
rect 18781 30953 18815 30987
rect 18709 30351 18743 30385
rect 18780 30351 18814 30385
rect 18851 30351 18885 30385
rect 18709 30267 18743 30301
rect 18777 30267 18811 30301
rect 18845 30267 18879 30301
rect 18709 30170 18743 30204
rect 18777 30170 18811 30204
rect 18715 30066 18749 30100
rect 18783 30066 18817 30100
rect 18851 30066 18885 30100
rect 18739 29982 18773 30016
rect 18819 29982 18853 30016
rect 18709 29896 18743 29930
rect 18780 29896 18814 29930
rect 18851 29896 18885 29930
rect 18717 29772 18751 29806
rect 18727 29573 18761 29607
rect 18717 29478 18751 29512
rect 18709 29394 18743 29428
rect 18777 29394 18811 29428
rect 18722 29155 18756 29189
rect 18717 29063 18751 29097
rect 18709 28979 18743 29013
rect 18717 28875 18751 28909
rect 18785 28875 18819 28909
rect 18733 28791 18767 28825
rect 18717 28707 18751 28741
rect 18785 28707 18819 28741
rect 18701 28165 18735 28199
rect 18772 28165 18806 28199
rect 18843 28165 18877 28199
rect 18701 28081 18735 28115
rect 18769 28081 18803 28115
rect 18837 28081 18871 28115
rect 18701 27984 18735 28018
rect 18769 27984 18803 28018
rect 18707 27880 18741 27914
rect 18775 27880 18809 27914
rect 18843 27880 18877 27914
rect 18731 27796 18765 27830
rect 18811 27796 18845 27830
rect 18701 27710 18735 27744
rect 18772 27710 18806 27744
rect 18843 27710 18877 27744
rect 18709 27586 18743 27620
rect 18719 27387 18753 27421
rect 18709 27292 18743 27326
rect 18701 27208 18735 27242
rect 18769 27208 18803 27242
rect 18714 26969 18748 27003
rect 18709 26877 18743 26911
rect 18701 26793 18735 26827
rect 18709 26689 18743 26723
rect 18777 26689 18811 26723
rect 18725 26605 18759 26639
rect 18709 26521 18743 26555
rect 18777 26521 18811 26555
rect 18705 25919 18739 25953
rect 18776 25919 18810 25953
rect 18847 25919 18881 25953
rect 18705 25835 18739 25869
rect 18773 25835 18807 25869
rect 18841 25835 18875 25869
rect 18705 25738 18739 25772
rect 18773 25738 18807 25772
rect 18711 25634 18745 25668
rect 18779 25634 18813 25668
rect 18847 25634 18881 25668
rect 18735 25550 18769 25584
rect 18815 25550 18849 25584
rect 18705 25464 18739 25498
rect 18776 25464 18810 25498
rect 18847 25464 18881 25498
rect 18713 25340 18747 25374
rect 18723 25141 18757 25175
rect 18713 25046 18747 25080
rect 18705 24962 18739 24996
rect 18773 24962 18807 24996
rect 18718 24723 18752 24757
rect 18713 24631 18747 24665
rect 18705 24547 18739 24581
rect 18713 24443 18747 24477
rect 18781 24443 18815 24477
rect 18729 24359 18763 24393
rect 18713 24275 18747 24309
rect 18781 24275 18815 24309
rect 7705 23271 7739 23305
rect 7705 23203 7739 23237
rect 7789 23255 7823 23289
rect 7873 23271 7907 23305
rect 7977 23279 8011 23313
rect 8061 23271 8095 23305
rect 8153 23266 8187 23300
rect 8392 23279 8426 23313
rect 7873 23203 7907 23237
rect 8392 23211 8426 23245
rect 8476 23271 8510 23305
rect 8571 23261 8605 23295
rect 8770 23271 8804 23305
rect 8894 23279 8928 23313
rect 8894 23208 8928 23242
rect 8894 23137 8928 23171
rect 8980 23249 9014 23283
rect 8980 23169 9014 23203
rect 9064 23273 9098 23307
rect 9064 23205 9098 23239
rect 9168 23279 9202 23313
rect 9168 23211 9202 23245
rect 9265 23279 9299 23313
rect 9265 23211 9299 23245
rect 9064 23137 9098 23171
rect 9265 23143 9299 23177
rect 9349 23279 9383 23313
rect 9349 23208 9383 23242
rect 9349 23137 9383 23171
rect 9951 23275 9985 23309
rect 9951 23207 9985 23241
rect 10035 23259 10069 23293
rect 10119 23275 10153 23309
rect 10223 23283 10257 23317
rect 10307 23275 10341 23309
rect 10399 23270 10433 23304
rect 10638 23283 10672 23317
rect 10119 23207 10153 23241
rect 10638 23215 10672 23249
rect 10722 23275 10756 23309
rect 10817 23265 10851 23299
rect 11016 23275 11050 23309
rect 11140 23283 11174 23317
rect 11140 23212 11174 23246
rect 11140 23141 11174 23175
rect 11226 23253 11260 23287
rect 11226 23173 11260 23207
rect 11310 23277 11344 23311
rect 11310 23209 11344 23243
rect 11414 23283 11448 23317
rect 11414 23215 11448 23249
rect 11511 23283 11545 23317
rect 11511 23215 11545 23249
rect 11310 23141 11344 23175
rect 11511 23147 11545 23181
rect 11595 23283 11629 23317
rect 11595 23212 11629 23246
rect 11595 23141 11629 23175
rect 12137 23267 12171 23301
rect 12137 23199 12171 23233
rect 12221 23251 12255 23285
rect 12305 23267 12339 23301
rect 12409 23275 12443 23309
rect 12493 23267 12527 23301
rect 12585 23262 12619 23296
rect 12824 23275 12858 23309
rect 12305 23199 12339 23233
rect 12824 23207 12858 23241
rect 12908 23267 12942 23301
rect 13003 23257 13037 23291
rect 13202 23267 13236 23301
rect 13326 23275 13360 23309
rect 13326 23204 13360 23238
rect 13326 23133 13360 23167
rect 13412 23245 13446 23279
rect 13412 23165 13446 23199
rect 13496 23269 13530 23303
rect 13496 23201 13530 23235
rect 13600 23275 13634 23309
rect 13600 23207 13634 23241
rect 13697 23275 13731 23309
rect 13697 23207 13731 23241
rect 13496 23133 13530 23167
rect 13697 23139 13731 23173
rect 13781 23275 13815 23309
rect 13781 23204 13815 23238
rect 13781 23133 13815 23167
rect 14383 23271 14417 23305
rect 14383 23203 14417 23237
rect 14467 23255 14501 23289
rect 14551 23271 14585 23305
rect 14655 23279 14689 23313
rect 14739 23271 14773 23305
rect 14831 23266 14865 23300
rect 15070 23279 15104 23313
rect 14551 23203 14585 23237
rect 15070 23211 15104 23245
rect 15154 23271 15188 23305
rect 15249 23261 15283 23295
rect 15448 23271 15482 23305
rect 15572 23279 15606 23313
rect 15572 23208 15606 23242
rect 15572 23137 15606 23171
rect 15658 23249 15692 23283
rect 15658 23169 15692 23203
rect 15742 23273 15776 23307
rect 15742 23205 15776 23239
rect 15846 23279 15880 23313
rect 15846 23211 15880 23245
rect 15943 23279 15977 23313
rect 15943 23211 15977 23245
rect 15742 23137 15776 23171
rect 15943 23143 15977 23177
rect 16027 23279 16061 23313
rect 16027 23208 16061 23242
rect 16027 23137 16061 23171
rect 16665 23271 16699 23305
rect 16665 23203 16699 23237
rect 16749 23255 16783 23289
rect 16833 23271 16867 23305
rect 16937 23279 16971 23313
rect 17021 23271 17055 23305
rect 17113 23266 17147 23300
rect 17352 23279 17386 23313
rect 16833 23203 16867 23237
rect 17352 23211 17386 23245
rect 17436 23271 17470 23305
rect 17531 23261 17565 23295
rect 17730 23271 17764 23305
rect 17854 23279 17888 23313
rect 17854 23208 17888 23242
rect 17854 23137 17888 23171
rect 17940 23249 17974 23283
rect 17940 23169 17974 23203
rect 18024 23273 18058 23307
rect 18024 23205 18058 23239
rect 18128 23279 18162 23313
rect 18128 23211 18162 23245
rect 18225 23279 18259 23313
rect 18225 23211 18259 23245
rect 18024 23137 18058 23171
rect 18225 23143 18259 23177
rect 18309 23279 18343 23313
rect 18309 23208 18343 23242
rect 18309 23137 18343 23171
rect 9512 17445 9546 17479
rect 9512 17377 9546 17411
rect 9512 17309 9546 17343
rect 9596 17445 9630 17479
rect 9596 17377 9630 17411
rect 9596 17309 9630 17343
rect 15649 17297 15683 17331
rect 15649 17229 15683 17263
rect 15649 17161 15683 17195
rect 15733 17297 15767 17331
rect 15733 17229 15767 17263
rect 16427 17335 16461 17369
rect 16427 17267 16461 17301
rect 15733 17161 15767 17195
rect 16427 17199 16461 17233
rect 16511 17335 16545 17369
rect 16511 17267 16545 17301
rect 16511 17199 16545 17233
rect 17301 17337 17335 17371
rect 17301 17269 17335 17303
rect 17301 17201 17335 17235
rect 17385 17337 17419 17371
rect 17385 17269 17419 17303
rect 17385 17201 17419 17235
rect 18069 17327 18103 17361
rect 18069 17259 18103 17293
rect 18069 17191 18103 17225
rect 18153 17327 18187 17361
rect 18153 17259 18187 17293
rect 18153 17191 18187 17225
rect 19191 17329 19225 17363
rect 19191 17261 19225 17295
rect 19191 17193 19225 17227
rect 19275 17329 19309 17363
rect 19275 17261 19309 17295
rect 19275 17193 19309 17227
rect 20065 17331 20099 17365
rect 20065 17263 20099 17297
rect 20065 17195 20099 17229
rect 20149 17331 20183 17365
rect 20149 17263 20183 17297
rect 20149 17195 20183 17229
rect 20833 17321 20867 17355
rect 20833 17253 20867 17287
rect 20833 17185 20867 17219
rect 20917 17321 20951 17355
rect 20917 17253 20951 17287
rect 20917 17185 20951 17219
rect 21447 17319 21481 17353
rect 21447 17251 21481 17285
rect 21447 17183 21481 17217
rect 21531 17319 21565 17353
rect 21531 17251 21565 17285
rect 21531 17183 21565 17217
rect 22321 17321 22355 17355
rect 22321 17253 22355 17287
rect 22321 17185 22355 17219
rect 22405 17321 22439 17355
rect 22405 17253 22439 17287
rect 22405 17185 22439 17219
rect 23089 17311 23123 17345
rect 23089 17243 23123 17277
rect 23089 17175 23123 17209
rect 23173 17311 23207 17345
rect 23173 17243 23207 17277
rect 23173 17175 23207 17209
rect 4511 16493 4545 16527
rect 4511 16425 4545 16459
rect 4679 16483 4713 16517
rect 4679 16415 4713 16449
rect 4763 16483 4797 16517
rect 4763 16415 4797 16449
rect 4847 16483 4881 16517
rect 4951 16483 4985 16517
rect 4951 16415 4985 16449
rect 5035 16485 5069 16519
rect 5035 16417 5069 16451
rect 5035 16349 5069 16383
rect 9377 16497 9411 16531
rect 9377 16429 9411 16463
rect 9545 16487 9579 16521
rect 9545 16419 9579 16453
rect 9629 16487 9663 16521
rect 9629 16419 9663 16453
rect 9713 16487 9747 16521
rect 9817 16487 9851 16521
rect 9817 16419 9851 16453
rect 9901 16489 9935 16523
rect 16412 16601 16446 16635
rect 16412 16533 16446 16567
rect 16412 16465 16446 16499
rect 9901 16421 9935 16455
rect 16496 16601 16530 16635
rect 16496 16533 16530 16567
rect 16496 16465 16530 16499
rect 17180 16591 17214 16625
rect 17180 16523 17214 16557
rect 17180 16455 17214 16489
rect 17264 16591 17298 16625
rect 17264 16523 17298 16557
rect 17264 16455 17298 16489
rect 18054 16593 18088 16627
rect 18054 16525 18088 16559
rect 18054 16457 18088 16491
rect 18138 16593 18172 16627
rect 18138 16525 18172 16559
rect 18138 16457 18172 16491
rect 18668 16591 18702 16625
rect 18668 16523 18702 16557
rect 18668 16455 18702 16489
rect 9901 16353 9935 16387
rect 18752 16591 18786 16625
rect 18752 16523 18786 16557
rect 18752 16455 18786 16489
rect 19436 16581 19470 16615
rect 19436 16513 19470 16547
rect 19436 16445 19470 16479
rect 19520 16581 19554 16615
rect 19520 16513 19554 16547
rect 19520 16445 19554 16479
rect 20310 16583 20344 16617
rect 20310 16515 20344 16549
rect 20310 16447 20344 16481
rect 20394 16583 20428 16617
rect 20394 16515 20428 16549
rect 20394 16447 20428 16481
rect 21432 16585 21466 16619
rect 21432 16517 21466 16551
rect 21432 16449 21466 16483
rect 21516 16585 21550 16619
rect 21516 16517 21550 16551
rect 21516 16449 21550 16483
rect 22200 16575 22234 16609
rect 22200 16507 22234 16541
rect 22200 16439 22234 16473
rect 22284 16575 22318 16609
rect 22284 16507 22318 16541
rect 22284 16439 22318 16473
rect 23074 16577 23108 16611
rect 23074 16509 23108 16543
rect 23074 16441 23108 16475
rect 23158 16577 23192 16611
rect 23158 16509 23192 16543
rect 23158 16441 23192 16475
rect 4637 15707 4671 15741
rect 4721 15707 4755 15741
rect 4829 15749 4863 15783
rect 4829 15681 4863 15715
rect 4933 15749 4967 15783
rect 4933 15681 4967 15715
rect 6643 15639 6677 15673
rect 6735 15631 6769 15665
rect 6837 15639 6871 15673
rect 6932 15631 6966 15665
rect 7083 15639 7117 15673
rect 7083 15571 7117 15605
rect 7183 15639 7217 15673
rect 7183 15571 7217 15605
rect 7183 15503 7217 15537
rect 9503 15711 9537 15745
rect 9587 15711 9621 15745
rect 9695 15753 9729 15787
rect 9695 15685 9729 15719
rect 9799 15753 9833 15787
rect 9799 15685 9833 15719
rect 11509 15643 11543 15677
rect 11601 15635 11635 15669
rect 11703 15643 11737 15677
rect 11798 15635 11832 15669
rect 11949 15643 11983 15677
rect 11949 15575 11983 15609
rect 12049 15643 12083 15677
rect 12049 15575 12083 15609
rect 12049 15507 12083 15541
rect 5821 15097 5855 15131
rect 5905 15097 5939 15131
rect 6013 15139 6047 15173
rect 6013 15071 6047 15105
rect 4521 14929 4555 14963
rect 4521 14861 4555 14895
rect 4689 14919 4723 14953
rect 4689 14851 4723 14885
rect 4773 14919 4807 14953
rect 4773 14851 4807 14885
rect 4857 14919 4891 14953
rect 4961 14919 4995 14953
rect 4961 14851 4995 14885
rect 5045 14921 5079 14955
rect 5045 14853 5079 14887
rect 6117 15139 6151 15173
rect 6117 15071 6151 15105
rect 10687 15101 10721 15135
rect 10771 15101 10805 15135
rect 10879 15143 10913 15177
rect 10879 15075 10913 15109
rect 5045 14785 5079 14819
rect 9387 14933 9421 14967
rect 9387 14865 9421 14899
rect 9555 14923 9589 14957
rect 9555 14855 9589 14889
rect 9639 14923 9673 14957
rect 9639 14855 9673 14889
rect 9723 14923 9757 14957
rect 9827 14923 9861 14957
rect 9827 14855 9861 14889
rect 9911 14925 9945 14959
rect 9911 14857 9945 14891
rect 10983 15143 11017 15177
rect 10983 15075 11017 15109
rect 9911 14789 9945 14823
rect 23519 14731 23553 14765
rect 23603 14739 23637 14773
rect 23687 14731 23721 14765
rect 23791 14663 23825 14697
rect 23875 14679 23909 14713
rect 24063 14731 24097 14765
rect 24147 14739 24181 14773
rect 23959 14663 23993 14697
rect 24249 14663 24283 14697
rect 24333 14679 24367 14713
rect 24512 14739 24546 14773
rect 24596 14731 24630 14765
rect 24700 14739 24734 14773
rect 24784 14731 24818 14765
rect 24888 14731 24922 14765
rect 24972 14739 25006 14773
rect 25263 14739 25297 14773
rect 25069 14679 25103 14713
rect 25347 14731 25381 14765
rect 4647 14143 4681 14177
rect 4731 14143 4765 14177
rect 4839 14185 4873 14219
rect 4839 14117 4873 14151
rect 4943 14185 4977 14219
rect 4943 14117 4977 14151
rect 5859 14173 5893 14207
rect 5951 14165 5985 14199
rect 6053 14173 6087 14207
rect 6148 14165 6182 14199
rect 6299 14173 6333 14207
rect 6299 14105 6333 14139
rect 6399 14173 6433 14207
rect 6399 14105 6433 14139
rect 8118 14157 8152 14191
rect 8118 14089 8152 14123
rect 6399 14037 6433 14071
rect 7757 14026 7791 14060
rect 8203 14126 8237 14160
rect 8203 14058 8237 14092
rect 9513 14147 9547 14181
rect 9597 14147 9631 14181
rect 9705 14189 9739 14223
rect 9705 14121 9739 14155
rect 7039 13783 7073 13817
rect 6870 13663 6904 13697
rect 7039 13715 7073 13749
rect 9809 14189 9843 14223
rect 9809 14121 9843 14155
rect 10725 14177 10759 14211
rect 10817 14169 10851 14203
rect 10919 14177 10953 14211
rect 11014 14169 11048 14203
rect 11165 14177 11199 14211
rect 11165 14109 11199 14143
rect 11265 14177 11299 14211
rect 11265 14109 11299 14143
rect 12984 14161 13018 14195
rect 12984 14093 13018 14127
rect 11265 14041 11299 14075
rect 12623 14030 12657 14064
rect 13069 14130 13103 14164
rect 13069 14062 13103 14096
rect 7139 13799 7173 13833
rect 7139 13731 7173 13765
rect 11905 13787 11939 13821
rect 11736 13667 11770 13701
rect 11905 13719 11939 13753
rect 12005 13803 12039 13837
rect 12005 13735 12039 13769
rect 4513 13261 4547 13295
rect 4513 13193 4547 13227
rect 4681 13251 4715 13285
rect 4681 13183 4715 13217
rect 4765 13251 4799 13285
rect 4765 13183 4799 13217
rect 4849 13251 4883 13285
rect 4953 13251 4987 13285
rect 4953 13183 4987 13217
rect 5037 13253 5071 13287
rect 5037 13185 5071 13219
rect 6255 13331 6289 13365
rect 5983 13192 6017 13226
rect 6067 13222 6101 13256
rect 6160 13203 6194 13237
rect 5037 13117 5071 13151
rect 6339 13317 6373 13351
rect 6339 13249 6373 13283
rect 9379 13265 9413 13299
rect 9379 13197 9413 13231
rect 9547 13255 9581 13289
rect 9547 13187 9581 13221
rect 9631 13255 9665 13289
rect 9631 13187 9665 13221
rect 9715 13255 9749 13289
rect 9819 13255 9853 13289
rect 9819 13187 9853 13221
rect 9903 13257 9937 13291
rect 9903 13189 9937 13223
rect 11121 13335 11155 13369
rect 10849 13196 10883 13230
rect 10933 13226 10967 13260
rect 11026 13207 11060 13241
rect 9903 13121 9937 13155
rect 11205 13321 11239 13355
rect 11205 13253 11239 13287
rect 4639 12475 4673 12509
rect 4723 12475 4757 12509
rect 4831 12517 4865 12551
rect 4831 12449 4865 12483
rect 4935 12517 4969 12551
rect 4935 12449 4969 12483
rect 9505 12479 9539 12513
rect 9589 12479 9623 12513
rect 9697 12521 9731 12555
rect 9697 12453 9731 12487
rect 6015 12269 6049 12303
rect 6099 12269 6133 12303
rect 6207 12311 6241 12345
rect 6207 12243 6241 12277
rect 6311 12311 6345 12345
rect 6311 12243 6345 12277
rect 9801 12521 9835 12555
rect 9801 12453 9835 12487
rect 10881 12273 10915 12307
rect 10965 12273 10999 12307
rect 11073 12315 11107 12349
rect 11073 12247 11107 12281
rect 11177 12315 11211 12349
rect 11177 12247 11211 12281
rect 4523 11697 4557 11731
rect 4523 11629 4557 11663
rect 4691 11687 4725 11721
rect 4691 11619 4725 11653
rect 4775 11687 4809 11721
rect 4775 11619 4809 11653
rect 4859 11687 4893 11721
rect 4963 11687 4997 11721
rect 4963 11619 4997 11653
rect 5047 11689 5081 11723
rect 5047 11621 5081 11655
rect 5047 11553 5081 11587
rect 9389 11701 9423 11735
rect 9389 11633 9423 11667
rect 9557 11691 9591 11725
rect 9557 11623 9591 11657
rect 9641 11691 9675 11725
rect 9641 11623 9675 11657
rect 9725 11691 9759 11725
rect 9829 11691 9863 11725
rect 9829 11623 9863 11657
rect 9913 11693 9947 11727
rect 9913 11625 9947 11659
rect 9913 11557 9947 11591
rect 4649 10911 4683 10945
rect 4733 10911 4767 10945
rect 4841 10953 4875 10987
rect 4841 10885 4875 10919
rect 4945 10953 4979 10987
rect 4945 10885 4979 10919
rect 9515 10915 9549 10949
rect 9599 10915 9633 10949
rect 9707 10957 9741 10991
rect 9707 10889 9741 10923
rect 9811 10957 9845 10991
rect 9811 10889 9845 10923
rect 6194 6251 6228 6285
rect 6194 6183 6228 6217
rect 6194 6115 6228 6149
rect 6278 6251 6312 6285
rect 6278 6183 6312 6217
rect 6278 6115 6312 6149
rect 1906 5179 1940 5213
rect 1906 5089 1940 5123
rect 1990 5059 2024 5093
rect 2257 5071 2291 5105
rect 2358 5076 2392 5110
rect 2442 5059 2476 5093
rect 2526 5076 2560 5110
rect 2610 5063 2644 5097
rect 2714 5076 2748 5110
rect 2798 5059 2832 5093
rect 2882 5076 2916 5110
rect 2966 5076 3000 5110
rect 3155 5067 3189 5101
rect 3239 5176 3273 5210
rect 3239 5082 3273 5116
rect 4040 5171 4074 5205
rect 4040 5081 4074 5115
rect 4124 5051 4158 5085
rect 4391 5063 4425 5097
rect 4492 5068 4526 5102
rect 4576 5051 4610 5085
rect 4660 5068 4694 5102
rect 4744 5055 4778 5089
rect 4848 5068 4882 5102
rect 4932 5051 4966 5085
rect 5016 5068 5050 5102
rect 5100 5068 5134 5102
rect 5289 5059 5323 5093
rect 5373 5168 5407 5202
rect 5373 5074 5407 5108
rect 5992 5171 6026 5205
rect 5992 5081 6026 5115
rect 6076 5051 6110 5085
rect 6343 5063 6377 5097
rect 6444 5068 6478 5102
rect 6528 5051 6562 5085
rect 6612 5068 6646 5102
rect 6696 5055 6730 5089
rect 6800 5068 6834 5102
rect 6884 5051 6918 5085
rect 6968 5068 7002 5102
rect 7052 5068 7086 5102
rect 7241 5059 7275 5093
rect 7325 5168 7359 5202
rect 7325 5074 7359 5108
rect 7994 5177 8028 5211
rect 7994 5087 8028 5121
rect 10088 5599 10122 5633
rect 10088 5509 10122 5543
rect 10172 5479 10206 5513
rect 10439 5491 10473 5525
rect 10540 5496 10574 5530
rect 10624 5479 10658 5513
rect 10708 5496 10742 5530
rect 10792 5483 10826 5517
rect 10896 5496 10930 5530
rect 10980 5479 11014 5513
rect 11064 5496 11098 5530
rect 11148 5496 11182 5530
rect 11337 5487 11371 5521
rect 11421 5596 11455 5630
rect 11421 5502 11455 5536
rect 12150 5587 12184 5621
rect 12150 5497 12184 5531
rect 12234 5467 12268 5501
rect 12501 5479 12535 5513
rect 12602 5484 12636 5518
rect 12686 5467 12720 5501
rect 12770 5484 12804 5518
rect 12854 5471 12888 5505
rect 12958 5484 12992 5518
rect 13042 5467 13076 5501
rect 13126 5484 13160 5518
rect 13210 5484 13244 5518
rect 13399 5475 13433 5509
rect 13483 5584 13517 5618
rect 13483 5490 13517 5524
rect 14108 5595 14142 5629
rect 14108 5505 14142 5539
rect 14192 5475 14226 5509
rect 14459 5487 14493 5521
rect 14560 5492 14594 5526
rect 14644 5475 14678 5509
rect 14728 5492 14762 5526
rect 14812 5479 14846 5513
rect 14916 5492 14950 5526
rect 15000 5475 15034 5509
rect 15084 5492 15118 5526
rect 15168 5492 15202 5526
rect 15357 5483 15391 5517
rect 15441 5592 15475 5626
rect 15441 5498 15475 5532
rect 16102 5601 16136 5635
rect 16102 5511 16136 5545
rect 16186 5481 16220 5515
rect 16453 5493 16487 5527
rect 16554 5498 16588 5532
rect 16638 5481 16672 5515
rect 16722 5498 16756 5532
rect 16806 5485 16840 5519
rect 16910 5498 16944 5532
rect 16994 5481 17028 5515
rect 17078 5498 17112 5532
rect 17162 5498 17196 5532
rect 17351 5489 17385 5523
rect 17435 5598 17469 5632
rect 17435 5504 17469 5538
rect 8078 5057 8112 5091
rect 8345 5069 8379 5103
rect 8446 5074 8480 5108
rect 8530 5057 8564 5091
rect 8614 5074 8648 5108
rect 8698 5061 8732 5095
rect 8802 5074 8836 5108
rect 8886 5057 8920 5091
rect 8970 5074 9004 5108
rect 9054 5074 9088 5108
rect 9243 5065 9277 5099
rect 9327 5174 9361 5208
rect 9327 5080 9361 5114
rect 10116 4725 10150 4759
rect 10116 4635 10150 4669
rect 10200 4605 10234 4639
rect 10467 4617 10501 4651
rect 10568 4622 10602 4656
rect 10652 4605 10686 4639
rect 10736 4622 10770 4656
rect 10820 4609 10854 4643
rect 10924 4622 10958 4656
rect 11008 4605 11042 4639
rect 11092 4622 11126 4656
rect 11176 4622 11210 4656
rect 11365 4613 11399 4647
rect 11449 4722 11483 4756
rect 11449 4628 11483 4662
rect 12386 4681 12420 4715
rect 12386 4591 12420 4625
rect 18977 5047 19011 5081
rect 12470 4561 12504 4595
rect 12737 4573 12771 4607
rect 12838 4578 12872 4612
rect 12922 4561 12956 4595
rect 13006 4578 13040 4612
rect 13090 4565 13124 4599
rect 13194 4578 13228 4612
rect 13278 4561 13312 4595
rect 13362 4578 13396 4612
rect 13446 4578 13480 4612
rect 13635 4569 13669 4603
rect 13719 4678 13753 4712
rect 13719 4584 13753 4618
rect 14388 4675 14422 4709
rect 14388 4585 14422 4619
rect 14472 4555 14506 4589
rect 14739 4567 14773 4601
rect 14840 4572 14874 4606
rect 14924 4555 14958 4589
rect 15008 4572 15042 4606
rect 15092 4559 15126 4593
rect 15196 4572 15230 4606
rect 15280 4555 15314 4589
rect 15364 4572 15398 4606
rect 15448 4572 15482 4606
rect 15637 4563 15671 4597
rect 15721 4672 15755 4706
rect 15721 4578 15755 4612
rect 16410 4657 16444 4691
rect 16410 4567 16444 4601
rect 18383 4971 18417 5005
rect 18469 4971 18503 5005
rect 18666 4971 18700 5005
rect 18741 4971 18775 5005
rect 18977 4979 19011 5013
rect 18977 4911 19011 4945
rect 19061 5047 19095 5081
rect 19061 4979 19095 5013
rect 19061 4911 19095 4945
rect 16494 4537 16528 4571
rect 16761 4549 16795 4583
rect 16862 4554 16896 4588
rect 16946 4537 16980 4571
rect 17030 4554 17064 4588
rect 17114 4541 17148 4575
rect 17218 4554 17252 4588
rect 17302 4537 17336 4571
rect 17386 4554 17420 4588
rect 17470 4554 17504 4588
rect 17659 4545 17693 4579
rect 17743 4654 17777 4688
rect 17743 4560 17777 4594
rect 6164 2991 6198 3025
rect 6164 2923 6198 2957
rect 6164 2855 6198 2889
rect 6248 2991 6282 3025
rect 6248 2923 6282 2957
rect 6248 2855 6282 2889
rect 1876 1919 1910 1953
rect 1876 1829 1910 1863
rect 1960 1799 1994 1833
rect 2227 1811 2261 1845
rect 2328 1816 2362 1850
rect 2412 1799 2446 1833
rect 2496 1816 2530 1850
rect 2580 1803 2614 1837
rect 2684 1816 2718 1850
rect 2768 1799 2802 1833
rect 2852 1816 2886 1850
rect 2936 1816 2970 1850
rect 3125 1807 3159 1841
rect 3209 1916 3243 1950
rect 3209 1822 3243 1856
rect 3946 1915 3980 1949
rect 3946 1825 3980 1859
rect 4030 1795 4064 1829
rect 4297 1807 4331 1841
rect 4398 1812 4432 1846
rect 4482 1795 4516 1829
rect 4566 1812 4600 1846
rect 4650 1799 4684 1833
rect 4754 1812 4788 1846
rect 4838 1795 4872 1829
rect 4922 1812 4956 1846
rect 5006 1812 5040 1846
rect 5195 1803 5229 1837
rect 5279 1912 5313 1946
rect 5279 1818 5313 1852
rect 5898 1915 5932 1949
rect 5898 1825 5932 1859
rect 5982 1795 6016 1829
rect 6249 1807 6283 1841
rect 6350 1812 6384 1846
rect 6434 1795 6468 1829
rect 6518 1812 6552 1846
rect 6602 1799 6636 1833
rect 6706 1812 6740 1846
rect 6790 1795 6824 1829
rect 6874 1812 6908 1846
rect 6958 1812 6992 1846
rect 7147 1803 7181 1837
rect 7231 1912 7265 1946
rect 7231 1818 7265 1852
rect 7900 1921 7934 1955
rect 7900 1831 7934 1865
rect 7984 1801 8018 1835
rect 8251 1813 8285 1847
rect 8352 1818 8386 1852
rect 8436 1801 8470 1835
rect 8520 1818 8554 1852
rect 8604 1805 8638 1839
rect 8708 1818 8742 1852
rect 8792 1801 8826 1835
rect 8876 1818 8910 1852
rect 8960 1818 8994 1852
rect 9149 1809 9183 1843
rect 9233 1918 9267 1952
rect 9233 1824 9267 1858
rect 9852 1921 9886 1955
rect 9852 1831 9886 1865
rect 9936 1801 9970 1835
rect 10203 1813 10237 1847
rect 10304 1818 10338 1852
rect 10388 1801 10422 1835
rect 10472 1818 10506 1852
rect 10556 1805 10590 1839
rect 10660 1818 10694 1852
rect 10744 1801 10778 1835
rect 10828 1818 10862 1852
rect 10912 1818 10946 1852
rect 11101 1809 11135 1843
rect 11185 1918 11219 1952
rect 11185 1824 11219 1858
rect 11844 1921 11878 1955
rect 11844 1831 11878 1865
rect 11928 1801 11962 1835
rect 12195 1813 12229 1847
rect 12296 1818 12330 1852
rect 12380 1801 12414 1835
rect 12464 1818 12498 1852
rect 12548 1805 12582 1839
rect 12652 1818 12686 1852
rect 12736 1801 12770 1835
rect 12820 1818 12854 1852
rect 12904 1818 12938 1852
rect 13093 1809 13127 1843
rect 13177 1918 13211 1952
rect 13177 1824 13211 1858
rect 13796 1921 13830 1955
rect 13796 1831 13830 1865
rect 13880 1801 13914 1835
rect 14147 1813 14181 1847
rect 14248 1818 14282 1852
rect 14332 1801 14366 1835
rect 14416 1818 14450 1852
rect 14500 1805 14534 1839
rect 14604 1818 14638 1852
rect 14688 1801 14722 1835
rect 14772 1818 14806 1852
rect 14856 1818 14890 1852
rect 15045 1809 15079 1843
rect 15129 1918 15163 1952
rect 15129 1824 15163 1858
rect 15860 1921 15894 1955
rect 15860 1831 15894 1865
rect 15944 1801 15978 1835
rect 16211 1813 16245 1847
rect 16312 1818 16346 1852
rect 16396 1801 16430 1835
rect 16480 1818 16514 1852
rect 16564 1805 16598 1839
rect 16668 1818 16702 1852
rect 16752 1801 16786 1835
rect 16836 1818 16870 1852
rect 16920 1818 16954 1852
rect 17109 1809 17143 1843
rect 17193 1918 17227 1952
rect 17193 1824 17227 1858
<< psubdiff >>
rect 18971 43447 18995 43481
rect 19029 43447 19076 43481
rect 18955 41461 18979 41495
rect 19013 41461 19060 41495
rect 18963 39665 18987 39699
rect 19021 39665 19068 39699
rect 18977 38403 19001 38437
rect 19035 38403 19082 38437
rect 18989 37249 19013 37283
rect 19047 37249 19094 37283
rect 18997 36365 19021 36399
rect 19055 36365 19102 36399
rect 19021 34977 19045 35011
rect 19079 34977 19126 35011
rect 19021 32695 19045 32729
rect 19079 32695 19126 32729
rect 19025 30449 19049 30483
rect 19083 30449 19130 30483
rect 19017 28263 19041 28297
rect 19075 28263 19122 28297
rect 19021 26017 19045 26051
rect 19079 26017 19126 26051
rect 9447 22973 9481 22997
rect 9447 22892 9481 22939
rect 11693 22977 11727 23001
rect 11693 22896 11727 22943
rect 13879 22969 13913 22993
rect 13879 22888 13913 22935
rect 16125 22973 16159 22997
rect 16125 22892 16159 22939
rect 18407 22973 18441 22997
rect 18407 22892 18441 22939
rect 9719 17683 9753 17730
rect 9719 17625 9753 17649
rect 15510 17535 15544 17582
rect 15510 17477 15544 17501
rect 16296 17573 16330 17620
rect 16296 17515 16330 17539
rect 17162 17575 17196 17622
rect 17162 17517 17196 17541
rect 17940 17565 17974 17612
rect 17940 17507 17974 17531
rect 19056 17567 19090 17614
rect 19056 17509 19090 17533
rect 19922 17569 19956 17616
rect 19922 17511 19956 17535
rect 20692 17559 20726 17606
rect 20692 17501 20726 17525
rect 21670 17557 21704 17604
rect 21670 17499 21704 17523
rect 22178 17559 22212 17606
rect 22178 17501 22212 17525
rect 23310 17549 23344 17596
rect 23310 17491 23344 17515
rect 16275 16295 16309 16319
rect 4405 16187 4439 16211
rect 4405 16106 4439 16153
rect 9271 16191 9305 16215
rect 9271 16110 9305 16157
rect 16275 16214 16309 16261
rect 17407 16285 17441 16309
rect 17407 16204 17441 16251
rect 17915 16287 17949 16311
rect 17915 16206 17949 16253
rect 18893 16285 18927 16309
rect 18893 16204 18927 16251
rect 19663 16275 19697 16299
rect 19663 16194 19697 16241
rect 20529 16277 20563 16301
rect 20529 16196 20563 16243
rect 21645 16279 21679 16303
rect 21645 16198 21679 16245
rect 22423 16269 22457 16293
rect 22423 16188 22457 16235
rect 23289 16271 23323 16295
rect 23289 16190 23323 16237
rect 4505 15443 4539 15467
rect 4505 15362 4539 15409
rect 9371 15447 9405 15471
rect 9371 15366 9405 15413
rect 7281 15333 7315 15357
rect 7281 15252 7315 15299
rect 12147 15337 12181 15361
rect 12147 15256 12181 15303
rect 6239 14833 6273 14857
rect 6239 14752 6273 14799
rect 11105 14837 11139 14861
rect 11105 14756 11139 14803
rect 4415 14623 4449 14647
rect 4415 14542 4449 14589
rect 9281 14627 9315 14651
rect 9281 14546 9315 14593
rect 25445 14433 25479 14457
rect 25445 14352 25479 14399
rect 4515 13879 4549 13903
rect 4515 13798 4549 13845
rect 5761 13867 5795 13891
rect 5761 13786 5795 13833
rect 9379 13883 9413 13907
rect 8303 13851 8337 13875
rect 8303 13770 8337 13817
rect 9379 13802 9413 13849
rect 10627 13871 10661 13895
rect 10627 13790 10661 13837
rect 13169 13855 13203 13879
rect 13169 13774 13203 13821
rect 7279 13493 7313 13517
rect 7279 13412 7313 13459
rect 5885 13025 5919 13049
rect 12147 13497 12181 13521
rect 12147 13416 12181 13463
rect 4407 12955 4441 12979
rect 4407 12874 4441 12921
rect 5885 12944 5919 12991
rect 10751 13029 10785 13053
rect 9273 12959 9307 12983
rect 9273 12878 9307 12925
rect 10751 12948 10785 12995
rect 4507 12211 4541 12235
rect 4507 12130 4541 12177
rect 5881 12005 5915 12029
rect 9371 12215 9405 12239
rect 9371 12134 9405 12181
rect 5881 11924 5915 11971
rect 10747 12009 10781 12033
rect 10747 11928 10781 11975
rect 4417 11391 4451 11415
rect 4417 11310 4451 11357
rect 9283 11395 9317 11419
rect 9283 11314 9317 11361
rect 4515 10647 4549 10671
rect 4515 10566 4549 10613
rect 9381 10651 9415 10675
rect 9381 10570 9415 10617
rect 6407 6489 6441 6536
rect 6407 6431 6441 6455
rect 9957 5857 9991 5904
rect 9957 5799 9991 5823
rect 1775 5437 1809 5484
rect 1775 5379 1809 5403
rect 3909 5429 3943 5476
rect 3909 5371 3943 5395
rect 5859 5429 5893 5476
rect 5859 5371 5893 5395
rect 7861 5435 7895 5482
rect 7861 5377 7895 5401
rect 12017 5845 12051 5892
rect 12017 5787 12051 5811
rect 13975 5853 14009 5900
rect 13975 5795 14009 5819
rect 15971 5859 16005 5906
rect 15971 5801 16005 5825
rect 11547 4983 11581 5030
rect 11547 4925 11581 4949
rect 12257 4939 12291 4986
rect 12257 4881 12291 4905
rect 19159 5285 19193 5332
rect 19159 5227 19193 5251
rect 14257 4933 14291 4980
rect 14257 4875 14291 4899
rect 16281 4915 16315 4962
rect 16281 4857 16315 4881
rect 6023 3229 6057 3276
rect 6023 3171 6057 3195
rect 1745 2177 1779 2224
rect 1745 2119 1779 2143
rect 3815 2173 3849 2220
rect 3815 2115 3849 2139
rect 5771 2173 5805 2220
rect 5771 2115 5805 2139
rect 7769 2179 7803 2226
rect 7769 2121 7803 2145
rect 9725 2179 9759 2226
rect 9725 2121 9759 2145
rect 11713 2179 11747 2226
rect 11713 2121 11747 2145
rect 13667 2179 13701 2226
rect 13667 2121 13701 2145
rect 15729 2179 15763 2226
rect 15729 2121 15763 2145
<< nsubdiff >>
rect 18660 43447 18684 43481
rect 18718 43447 18777 43481
rect 18811 43447 18835 43481
rect 18644 41461 18668 41495
rect 18702 41461 18761 41495
rect 18795 41461 18819 41495
rect 18652 39665 18676 39699
rect 18710 39665 18769 39699
rect 18803 39665 18827 39699
rect 18666 38403 18690 38437
rect 18724 38403 18783 38437
rect 18817 38403 18841 38437
rect 18678 37249 18702 37283
rect 18736 37249 18795 37283
rect 18829 37249 18853 37283
rect 18686 36365 18710 36399
rect 18744 36365 18803 36399
rect 18837 36365 18861 36399
rect 18710 34977 18734 35011
rect 18768 34977 18827 35011
rect 18861 34977 18885 35011
rect 18710 32695 18734 32729
rect 18768 32695 18827 32729
rect 18861 32695 18885 32729
rect 18714 30449 18738 30483
rect 18772 30449 18831 30483
rect 18865 30449 18889 30483
rect 18706 28263 18730 28297
rect 18764 28263 18823 28297
rect 18857 28263 18881 28297
rect 18710 26017 18734 26051
rect 18768 26017 18827 26051
rect 18861 26017 18885 26051
rect 9447 23284 9481 23308
rect 9447 23191 9481 23250
rect 9447 23133 9481 23157
rect 11693 23288 11727 23312
rect 11693 23195 11727 23254
rect 11693 23137 11727 23161
rect 13879 23280 13913 23304
rect 13879 23187 13913 23246
rect 13879 23129 13913 23153
rect 16125 23284 16159 23308
rect 16125 23191 16159 23250
rect 16125 23133 16159 23157
rect 18407 23284 18441 23308
rect 18407 23191 18441 23250
rect 18407 23133 18441 23157
rect 9719 17465 9753 17489
rect 9719 17372 9753 17431
rect 16296 17355 16330 17379
rect 9719 17314 9753 17338
rect 15510 17317 15544 17341
rect 15510 17224 15544 17283
rect 15510 17166 15544 17190
rect 16296 17262 16330 17321
rect 16296 17204 16330 17228
rect 17162 17357 17196 17381
rect 17162 17264 17196 17323
rect 17162 17206 17196 17230
rect 17940 17347 17974 17371
rect 17940 17254 17974 17313
rect 17940 17196 17974 17220
rect 19056 17349 19090 17373
rect 19056 17256 19090 17315
rect 19056 17198 19090 17222
rect 19922 17351 19956 17375
rect 19922 17258 19956 17317
rect 19922 17200 19956 17224
rect 20692 17341 20726 17365
rect 20692 17248 20726 17307
rect 20692 17190 20726 17214
rect 21670 17339 21704 17363
rect 21670 17246 21704 17305
rect 21670 17188 21704 17212
rect 22178 17341 22212 17365
rect 22178 17248 22212 17307
rect 22178 17190 22212 17214
rect 23310 17331 23344 17355
rect 23310 17238 23344 17297
rect 23310 17180 23344 17204
rect 16275 16606 16309 16630
rect 4405 16498 4439 16522
rect 4405 16405 4439 16464
rect 4405 16347 4439 16371
rect 9271 16502 9305 16526
rect 9271 16409 9305 16468
rect 9271 16351 9305 16375
rect 16275 16513 16309 16572
rect 16275 16455 16309 16479
rect 17407 16596 17441 16620
rect 17407 16503 17441 16562
rect 17407 16445 17441 16469
rect 17915 16598 17949 16622
rect 17915 16505 17949 16564
rect 17915 16447 17949 16471
rect 18893 16596 18927 16620
rect 18893 16503 18927 16562
rect 18893 16445 18927 16469
rect 19663 16586 19697 16610
rect 19663 16493 19697 16552
rect 19663 16435 19697 16459
rect 20529 16588 20563 16612
rect 20529 16495 20563 16554
rect 20529 16437 20563 16461
rect 21645 16590 21679 16614
rect 21645 16497 21679 16556
rect 21645 16439 21679 16463
rect 22423 16580 22457 16604
rect 22423 16487 22457 16546
rect 22423 16429 22457 16453
rect 23289 16582 23323 16606
rect 23289 16489 23323 16548
rect 23289 16431 23323 16455
rect 4505 15754 4539 15778
rect 4505 15661 4539 15720
rect 4505 15603 4539 15627
rect 9371 15758 9405 15782
rect 7281 15644 7315 15668
rect 7281 15551 7315 15610
rect 9371 15665 9405 15724
rect 9371 15607 9405 15631
rect 7281 15493 7315 15517
rect 12147 15648 12181 15672
rect 12147 15555 12181 15614
rect 12147 15497 12181 15521
rect 4415 14934 4449 14958
rect 4415 14841 4449 14900
rect 4415 14783 4449 14807
rect 6239 15144 6273 15168
rect 6239 15051 6273 15110
rect 6239 14993 6273 15017
rect 9281 14938 9315 14962
rect 9281 14845 9315 14904
rect 9281 14787 9315 14811
rect 11105 15148 11139 15172
rect 11105 15055 11139 15114
rect 11105 14997 11139 15021
rect 25445 14744 25479 14768
rect 25445 14651 25479 14710
rect 25445 14593 25479 14617
rect 4515 14190 4549 14214
rect 4515 14097 4549 14156
rect 4515 14039 4549 14063
rect 5761 14178 5795 14202
rect 5761 14085 5795 14144
rect 5761 14027 5795 14051
rect 9379 14194 9413 14218
rect 8303 14162 8337 14186
rect 8303 14069 8337 14128
rect 9379 14101 9413 14160
rect 9379 14043 9413 14067
rect 8303 14011 8337 14035
rect 10627 14182 10661 14206
rect 10627 14089 10661 14148
rect 10627 14031 10661 14055
rect 13169 14166 13203 14190
rect 13169 14073 13203 14132
rect 13169 14015 13203 14039
rect 7279 13804 7313 13828
rect 7279 13711 7313 13770
rect 7279 13653 7313 13677
rect 12147 13808 12181 13832
rect 12147 13715 12181 13774
rect 12147 13657 12181 13681
rect 5885 13336 5919 13360
rect 4407 13266 4441 13290
rect 4407 13173 4441 13232
rect 4407 13115 4441 13139
rect 5885 13243 5919 13302
rect 5885 13185 5919 13209
rect 10751 13340 10785 13364
rect 9273 13270 9307 13294
rect 9273 13177 9307 13236
rect 9273 13119 9307 13143
rect 10751 13247 10785 13306
rect 10751 13189 10785 13213
rect 4507 12522 4541 12546
rect 4507 12429 4541 12488
rect 4507 12371 4541 12395
rect 9371 12526 9405 12550
rect 9371 12433 9405 12492
rect 9371 12375 9405 12399
rect 5881 12316 5915 12340
rect 5881 12223 5915 12282
rect 5881 12165 5915 12189
rect 10747 12320 10781 12344
rect 10747 12227 10781 12286
rect 10747 12169 10781 12193
rect 4417 11702 4451 11726
rect 4417 11609 4451 11668
rect 4417 11551 4451 11575
rect 9283 11706 9317 11730
rect 9283 11613 9317 11672
rect 9283 11555 9317 11579
rect 4515 10958 4549 10982
rect 4515 10865 4549 10924
rect 4515 10807 4549 10831
rect 9381 10962 9415 10986
rect 9381 10869 9415 10928
rect 9381 10811 9415 10835
rect 6407 6271 6441 6295
rect 6407 6178 6441 6237
rect 6407 6120 6441 6144
rect 9957 5639 9991 5663
rect 9957 5546 9991 5605
rect 1775 5219 1809 5243
rect 1775 5126 1809 5185
rect 1775 5068 1809 5092
rect 3909 5211 3943 5235
rect 3909 5118 3943 5177
rect 3909 5060 3943 5084
rect 5859 5211 5893 5235
rect 5859 5118 5893 5177
rect 5859 5060 5893 5084
rect 7861 5217 7895 5241
rect 7861 5124 7895 5183
rect 7861 5066 7895 5090
rect 9957 5488 9991 5512
rect 12017 5627 12051 5651
rect 12017 5534 12051 5593
rect 12017 5476 12051 5500
rect 13975 5635 14009 5659
rect 13975 5542 14009 5601
rect 13975 5484 14009 5508
rect 15971 5641 16005 5665
rect 15971 5548 16005 5607
rect 15971 5490 16005 5514
rect 11547 4765 11581 4789
rect 11547 4672 11581 4731
rect 11547 4614 11581 4638
rect 12257 4721 12291 4745
rect 12257 4628 12291 4687
rect 12257 4570 12291 4594
rect 14257 4715 14291 4739
rect 14257 4622 14291 4681
rect 14257 4564 14291 4588
rect 16281 4697 16315 4721
rect 16281 4604 16315 4663
rect 16281 4546 16315 4570
rect 19159 5067 19193 5091
rect 19159 4974 19193 5033
rect 19159 4916 19193 4940
rect 6023 3011 6057 3035
rect 6023 2918 6057 2977
rect 6023 2860 6057 2884
rect 1745 1959 1779 1983
rect 1745 1866 1779 1925
rect 1745 1808 1779 1832
rect 3815 1955 3849 1979
rect 3815 1862 3849 1921
rect 3815 1804 3849 1828
rect 5771 1955 5805 1979
rect 5771 1862 5805 1921
rect 5771 1804 5805 1828
rect 7769 1961 7803 1985
rect 7769 1868 7803 1927
rect 7769 1810 7803 1834
rect 9725 1961 9759 1985
rect 9725 1868 9759 1927
rect 9725 1810 9759 1834
rect 11713 1961 11747 1985
rect 11713 1868 11747 1927
rect 11713 1810 11747 1834
rect 13667 1961 13701 1985
rect 13667 1868 13701 1927
rect 13667 1810 13701 1834
rect 15729 1961 15763 1985
rect 15729 1868 15763 1927
rect 15729 1810 15763 1834
<< psubdiffcont >>
rect 18995 43447 19029 43481
rect 18979 41461 19013 41495
rect 18987 39665 19021 39699
rect 19001 38403 19035 38437
rect 19013 37249 19047 37283
rect 19021 36365 19055 36399
rect 19045 34977 19079 35011
rect 19045 32695 19079 32729
rect 19049 30449 19083 30483
rect 19041 28263 19075 28297
rect 19045 26017 19079 26051
rect 9447 22939 9481 22973
rect 11693 22943 11727 22977
rect 13879 22935 13913 22969
rect 16125 22939 16159 22973
rect 18407 22939 18441 22973
rect 9719 17649 9753 17683
rect 15510 17501 15544 17535
rect 16296 17539 16330 17573
rect 17162 17541 17196 17575
rect 17940 17531 17974 17565
rect 19056 17533 19090 17567
rect 19922 17535 19956 17569
rect 20692 17525 20726 17559
rect 21670 17523 21704 17557
rect 22178 17525 22212 17559
rect 23310 17515 23344 17549
rect 16275 16261 16309 16295
rect 4405 16153 4439 16187
rect 9271 16157 9305 16191
rect 17407 16251 17441 16285
rect 17915 16253 17949 16287
rect 18893 16251 18927 16285
rect 19663 16241 19697 16275
rect 20529 16243 20563 16277
rect 21645 16245 21679 16279
rect 22423 16235 22457 16269
rect 23289 16237 23323 16271
rect 4505 15409 4539 15443
rect 9371 15413 9405 15447
rect 7281 15299 7315 15333
rect 12147 15303 12181 15337
rect 6239 14799 6273 14833
rect 11105 14803 11139 14837
rect 4415 14589 4449 14623
rect 9281 14593 9315 14627
rect 25445 14399 25479 14433
rect 4515 13845 4549 13879
rect 5761 13833 5795 13867
rect 8303 13817 8337 13851
rect 9379 13849 9413 13883
rect 10627 13837 10661 13871
rect 13169 13821 13203 13855
rect 7279 13459 7313 13493
rect 5885 12991 5919 13025
rect 12147 13463 12181 13497
rect 4407 12921 4441 12955
rect 10751 12995 10785 13029
rect 9273 12925 9307 12959
rect 4507 12177 4541 12211
rect 9371 12181 9405 12215
rect 5881 11971 5915 12005
rect 10747 11975 10781 12009
rect 4417 11357 4451 11391
rect 9283 11361 9317 11395
rect 4515 10613 4549 10647
rect 9381 10617 9415 10651
rect 6407 6455 6441 6489
rect 9957 5823 9991 5857
rect 1775 5403 1809 5437
rect 3909 5395 3943 5429
rect 5859 5395 5893 5429
rect 7861 5401 7895 5435
rect 12017 5811 12051 5845
rect 13975 5819 14009 5853
rect 15971 5825 16005 5859
rect 11547 4949 11581 4983
rect 12257 4905 12291 4939
rect 19159 5251 19193 5285
rect 14257 4899 14291 4933
rect 16281 4881 16315 4915
rect 6023 3195 6057 3229
rect 1745 2143 1779 2177
rect 3815 2139 3849 2173
rect 5771 2139 5805 2173
rect 7769 2145 7803 2179
rect 9725 2145 9759 2179
rect 11713 2145 11747 2179
rect 13667 2145 13701 2179
rect 15729 2145 15763 2179
<< nsubdiffcont >>
rect 18684 43447 18718 43481
rect 18777 43447 18811 43481
rect 18668 41461 18702 41495
rect 18761 41461 18795 41495
rect 18676 39665 18710 39699
rect 18769 39665 18803 39699
rect 18690 38403 18724 38437
rect 18783 38403 18817 38437
rect 18702 37249 18736 37283
rect 18795 37249 18829 37283
rect 18710 36365 18744 36399
rect 18803 36365 18837 36399
rect 18734 34977 18768 35011
rect 18827 34977 18861 35011
rect 18734 32695 18768 32729
rect 18827 32695 18861 32729
rect 18738 30449 18772 30483
rect 18831 30449 18865 30483
rect 18730 28263 18764 28297
rect 18823 28263 18857 28297
rect 18734 26017 18768 26051
rect 18827 26017 18861 26051
rect 9447 23250 9481 23284
rect 9447 23157 9481 23191
rect 11693 23254 11727 23288
rect 11693 23161 11727 23195
rect 13879 23246 13913 23280
rect 13879 23153 13913 23187
rect 16125 23250 16159 23284
rect 16125 23157 16159 23191
rect 18407 23250 18441 23284
rect 18407 23157 18441 23191
rect 9719 17431 9753 17465
rect 9719 17338 9753 17372
rect 15510 17283 15544 17317
rect 15510 17190 15544 17224
rect 16296 17321 16330 17355
rect 16296 17228 16330 17262
rect 17162 17323 17196 17357
rect 17162 17230 17196 17264
rect 17940 17313 17974 17347
rect 17940 17220 17974 17254
rect 19056 17315 19090 17349
rect 19056 17222 19090 17256
rect 19922 17317 19956 17351
rect 19922 17224 19956 17258
rect 20692 17307 20726 17341
rect 20692 17214 20726 17248
rect 21670 17305 21704 17339
rect 21670 17212 21704 17246
rect 22178 17307 22212 17341
rect 22178 17214 22212 17248
rect 23310 17297 23344 17331
rect 23310 17204 23344 17238
rect 16275 16572 16309 16606
rect 4405 16464 4439 16498
rect 4405 16371 4439 16405
rect 9271 16468 9305 16502
rect 9271 16375 9305 16409
rect 16275 16479 16309 16513
rect 17407 16562 17441 16596
rect 17407 16469 17441 16503
rect 17915 16564 17949 16598
rect 17915 16471 17949 16505
rect 18893 16562 18927 16596
rect 18893 16469 18927 16503
rect 19663 16552 19697 16586
rect 19663 16459 19697 16493
rect 20529 16554 20563 16588
rect 20529 16461 20563 16495
rect 21645 16556 21679 16590
rect 21645 16463 21679 16497
rect 22423 16546 22457 16580
rect 22423 16453 22457 16487
rect 23289 16548 23323 16582
rect 23289 16455 23323 16489
rect 4505 15720 4539 15754
rect 4505 15627 4539 15661
rect 9371 15724 9405 15758
rect 7281 15610 7315 15644
rect 9371 15631 9405 15665
rect 7281 15517 7315 15551
rect 12147 15614 12181 15648
rect 12147 15521 12181 15555
rect 4415 14900 4449 14934
rect 4415 14807 4449 14841
rect 6239 15110 6273 15144
rect 6239 15017 6273 15051
rect 9281 14904 9315 14938
rect 9281 14811 9315 14845
rect 11105 15114 11139 15148
rect 11105 15021 11139 15055
rect 25445 14710 25479 14744
rect 25445 14617 25479 14651
rect 4515 14156 4549 14190
rect 4515 14063 4549 14097
rect 5761 14144 5795 14178
rect 5761 14051 5795 14085
rect 8303 14128 8337 14162
rect 8303 14035 8337 14069
rect 9379 14160 9413 14194
rect 9379 14067 9413 14101
rect 10627 14148 10661 14182
rect 10627 14055 10661 14089
rect 13169 14132 13203 14166
rect 13169 14039 13203 14073
rect 7279 13770 7313 13804
rect 7279 13677 7313 13711
rect 12147 13774 12181 13808
rect 12147 13681 12181 13715
rect 4407 13232 4441 13266
rect 4407 13139 4441 13173
rect 5885 13302 5919 13336
rect 5885 13209 5919 13243
rect 9273 13236 9307 13270
rect 9273 13143 9307 13177
rect 10751 13306 10785 13340
rect 10751 13213 10785 13247
rect 4507 12488 4541 12522
rect 4507 12395 4541 12429
rect 9371 12492 9405 12526
rect 9371 12399 9405 12433
rect 5881 12282 5915 12316
rect 5881 12189 5915 12223
rect 10747 12286 10781 12320
rect 10747 12193 10781 12227
rect 4417 11668 4451 11702
rect 4417 11575 4451 11609
rect 9283 11672 9317 11706
rect 9283 11579 9317 11613
rect 4515 10924 4549 10958
rect 4515 10831 4549 10865
rect 9381 10928 9415 10962
rect 9381 10835 9415 10869
rect 6407 6237 6441 6271
rect 6407 6144 6441 6178
rect 9957 5605 9991 5639
rect 1775 5185 1809 5219
rect 1775 5092 1809 5126
rect 9957 5512 9991 5546
rect 3909 5177 3943 5211
rect 3909 5084 3943 5118
rect 5859 5177 5893 5211
rect 5859 5084 5893 5118
rect 7861 5183 7895 5217
rect 7861 5090 7895 5124
rect 12017 5593 12051 5627
rect 12017 5500 12051 5534
rect 13975 5601 14009 5635
rect 13975 5508 14009 5542
rect 15971 5607 16005 5641
rect 15971 5514 16005 5548
rect 11547 4731 11581 4765
rect 11547 4638 11581 4672
rect 12257 4687 12291 4721
rect 12257 4594 12291 4628
rect 14257 4681 14291 4715
rect 14257 4588 14291 4622
rect 16281 4663 16315 4697
rect 16281 4570 16315 4604
rect 19159 5033 19193 5067
rect 19159 4940 19193 4974
rect 6023 2977 6057 3011
rect 6023 2884 6057 2918
rect 1745 1925 1779 1959
rect 1745 1832 1779 1866
rect 3815 1921 3849 1955
rect 3815 1828 3849 1862
rect 5771 1921 5805 1955
rect 5771 1828 5805 1862
rect 7769 1927 7803 1961
rect 7769 1834 7803 1868
rect 9725 1927 9759 1961
rect 9725 1834 9759 1868
rect 11713 1927 11747 1961
rect 11713 1834 11747 1868
rect 13667 1927 13701 1961
rect 13667 1834 13701 1868
rect 15729 1927 15763 1961
rect 15729 1834 15763 1868
<< poly >>
rect 18617 43300 18643 43330
rect 18843 43300 18963 43330
rect 19093 43300 19119 43330
rect 18875 43246 18941 43300
rect 18617 43216 18643 43246
rect 18843 43216 18963 43246
rect 19093 43216 19119 43246
rect 18875 43162 18941 43216
rect 18617 43132 18643 43162
rect 18843 43132 18963 43162
rect 19093 43132 19119 43162
rect 18875 43078 18941 43132
rect 18617 43048 18643 43078
rect 18843 43048 18963 43078
rect 19093 43048 19119 43078
rect 18875 43037 18941 43048
rect 18875 43003 18891 43037
rect 18925 43003 18941 43037
rect 18875 42994 18941 43003
rect 18617 42964 18643 42994
rect 18843 42964 18963 42994
rect 19093 42964 19119 42994
rect 18875 42910 18941 42964
rect 18617 42880 18643 42910
rect 18843 42880 18963 42910
rect 19093 42880 19119 42910
rect 18875 42870 18941 42880
rect 18875 42836 18891 42870
rect 18925 42836 18941 42870
rect 18875 42826 18941 42836
rect 18617 42796 18643 42826
rect 18843 42796 18963 42826
rect 19093 42796 19119 42826
rect 18875 42742 18941 42796
rect 18617 42712 18643 42742
rect 18843 42712 18963 42742
rect 19093 42712 19119 42742
rect 18875 42702 18941 42712
rect 18875 42668 18891 42702
rect 18925 42668 18941 42702
rect 18875 42658 18941 42668
rect 18617 42628 18643 42658
rect 18843 42628 18963 42658
rect 19093 42628 19119 42658
rect 18875 42574 18941 42628
rect 18617 42544 18643 42574
rect 18843 42544 18963 42574
rect 19093 42544 19119 42574
rect 18875 42535 18941 42544
rect 18875 42501 18891 42535
rect 18925 42501 18941 42535
rect 18875 42490 18941 42501
rect 18617 42460 18643 42490
rect 18843 42460 18963 42490
rect 19093 42460 19119 42490
rect 18875 42406 18941 42460
rect 18617 42376 18643 42406
rect 18843 42376 18963 42406
rect 19093 42376 19119 42406
rect 18875 42366 18941 42376
rect 18875 42332 18891 42366
rect 18925 42332 18941 42366
rect 18875 42322 18941 42332
rect 18617 42292 18643 42322
rect 18843 42292 18963 42322
rect 19093 42292 19119 42322
rect 18875 42238 18941 42292
rect 18617 42208 18643 42238
rect 18843 42208 18963 42238
rect 19093 42208 19119 42238
rect 18875 42198 18941 42208
rect 18875 42164 18891 42198
rect 18925 42164 18941 42198
rect 18875 42154 18941 42164
rect 18617 42124 18643 42154
rect 18843 42124 18963 42154
rect 19093 42124 19119 42154
rect 18875 42070 18941 42124
rect 18617 42040 18643 42070
rect 18843 42040 18963 42070
rect 19093 42040 19119 42070
rect 18875 42024 18941 42040
rect 18875 41990 18891 42024
rect 18925 41990 18941 42024
rect 18875 41974 18941 41990
rect 18601 41272 18627 41302
rect 18827 41272 18947 41302
rect 19077 41272 19103 41302
rect 18859 41262 18925 41272
rect 18859 41228 18875 41262
rect 18909 41228 18925 41262
rect 18859 41218 18925 41228
rect 18601 41188 18627 41218
rect 18827 41188 18947 41218
rect 19077 41188 19103 41218
rect 18859 41178 18925 41188
rect 18859 41144 18875 41178
rect 18909 41144 18925 41178
rect 18859 41134 18925 41144
rect 18601 41104 18627 41134
rect 18827 41104 18947 41134
rect 19077 41104 19103 41134
rect 18859 41094 18925 41104
rect 18859 41060 18875 41094
rect 18909 41060 18925 41094
rect 18859 41050 18925 41060
rect 18601 41020 18627 41050
rect 18827 41020 18947 41050
rect 19077 41020 19103 41050
rect 18859 41010 18925 41020
rect 18859 40976 18875 41010
rect 18909 40976 18925 41010
rect 18859 40966 18925 40976
rect 18601 40936 18627 40966
rect 18827 40936 18947 40966
rect 19077 40936 19103 40966
rect 18859 40926 18925 40936
rect 18859 40892 18875 40926
rect 18909 40892 18925 40926
rect 18859 40882 18925 40892
rect 18601 40852 18627 40882
rect 18827 40852 18947 40882
rect 19077 40852 19103 40882
rect 18859 40842 18925 40852
rect 18859 40808 18875 40842
rect 18909 40808 18925 40842
rect 18859 40798 18925 40808
rect 18601 40768 18627 40798
rect 18827 40768 18947 40798
rect 19077 40768 19103 40798
rect 18859 40758 18925 40768
rect 18859 40724 18875 40758
rect 18909 40724 18925 40758
rect 18859 40714 18925 40724
rect 18601 40684 18627 40714
rect 18827 40684 18947 40714
rect 19077 40684 19103 40714
rect 18859 40674 18925 40684
rect 18859 40640 18875 40674
rect 18909 40640 18925 40674
rect 18859 40630 18925 40640
rect 18601 40600 18627 40630
rect 18827 40600 18947 40630
rect 19077 40600 19103 40630
rect 18859 40590 18925 40600
rect 18859 40556 18875 40590
rect 18909 40556 18925 40590
rect 18859 40546 18925 40556
rect 18601 40516 18627 40546
rect 18827 40516 18947 40546
rect 19077 40516 19103 40546
rect 18859 40506 18925 40516
rect 18859 40472 18875 40506
rect 18909 40472 18925 40506
rect 18859 40462 18925 40472
rect 18601 40432 18627 40462
rect 18827 40432 18947 40462
rect 19077 40432 19103 40462
rect 18859 40422 18925 40432
rect 18859 40388 18875 40422
rect 18909 40388 18925 40422
rect 18859 40378 18925 40388
rect 18601 40348 18627 40378
rect 18827 40348 18947 40378
rect 19077 40348 19103 40378
rect 18609 39508 18635 39538
rect 18835 39508 18955 39538
rect 19085 39508 19111 39538
rect 18867 39498 18933 39508
rect 18867 39464 18883 39498
rect 18917 39464 18933 39498
rect 18867 39454 18933 39464
rect 18609 39424 18635 39454
rect 18835 39424 18955 39454
rect 19085 39424 19111 39454
rect 18867 39414 18933 39424
rect 18867 39380 18883 39414
rect 18917 39380 18933 39414
rect 18867 39370 18933 39380
rect 18609 39340 18635 39370
rect 18835 39340 18955 39370
rect 19085 39340 19111 39370
rect 18867 39330 18933 39340
rect 18867 39296 18883 39330
rect 18917 39296 18933 39330
rect 18867 39286 18933 39296
rect 18609 39256 18635 39286
rect 18835 39256 18955 39286
rect 19085 39256 19111 39286
rect 18867 39246 18933 39256
rect 18867 39212 18883 39246
rect 18917 39212 18933 39246
rect 18867 39202 18933 39212
rect 18609 39172 18635 39202
rect 18835 39172 18955 39202
rect 19085 39172 19111 39202
rect 18867 39162 18933 39172
rect 18867 39128 18883 39162
rect 18917 39128 18933 39162
rect 18867 39118 18933 39128
rect 18609 39088 18635 39118
rect 18835 39088 18955 39118
rect 19085 39088 19111 39118
rect 18867 39078 18933 39088
rect 18867 39044 18883 39078
rect 18917 39044 18933 39078
rect 18867 39034 18933 39044
rect 18609 39004 18635 39034
rect 18835 39004 18955 39034
rect 19085 39004 19111 39034
rect 18867 38994 18933 39004
rect 18867 38960 18883 38994
rect 18917 38960 18933 38994
rect 18867 38950 18933 38960
rect 18609 38920 18635 38950
rect 18835 38920 18955 38950
rect 19085 38920 19111 38950
rect 18623 38263 18649 38293
rect 18849 38263 18969 38293
rect 19099 38263 19125 38293
rect 18881 38237 18947 38263
rect 18881 38209 18897 38237
rect 18623 38179 18649 38209
rect 18849 38203 18897 38209
rect 18931 38209 18947 38237
rect 18931 38203 18969 38209
rect 18849 38179 18969 38203
rect 19099 38179 19125 38209
rect 18881 38153 18947 38179
rect 18881 38125 18897 38153
rect 18623 38095 18649 38125
rect 18849 38119 18897 38125
rect 18931 38125 18947 38153
rect 18931 38119 18969 38125
rect 18849 38095 18969 38119
rect 19099 38095 19125 38125
rect 18881 38069 18947 38095
rect 18881 38041 18897 38069
rect 18623 38011 18649 38041
rect 18849 38035 18897 38041
rect 18931 38041 18947 38069
rect 18931 38035 18969 38041
rect 18849 38011 18969 38035
rect 19099 38011 19125 38041
rect 18881 37957 18947 38011
rect 18623 37927 18649 37957
rect 18849 37927 18969 37957
rect 19099 37927 19125 37957
rect 18881 37873 18947 37927
rect 18623 37843 18649 37873
rect 18849 37843 18969 37873
rect 19099 37843 19125 37873
rect 18881 37801 18947 37843
rect 18881 37767 18897 37801
rect 18931 37767 18947 37801
rect 18881 37751 18947 37767
rect 18635 37105 18661 37135
rect 18861 37105 18981 37135
rect 19111 37105 19137 37135
rect 18893 37095 18959 37105
rect 18893 37061 18909 37095
rect 18943 37061 18959 37095
rect 18893 37051 18959 37061
rect 18635 37021 18661 37051
rect 18861 37021 18981 37051
rect 19111 37021 19137 37051
rect 18893 37011 18959 37021
rect 18893 36977 18909 37011
rect 18943 36977 18959 37011
rect 18893 36967 18959 36977
rect 18635 36937 18661 36967
rect 18861 36937 18981 36967
rect 19111 36937 19137 36967
rect 18893 36927 18959 36937
rect 18893 36893 18909 36927
rect 18943 36893 18959 36927
rect 18893 36883 18959 36893
rect 18635 36853 18661 36883
rect 18861 36853 18981 36883
rect 19111 36853 19137 36883
rect 18893 36835 18959 36853
rect 18893 36801 18909 36835
rect 18943 36801 18959 36835
rect 18893 36785 18959 36801
rect 18643 36225 18669 36255
rect 18869 36225 18989 36255
rect 19119 36225 19145 36255
rect 18901 36171 18967 36225
rect 18643 36141 18669 36171
rect 18869 36141 18989 36171
rect 19119 36141 19145 36171
rect 18901 36131 18967 36141
rect 18901 36097 18917 36131
rect 18951 36097 18967 36131
rect 18901 36081 18967 36097
rect 18667 34839 18693 34869
rect 18893 34849 19013 34869
rect 18893 34839 18941 34849
rect 18925 34815 18941 34839
rect 18975 34839 19013 34849
rect 19143 34839 19169 34869
rect 18975 34815 18991 34839
rect 18925 34805 18991 34815
rect 18667 34742 18693 34772
rect 18821 34763 18887 34772
rect 19020 34763 19059 34774
rect 18821 34744 19059 34763
rect 19143 34744 19169 34774
rect 18821 34742 19044 34744
rect 18857 34733 19044 34742
rect 18925 34588 18991 34733
rect 18925 34584 18941 34588
rect 18667 34554 18693 34584
rect 18893 34554 18941 34584
rect 18975 34586 18991 34588
rect 18975 34556 19013 34586
rect 19143 34556 19169 34586
rect 18975 34554 18991 34556
rect 18925 34544 18991 34554
rect 18925 34500 19013 34502
rect 18667 34470 18693 34500
rect 18893 34472 19013 34500
rect 19143 34472 19169 34502
rect 18893 34470 18991 34472
rect 18925 34404 18991 34470
rect 18925 34370 18941 34404
rect 18975 34370 18991 34404
rect 18925 34360 18991 34370
rect 18809 34330 18875 34340
rect 18809 34296 18825 34330
rect 18859 34312 18875 34330
rect 18859 34296 19059 34312
rect 18809 34289 19059 34296
rect 18667 34259 18693 34289
rect 18777 34282 19059 34289
rect 19143 34282 19169 34312
rect 18777 34259 18875 34282
rect 18815 34194 18869 34210
rect 18815 34175 18825 34194
rect 18667 34145 18693 34175
rect 18777 34160 18825 34175
rect 18859 34160 18869 34194
rect 18777 34145 18869 34160
rect 18815 34144 18869 34145
rect 18911 34187 19071 34217
rect 19143 34187 19169 34217
rect 18911 34102 18941 34187
rect 18875 34092 18941 34102
rect 18875 34091 18891 34092
rect 18667 34061 18693 34091
rect 18777 34061 18891 34091
rect 18875 34058 18891 34061
rect 18925 34058 18941 34092
rect 18983 34135 19049 34145
rect 18983 34101 18999 34135
rect 19033 34111 19049 34135
rect 19033 34101 19071 34111
rect 18983 34081 19071 34101
rect 19143 34081 19169 34111
rect 18875 34048 18941 34058
rect 18970 33996 19015 34010
rect 18667 33966 18693 33996
rect 18843 33980 19015 33996
rect 19143 33980 19169 34010
rect 18843 33966 19000 33980
rect 18881 33956 18935 33966
rect 18881 33922 18891 33956
rect 18925 33922 18935 33956
rect 18881 33906 18935 33922
rect 18977 33892 19031 33908
rect 18977 33864 18987 33892
rect 18667 33834 18693 33864
rect 18777 33858 18987 33864
rect 19021 33891 19031 33892
rect 19021 33861 19059 33891
rect 19143 33861 19169 33891
rect 19021 33858 19031 33861
rect 18777 33834 19031 33858
rect 18809 33782 18875 33792
rect 18809 33761 18825 33782
rect 18667 33731 18693 33761
rect 18777 33748 18825 33761
rect 18859 33748 18875 33782
rect 18777 33731 18875 33748
rect 18917 33762 19071 33792
rect 19143 33762 19169 33792
rect 18917 33689 18947 33762
rect 18893 33673 18947 33689
rect 18893 33666 18903 33673
rect 18667 33636 18693 33666
rect 18777 33639 18903 33666
rect 18937 33639 18947 33673
rect 18989 33693 19043 33709
rect 18989 33659 18999 33693
rect 19033 33663 19071 33693
rect 19143 33663 19169 33693
rect 19033 33659 19043 33663
rect 18989 33643 19043 33659
rect 18777 33636 18947 33639
rect 18893 33623 18947 33636
rect 18667 33551 18693 33581
rect 18777 33551 19059 33581
rect 19143 33551 19169 33581
rect 18857 33530 18923 33551
rect 18857 33496 18873 33530
rect 18907 33496 18923 33530
rect 18857 33486 18923 33496
rect 18673 33363 18699 33393
rect 18827 33368 19059 33393
rect 18827 33363 18926 33368
rect 18916 33334 18926 33363
rect 18960 33363 19059 33368
rect 19143 33363 19169 33393
rect 18960 33334 18970 33363
rect 18916 33318 18970 33334
rect 18673 33279 18699 33309
rect 18827 33279 18872 33309
rect 18842 33276 18872 33279
rect 19014 33279 19059 33309
rect 19143 33279 19169 33309
rect 19014 33276 19044 33279
rect 18842 33266 19044 33276
rect 18842 33246 18941 33266
rect 18925 33232 18941 33246
rect 18975 33246 19044 33266
rect 18975 33232 18991 33246
rect 18925 33222 18991 33232
rect 18667 32557 18693 32587
rect 18893 32567 19013 32587
rect 18893 32557 18941 32567
rect 18925 32533 18941 32557
rect 18975 32557 19013 32567
rect 19143 32557 19169 32587
rect 18975 32533 18991 32557
rect 18925 32523 18991 32533
rect 18667 32460 18693 32490
rect 18821 32481 18887 32490
rect 19020 32481 19059 32492
rect 18821 32462 19059 32481
rect 19143 32462 19169 32492
rect 18821 32460 19044 32462
rect 18857 32451 19044 32460
rect 18925 32306 18991 32451
rect 18925 32302 18941 32306
rect 18667 32272 18693 32302
rect 18893 32272 18941 32302
rect 18975 32304 18991 32306
rect 18975 32274 19013 32304
rect 19143 32274 19169 32304
rect 18975 32272 18991 32274
rect 18925 32262 18991 32272
rect 18925 32218 19013 32220
rect 18667 32188 18693 32218
rect 18893 32190 19013 32218
rect 19143 32190 19169 32220
rect 18893 32188 18991 32190
rect 18925 32122 18991 32188
rect 18925 32088 18941 32122
rect 18975 32088 18991 32122
rect 18925 32078 18991 32088
rect 18809 32048 18875 32058
rect 18809 32014 18825 32048
rect 18859 32030 18875 32048
rect 18859 32014 19059 32030
rect 18809 32007 19059 32014
rect 18667 31977 18693 32007
rect 18777 32000 19059 32007
rect 19143 32000 19169 32030
rect 18777 31977 18875 32000
rect 18815 31912 18869 31928
rect 18815 31893 18825 31912
rect 18667 31863 18693 31893
rect 18777 31878 18825 31893
rect 18859 31878 18869 31912
rect 18777 31863 18869 31878
rect 18815 31862 18869 31863
rect 18911 31905 19071 31935
rect 19143 31905 19169 31935
rect 18911 31820 18941 31905
rect 18875 31810 18941 31820
rect 18875 31809 18891 31810
rect 18667 31779 18693 31809
rect 18777 31779 18891 31809
rect 18875 31776 18891 31779
rect 18925 31776 18941 31810
rect 18983 31853 19049 31863
rect 18983 31819 18999 31853
rect 19033 31829 19049 31853
rect 19033 31819 19071 31829
rect 18983 31799 19071 31819
rect 19143 31799 19169 31829
rect 18875 31766 18941 31776
rect 18970 31714 19015 31728
rect 18667 31684 18693 31714
rect 18843 31698 19015 31714
rect 19143 31698 19169 31728
rect 18843 31684 19000 31698
rect 18881 31674 18935 31684
rect 18881 31640 18891 31674
rect 18925 31640 18935 31674
rect 18881 31624 18935 31640
rect 18977 31610 19031 31626
rect 18977 31582 18987 31610
rect 18667 31552 18693 31582
rect 18777 31576 18987 31582
rect 19021 31609 19031 31610
rect 19021 31579 19059 31609
rect 19143 31579 19169 31609
rect 19021 31576 19031 31579
rect 18777 31552 19031 31576
rect 18809 31500 18875 31510
rect 18809 31479 18825 31500
rect 18667 31449 18693 31479
rect 18777 31466 18825 31479
rect 18859 31466 18875 31500
rect 18777 31449 18875 31466
rect 18917 31480 19071 31510
rect 19143 31480 19169 31510
rect 18917 31407 18947 31480
rect 18893 31391 18947 31407
rect 18893 31384 18903 31391
rect 18667 31354 18693 31384
rect 18777 31357 18903 31384
rect 18937 31357 18947 31391
rect 18989 31411 19043 31427
rect 18989 31377 18999 31411
rect 19033 31381 19071 31411
rect 19143 31381 19169 31411
rect 19033 31377 19043 31381
rect 18989 31361 19043 31377
rect 18777 31354 18947 31357
rect 18893 31341 18947 31354
rect 18667 31269 18693 31299
rect 18777 31269 19059 31299
rect 19143 31269 19169 31299
rect 18857 31248 18923 31269
rect 18857 31214 18873 31248
rect 18907 31214 18923 31248
rect 18857 31204 18923 31214
rect 18673 31081 18699 31111
rect 18827 31086 19059 31111
rect 18827 31081 18926 31086
rect 18916 31052 18926 31081
rect 18960 31081 19059 31086
rect 19143 31081 19169 31111
rect 18960 31052 18970 31081
rect 18916 31036 18970 31052
rect 18673 30997 18699 31027
rect 18827 30997 18872 31027
rect 18842 30994 18872 30997
rect 19014 30997 19059 31027
rect 19143 30997 19169 31027
rect 19014 30994 19044 30997
rect 18842 30984 19044 30994
rect 18842 30964 18941 30984
rect 18925 30950 18941 30964
rect 18975 30964 19044 30984
rect 18975 30950 18991 30964
rect 18925 30940 18991 30950
rect 18671 30311 18697 30341
rect 18897 30321 19017 30341
rect 18897 30311 18945 30321
rect 18929 30287 18945 30311
rect 18979 30311 19017 30321
rect 19147 30311 19173 30341
rect 18979 30287 18995 30311
rect 18929 30277 18995 30287
rect 18671 30214 18697 30244
rect 18825 30235 18891 30244
rect 19024 30235 19063 30246
rect 18825 30216 19063 30235
rect 19147 30216 19173 30246
rect 18825 30214 19048 30216
rect 18861 30205 19048 30214
rect 18929 30060 18995 30205
rect 18929 30056 18945 30060
rect 18671 30026 18697 30056
rect 18897 30026 18945 30056
rect 18979 30058 18995 30060
rect 18979 30028 19017 30058
rect 19147 30028 19173 30058
rect 18979 30026 18995 30028
rect 18929 30016 18995 30026
rect 18929 29972 19017 29974
rect 18671 29942 18697 29972
rect 18897 29944 19017 29972
rect 19147 29944 19173 29974
rect 18897 29942 18995 29944
rect 18929 29876 18995 29942
rect 18929 29842 18945 29876
rect 18979 29842 18995 29876
rect 18929 29832 18995 29842
rect 18813 29802 18879 29812
rect 18813 29768 18829 29802
rect 18863 29784 18879 29802
rect 18863 29768 19063 29784
rect 18813 29761 19063 29768
rect 18671 29731 18697 29761
rect 18781 29754 19063 29761
rect 19147 29754 19173 29784
rect 18781 29731 18879 29754
rect 18819 29666 18873 29682
rect 18819 29647 18829 29666
rect 18671 29617 18697 29647
rect 18781 29632 18829 29647
rect 18863 29632 18873 29666
rect 18781 29617 18873 29632
rect 18819 29616 18873 29617
rect 18915 29659 19075 29689
rect 19147 29659 19173 29689
rect 18915 29574 18945 29659
rect 18879 29564 18945 29574
rect 18879 29563 18895 29564
rect 18671 29533 18697 29563
rect 18781 29533 18895 29563
rect 18879 29530 18895 29533
rect 18929 29530 18945 29564
rect 18987 29607 19053 29617
rect 18987 29573 19003 29607
rect 19037 29583 19053 29607
rect 19037 29573 19075 29583
rect 18987 29553 19075 29573
rect 19147 29553 19173 29583
rect 18879 29520 18945 29530
rect 18974 29468 19019 29482
rect 18671 29438 18697 29468
rect 18847 29452 19019 29468
rect 19147 29452 19173 29482
rect 18847 29438 19004 29452
rect 18885 29428 18939 29438
rect 18885 29394 18895 29428
rect 18929 29394 18939 29428
rect 18885 29378 18939 29394
rect 18981 29364 19035 29380
rect 18981 29336 18991 29364
rect 18671 29306 18697 29336
rect 18781 29330 18991 29336
rect 19025 29363 19035 29364
rect 19025 29333 19063 29363
rect 19147 29333 19173 29363
rect 19025 29330 19035 29333
rect 18781 29306 19035 29330
rect 18813 29254 18879 29264
rect 18813 29233 18829 29254
rect 18671 29203 18697 29233
rect 18781 29220 18829 29233
rect 18863 29220 18879 29254
rect 18781 29203 18879 29220
rect 18921 29234 19075 29264
rect 19147 29234 19173 29264
rect 18921 29161 18951 29234
rect 18897 29145 18951 29161
rect 18897 29138 18907 29145
rect 18671 29108 18697 29138
rect 18781 29111 18907 29138
rect 18941 29111 18951 29145
rect 18993 29165 19047 29181
rect 18993 29131 19003 29165
rect 19037 29135 19075 29165
rect 19147 29135 19173 29165
rect 19037 29131 19047 29135
rect 18993 29115 19047 29131
rect 18781 29108 18951 29111
rect 18897 29095 18951 29108
rect 18671 29023 18697 29053
rect 18781 29023 19063 29053
rect 19147 29023 19173 29053
rect 18861 29002 18927 29023
rect 18861 28968 18877 29002
rect 18911 28968 18927 29002
rect 18861 28958 18927 28968
rect 18677 28835 18703 28865
rect 18831 28840 19063 28865
rect 18831 28835 18930 28840
rect 18920 28806 18930 28835
rect 18964 28835 19063 28840
rect 19147 28835 19173 28865
rect 18964 28806 18974 28835
rect 18920 28790 18974 28806
rect 18677 28751 18703 28781
rect 18831 28751 18876 28781
rect 18846 28748 18876 28751
rect 19018 28751 19063 28781
rect 19147 28751 19173 28781
rect 19018 28748 19048 28751
rect 18846 28738 19048 28748
rect 18846 28718 18945 28738
rect 18929 28704 18945 28718
rect 18979 28718 19048 28738
rect 18979 28704 18995 28718
rect 18929 28694 18995 28704
rect 18663 28125 18689 28155
rect 18889 28135 19009 28155
rect 18889 28125 18937 28135
rect 18921 28101 18937 28125
rect 18971 28125 19009 28135
rect 19139 28125 19165 28155
rect 18971 28101 18987 28125
rect 18921 28091 18987 28101
rect 18663 28028 18689 28058
rect 18817 28049 18883 28058
rect 19016 28049 19055 28060
rect 18817 28030 19055 28049
rect 19139 28030 19165 28060
rect 18817 28028 19040 28030
rect 18853 28019 19040 28028
rect 18921 27874 18987 28019
rect 18921 27870 18937 27874
rect 18663 27840 18689 27870
rect 18889 27840 18937 27870
rect 18971 27872 18987 27874
rect 18971 27842 19009 27872
rect 19139 27842 19165 27872
rect 18971 27840 18987 27842
rect 18921 27830 18987 27840
rect 18921 27786 19009 27788
rect 18663 27756 18689 27786
rect 18889 27758 19009 27786
rect 19139 27758 19165 27788
rect 18889 27756 18987 27758
rect 18921 27690 18987 27756
rect 18921 27656 18937 27690
rect 18971 27656 18987 27690
rect 18921 27646 18987 27656
rect 18805 27616 18871 27626
rect 18805 27582 18821 27616
rect 18855 27598 18871 27616
rect 18855 27582 19055 27598
rect 18805 27575 19055 27582
rect 18663 27545 18689 27575
rect 18773 27568 19055 27575
rect 19139 27568 19165 27598
rect 18773 27545 18871 27568
rect 18811 27480 18865 27496
rect 18811 27461 18821 27480
rect 18663 27431 18689 27461
rect 18773 27446 18821 27461
rect 18855 27446 18865 27480
rect 18773 27431 18865 27446
rect 18811 27430 18865 27431
rect 18907 27473 19067 27503
rect 19139 27473 19165 27503
rect 18907 27388 18937 27473
rect 18871 27378 18937 27388
rect 18871 27377 18887 27378
rect 18663 27347 18689 27377
rect 18773 27347 18887 27377
rect 18871 27344 18887 27347
rect 18921 27344 18937 27378
rect 18979 27421 19045 27431
rect 18979 27387 18995 27421
rect 19029 27397 19045 27421
rect 19029 27387 19067 27397
rect 18979 27367 19067 27387
rect 19139 27367 19165 27397
rect 18871 27334 18937 27344
rect 18966 27282 19011 27296
rect 18663 27252 18689 27282
rect 18839 27266 19011 27282
rect 19139 27266 19165 27296
rect 18839 27252 18996 27266
rect 18877 27242 18931 27252
rect 18877 27208 18887 27242
rect 18921 27208 18931 27242
rect 18877 27192 18931 27208
rect 18973 27178 19027 27194
rect 18973 27150 18983 27178
rect 18663 27120 18689 27150
rect 18773 27144 18983 27150
rect 19017 27177 19027 27178
rect 19017 27147 19055 27177
rect 19139 27147 19165 27177
rect 19017 27144 19027 27147
rect 18773 27120 19027 27144
rect 18805 27068 18871 27078
rect 18805 27047 18821 27068
rect 18663 27017 18689 27047
rect 18773 27034 18821 27047
rect 18855 27034 18871 27068
rect 18773 27017 18871 27034
rect 18913 27048 19067 27078
rect 19139 27048 19165 27078
rect 18913 26975 18943 27048
rect 18889 26959 18943 26975
rect 18889 26952 18899 26959
rect 18663 26922 18689 26952
rect 18773 26925 18899 26952
rect 18933 26925 18943 26959
rect 18985 26979 19039 26995
rect 18985 26945 18995 26979
rect 19029 26949 19067 26979
rect 19139 26949 19165 26979
rect 19029 26945 19039 26949
rect 18985 26929 19039 26945
rect 18773 26922 18943 26925
rect 18889 26909 18943 26922
rect 18663 26837 18689 26867
rect 18773 26837 19055 26867
rect 19139 26837 19165 26867
rect 18853 26816 18919 26837
rect 18853 26782 18869 26816
rect 18903 26782 18919 26816
rect 18853 26772 18919 26782
rect 18669 26649 18695 26679
rect 18823 26654 19055 26679
rect 18823 26649 18922 26654
rect 18912 26620 18922 26649
rect 18956 26649 19055 26654
rect 19139 26649 19165 26679
rect 18956 26620 18966 26649
rect 18912 26604 18966 26620
rect 18669 26565 18695 26595
rect 18823 26565 18868 26595
rect 18838 26562 18868 26565
rect 19010 26565 19055 26595
rect 19139 26565 19165 26595
rect 19010 26562 19040 26565
rect 18838 26552 19040 26562
rect 18838 26532 18937 26552
rect 18921 26518 18937 26532
rect 18971 26532 19040 26552
rect 18971 26518 18987 26532
rect 18921 26508 18987 26518
rect 18667 25879 18693 25909
rect 18893 25889 19013 25909
rect 18893 25879 18941 25889
rect 18925 25855 18941 25879
rect 18975 25879 19013 25889
rect 19143 25879 19169 25909
rect 18975 25855 18991 25879
rect 18925 25845 18991 25855
rect 18667 25782 18693 25812
rect 18821 25803 18887 25812
rect 19020 25803 19059 25814
rect 18821 25784 19059 25803
rect 19143 25784 19169 25814
rect 18821 25782 19044 25784
rect 18857 25773 19044 25782
rect 18925 25628 18991 25773
rect 18925 25624 18941 25628
rect 18667 25594 18693 25624
rect 18893 25594 18941 25624
rect 18975 25626 18991 25628
rect 18975 25596 19013 25626
rect 19143 25596 19169 25626
rect 18975 25594 18991 25596
rect 18925 25584 18991 25594
rect 18925 25540 19013 25542
rect 18667 25510 18693 25540
rect 18893 25512 19013 25540
rect 19143 25512 19169 25542
rect 18893 25510 18991 25512
rect 18925 25444 18991 25510
rect 18925 25410 18941 25444
rect 18975 25410 18991 25444
rect 18925 25400 18991 25410
rect 18809 25370 18875 25380
rect 18809 25336 18825 25370
rect 18859 25352 18875 25370
rect 18859 25336 19059 25352
rect 18809 25329 19059 25336
rect 18667 25299 18693 25329
rect 18777 25322 19059 25329
rect 19143 25322 19169 25352
rect 18777 25299 18875 25322
rect 18815 25234 18869 25250
rect 18815 25215 18825 25234
rect 18667 25185 18693 25215
rect 18777 25200 18825 25215
rect 18859 25200 18869 25234
rect 18777 25185 18869 25200
rect 18815 25184 18869 25185
rect 18911 25227 19071 25257
rect 19143 25227 19169 25257
rect 18911 25142 18941 25227
rect 18875 25132 18941 25142
rect 18875 25131 18891 25132
rect 18667 25101 18693 25131
rect 18777 25101 18891 25131
rect 18875 25098 18891 25101
rect 18925 25098 18941 25132
rect 18983 25175 19049 25185
rect 18983 25141 18999 25175
rect 19033 25151 19049 25175
rect 19033 25141 19071 25151
rect 18983 25121 19071 25141
rect 19143 25121 19169 25151
rect 18875 25088 18941 25098
rect 18970 25036 19015 25050
rect 18667 25006 18693 25036
rect 18843 25020 19015 25036
rect 19143 25020 19169 25050
rect 18843 25006 19000 25020
rect 18881 24996 18935 25006
rect 18881 24962 18891 24996
rect 18925 24962 18935 24996
rect 18881 24946 18935 24962
rect 18977 24932 19031 24948
rect 18977 24904 18987 24932
rect 18667 24874 18693 24904
rect 18777 24898 18987 24904
rect 19021 24931 19031 24932
rect 19021 24901 19059 24931
rect 19143 24901 19169 24931
rect 19021 24898 19031 24901
rect 18777 24874 19031 24898
rect 18809 24822 18875 24832
rect 18809 24801 18825 24822
rect 18667 24771 18693 24801
rect 18777 24788 18825 24801
rect 18859 24788 18875 24822
rect 18777 24771 18875 24788
rect 18917 24802 19071 24832
rect 19143 24802 19169 24832
rect 18917 24729 18947 24802
rect 18893 24713 18947 24729
rect 18893 24706 18903 24713
rect 18667 24676 18693 24706
rect 18777 24679 18903 24706
rect 18937 24679 18947 24713
rect 18989 24733 19043 24749
rect 18989 24699 18999 24733
rect 19033 24703 19071 24733
rect 19143 24703 19169 24733
rect 19033 24699 19043 24703
rect 18989 24683 19043 24699
rect 18777 24676 18947 24679
rect 18893 24663 18947 24676
rect 18667 24591 18693 24621
rect 18777 24591 19059 24621
rect 19143 24591 19169 24621
rect 18857 24570 18923 24591
rect 18857 24536 18873 24570
rect 18907 24536 18923 24570
rect 18857 24526 18923 24536
rect 18673 24403 18699 24433
rect 18827 24408 19059 24433
rect 18827 24403 18926 24408
rect 18916 24374 18926 24403
rect 18960 24403 19059 24408
rect 19143 24403 19169 24433
rect 18960 24374 18970 24403
rect 18916 24358 18970 24374
rect 18673 24319 18699 24349
rect 18827 24319 18872 24349
rect 18842 24316 18872 24319
rect 19014 24319 19059 24349
rect 19143 24319 19169 24349
rect 19014 24316 19044 24319
rect 18842 24306 19044 24316
rect 18842 24286 18941 24306
rect 18925 24272 18941 24286
rect 18975 24286 19044 24306
rect 18975 24272 18991 24286
rect 18925 24262 18991 24272
rect 7749 23319 7779 23345
rect 7833 23319 7863 23345
rect 8021 23325 8051 23351
rect 8106 23325 8136 23351
rect 8201 23325 8231 23351
rect 8304 23325 8334 23351
rect 8436 23325 8466 23351
rect 8531 23325 8561 23351
rect 8615 23325 8645 23351
rect 8729 23325 8759 23351
rect 8940 23325 8970 23351
rect 9024 23325 9054 23351
rect 9212 23325 9242 23351
rect 9309 23325 9339 23351
rect 7749 23176 7779 23191
rect 7716 23146 7779 23176
rect 7716 23093 7746 23146
rect 7833 23102 7863 23191
rect 8021 23161 8051 23241
rect 7692 23077 7746 23093
rect 7692 23043 7702 23077
rect 7736 23043 7746 23077
rect 7788 23092 7863 23102
rect 7956 23145 8051 23161
rect 7956 23111 7966 23145
rect 8000 23111 8051 23145
rect 8106 23125 8136 23241
rect 8201 23209 8231 23241
rect 8201 23193 8262 23209
rect 8201 23159 8218 23193
rect 8252 23159 8262 23193
rect 8201 23143 8262 23159
rect 7956 23095 8051 23111
rect 7788 23058 7804 23092
rect 7838 23058 7863 23092
rect 7788 23048 7863 23058
rect 7692 23027 7746 23043
rect 7716 23004 7746 23027
rect 7716 22974 7779 23004
rect 7749 22959 7779 22974
rect 7833 22959 7863 23048
rect 8021 22959 8051 23095
rect 8093 23115 8159 23125
rect 8093 23081 8109 23115
rect 8143 23101 8159 23115
rect 8143 23081 8262 23101
rect 8093 23071 8262 23081
rect 8113 23019 8179 23029
rect 8113 22985 8129 23019
rect 8163 22985 8179 23019
rect 8113 22975 8179 22985
rect 8133 22947 8163 22975
rect 8232 22947 8262 23071
rect 8304 23041 8334 23241
rect 8436 23137 8466 23175
rect 8531 23143 8561 23241
rect 8615 23203 8645 23241
rect 8729 23209 8759 23241
rect 8614 23193 8680 23203
rect 8614 23159 8630 23193
rect 8664 23159 8680 23193
rect 8614 23149 8680 23159
rect 8729 23193 8810 23209
rect 8729 23159 8766 23193
rect 8800 23159 8810 23193
rect 8729 23143 8810 23159
rect 8376 23127 8466 23137
rect 8376 23093 8392 23127
rect 8426 23093 8466 23127
rect 8376 23083 8466 23093
rect 8436 23048 8466 23083
rect 8518 23127 8572 23143
rect 8518 23093 8528 23127
rect 8562 23107 8572 23127
rect 8562 23093 8687 23107
rect 8518 23077 8687 23093
rect 8304 23031 8378 23041
rect 8304 22997 8328 23031
rect 8362 22997 8378 23031
rect 8436 23018 8480 23048
rect 8450 23003 8480 23018
rect 8551 23019 8615 23035
rect 8304 22987 8378 22997
rect 8331 22959 8361 22987
rect 8551 22985 8571 23019
rect 8605 22985 8615 23019
rect 8551 22969 8615 22985
rect 8551 22947 8581 22969
rect 8657 22947 8687 23077
rect 8752 22959 8782 23143
rect 9212 23161 9242 23197
rect 9203 23131 9242 23161
rect 8940 23093 8970 23125
rect 9024 23093 9054 23125
rect 9203 23093 9233 23131
rect 9995 23323 10025 23349
rect 10079 23323 10109 23349
rect 10267 23329 10297 23355
rect 10352 23329 10382 23355
rect 10447 23329 10477 23355
rect 10550 23329 10580 23355
rect 10682 23329 10712 23355
rect 10777 23329 10807 23355
rect 10861 23329 10891 23355
rect 10975 23329 11005 23355
rect 11186 23329 11216 23355
rect 11270 23329 11300 23355
rect 11458 23329 11488 23355
rect 11555 23329 11585 23355
rect 9995 23180 10025 23195
rect 9962 23150 10025 23180
rect 9309 23093 9339 23125
rect 9962 23097 9992 23150
rect 10079 23106 10109 23195
rect 10267 23165 10297 23245
rect 8830 23077 8972 23093
rect 8830 23043 8840 23077
rect 8874 23043 8972 23077
rect 8830 23027 8972 23043
rect 9014 23077 9233 23093
rect 9014 23043 9024 23077
rect 9058 23043 9233 23077
rect 9014 23027 9233 23043
rect 9275 23077 9339 23093
rect 9275 23043 9285 23077
rect 9319 23043 9339 23077
rect 9275 23027 9339 23043
rect 9938 23081 9992 23097
rect 9938 23047 9948 23081
rect 9982 23047 9992 23081
rect 10034 23096 10109 23106
rect 10202 23149 10297 23165
rect 10202 23115 10212 23149
rect 10246 23115 10297 23149
rect 10352 23129 10382 23245
rect 10447 23213 10477 23245
rect 10447 23197 10508 23213
rect 10447 23163 10464 23197
rect 10498 23163 10508 23197
rect 10447 23147 10508 23163
rect 10202 23099 10297 23115
rect 10034 23062 10050 23096
rect 10084 23062 10109 23096
rect 10034 23052 10109 23062
rect 9938 23031 9992 23047
rect 8942 23005 8972 23027
rect 9026 23005 9056 23027
rect 9203 22998 9233 23027
rect 9309 23005 9339 23027
rect 9962 23008 9992 23031
rect 9203 22974 9244 22998
rect 9214 22959 9244 22974
rect 9962 22978 10025 23008
rect 9995 22963 10025 22978
rect 10079 22963 10109 23052
rect 10267 22963 10297 23099
rect 10339 23119 10405 23129
rect 10339 23085 10355 23119
rect 10389 23105 10405 23119
rect 10389 23085 10508 23105
rect 10339 23075 10508 23085
rect 10359 23023 10425 23033
rect 10359 22989 10375 23023
rect 10409 22989 10425 23023
rect 10359 22979 10425 22989
rect 10379 22951 10409 22979
rect 10478 22951 10508 23075
rect 10550 23045 10580 23245
rect 10682 23141 10712 23179
rect 10777 23147 10807 23245
rect 10861 23207 10891 23245
rect 10975 23213 11005 23245
rect 10860 23197 10926 23207
rect 10860 23163 10876 23197
rect 10910 23163 10926 23197
rect 10860 23153 10926 23163
rect 10975 23197 11056 23213
rect 10975 23163 11012 23197
rect 11046 23163 11056 23197
rect 10975 23147 11056 23163
rect 10622 23131 10712 23141
rect 10622 23097 10638 23131
rect 10672 23097 10712 23131
rect 10622 23087 10712 23097
rect 10682 23052 10712 23087
rect 10764 23131 10818 23147
rect 10764 23097 10774 23131
rect 10808 23111 10818 23131
rect 10808 23097 10933 23111
rect 10764 23081 10933 23097
rect 10550 23035 10624 23045
rect 10550 23001 10574 23035
rect 10608 23001 10624 23035
rect 10682 23022 10726 23052
rect 10696 23007 10726 23022
rect 10797 23023 10861 23039
rect 10550 22991 10624 23001
rect 10577 22963 10607 22991
rect 10797 22989 10817 23023
rect 10851 22989 10861 23023
rect 10797 22973 10861 22989
rect 10797 22951 10827 22973
rect 10903 22951 10933 23081
rect 10998 22963 11028 23147
rect 11458 23165 11488 23201
rect 11449 23135 11488 23165
rect 11186 23097 11216 23129
rect 11270 23097 11300 23129
rect 11449 23097 11479 23135
rect 12181 23315 12211 23341
rect 12265 23315 12295 23341
rect 12453 23321 12483 23347
rect 12538 23321 12568 23347
rect 12633 23321 12663 23347
rect 12736 23321 12766 23347
rect 12868 23321 12898 23347
rect 12963 23321 12993 23347
rect 13047 23321 13077 23347
rect 13161 23321 13191 23347
rect 13372 23321 13402 23347
rect 13456 23321 13486 23347
rect 13644 23321 13674 23347
rect 13741 23321 13771 23347
rect 12181 23172 12211 23187
rect 12148 23142 12211 23172
rect 11555 23097 11585 23129
rect 11076 23081 11218 23097
rect 11076 23047 11086 23081
rect 11120 23047 11218 23081
rect 11076 23031 11218 23047
rect 11260 23081 11479 23097
rect 11260 23047 11270 23081
rect 11304 23047 11479 23081
rect 11260 23031 11479 23047
rect 11521 23081 11585 23097
rect 12148 23089 12178 23142
rect 12265 23098 12295 23187
rect 12453 23157 12483 23237
rect 11521 23047 11531 23081
rect 11565 23047 11585 23081
rect 11521 23031 11585 23047
rect 11188 23009 11218 23031
rect 11272 23009 11302 23031
rect 11449 23002 11479 23031
rect 11555 23009 11585 23031
rect 12124 23073 12178 23089
rect 12124 23039 12134 23073
rect 12168 23039 12178 23073
rect 12220 23088 12295 23098
rect 12388 23141 12483 23157
rect 12388 23107 12398 23141
rect 12432 23107 12483 23141
rect 12538 23121 12568 23237
rect 12633 23205 12663 23237
rect 12633 23189 12694 23205
rect 12633 23155 12650 23189
rect 12684 23155 12694 23189
rect 12633 23139 12694 23155
rect 12388 23091 12483 23107
rect 12220 23054 12236 23088
rect 12270 23054 12295 23088
rect 12220 23044 12295 23054
rect 12124 23023 12178 23039
rect 11449 22978 11490 23002
rect 11460 22963 11490 22978
rect 12148 23000 12178 23023
rect 12148 22970 12211 23000
rect 12181 22955 12211 22970
rect 12265 22955 12295 23044
rect 12453 22955 12483 23091
rect 12525 23111 12591 23121
rect 12525 23077 12541 23111
rect 12575 23097 12591 23111
rect 12575 23077 12694 23097
rect 12525 23067 12694 23077
rect 12545 23015 12611 23025
rect 12545 22981 12561 23015
rect 12595 22981 12611 23015
rect 12545 22971 12611 22981
rect 7749 22849 7779 22875
rect 7833 22849 7863 22875
rect 8021 22849 8051 22875
rect 8133 22849 8163 22875
rect 8232 22849 8262 22875
rect 8331 22849 8361 22875
rect 8450 22849 8480 22875
rect 8551 22849 8581 22875
rect 8657 22849 8687 22875
rect 8752 22849 8782 22875
rect 8942 22849 8972 22875
rect 9026 22849 9056 22875
rect 9214 22849 9244 22875
rect 9309 22849 9339 22875
rect 9995 22853 10025 22879
rect 10079 22853 10109 22879
rect 10267 22853 10297 22879
rect 10379 22853 10409 22879
rect 10478 22853 10508 22879
rect 10577 22853 10607 22879
rect 10696 22853 10726 22879
rect 10797 22853 10827 22879
rect 10903 22853 10933 22879
rect 10998 22853 11028 22879
rect 11188 22853 11218 22879
rect 11272 22853 11302 22879
rect 11460 22853 11490 22879
rect 11555 22853 11585 22879
rect 12565 22943 12595 22971
rect 12664 22943 12694 23067
rect 12736 23037 12766 23237
rect 12868 23133 12898 23171
rect 12963 23139 12993 23237
rect 13047 23199 13077 23237
rect 13161 23205 13191 23237
rect 13046 23189 13112 23199
rect 13046 23155 13062 23189
rect 13096 23155 13112 23189
rect 13046 23145 13112 23155
rect 13161 23189 13242 23205
rect 13161 23155 13198 23189
rect 13232 23155 13242 23189
rect 13161 23139 13242 23155
rect 12808 23123 12898 23133
rect 12808 23089 12824 23123
rect 12858 23089 12898 23123
rect 12808 23079 12898 23089
rect 12868 23044 12898 23079
rect 12950 23123 13004 23139
rect 12950 23089 12960 23123
rect 12994 23103 13004 23123
rect 12994 23089 13119 23103
rect 12950 23073 13119 23089
rect 12736 23027 12810 23037
rect 12736 22993 12760 23027
rect 12794 22993 12810 23027
rect 12868 23014 12912 23044
rect 12882 22999 12912 23014
rect 12983 23015 13047 23031
rect 12736 22983 12810 22993
rect 12763 22955 12793 22983
rect 12983 22981 13003 23015
rect 13037 22981 13047 23015
rect 12983 22965 13047 22981
rect 12983 22943 13013 22965
rect 13089 22943 13119 23073
rect 13184 22955 13214 23139
rect 13644 23157 13674 23193
rect 13635 23127 13674 23157
rect 13372 23089 13402 23121
rect 13456 23089 13486 23121
rect 13635 23089 13665 23127
rect 14427 23319 14457 23345
rect 14511 23319 14541 23345
rect 14699 23325 14729 23351
rect 14784 23325 14814 23351
rect 14879 23325 14909 23351
rect 14982 23325 15012 23351
rect 15114 23325 15144 23351
rect 15209 23325 15239 23351
rect 15293 23325 15323 23351
rect 15407 23325 15437 23351
rect 15618 23325 15648 23351
rect 15702 23325 15732 23351
rect 15890 23325 15920 23351
rect 15987 23325 16017 23351
rect 14427 23176 14457 23191
rect 14394 23146 14457 23176
rect 13741 23089 13771 23121
rect 14394 23093 14424 23146
rect 14511 23102 14541 23191
rect 14699 23161 14729 23241
rect 13262 23073 13404 23089
rect 13262 23039 13272 23073
rect 13306 23039 13404 23073
rect 13262 23023 13404 23039
rect 13446 23073 13665 23089
rect 13446 23039 13456 23073
rect 13490 23039 13665 23073
rect 13446 23023 13665 23039
rect 13707 23073 13771 23089
rect 13707 23039 13717 23073
rect 13751 23039 13771 23073
rect 13707 23023 13771 23039
rect 14370 23077 14424 23093
rect 14370 23043 14380 23077
rect 14414 23043 14424 23077
rect 14466 23092 14541 23102
rect 14634 23145 14729 23161
rect 14634 23111 14644 23145
rect 14678 23111 14729 23145
rect 14784 23125 14814 23241
rect 14879 23209 14909 23241
rect 14879 23193 14940 23209
rect 14879 23159 14896 23193
rect 14930 23159 14940 23193
rect 14879 23143 14940 23159
rect 14634 23095 14729 23111
rect 14466 23058 14482 23092
rect 14516 23058 14541 23092
rect 14466 23048 14541 23058
rect 14370 23027 14424 23043
rect 13374 23001 13404 23023
rect 13458 23001 13488 23023
rect 13635 22994 13665 23023
rect 13741 23001 13771 23023
rect 14394 23004 14424 23027
rect 13635 22970 13676 22994
rect 13646 22955 13676 22970
rect 14394 22974 14457 23004
rect 14427 22959 14457 22974
rect 14511 22959 14541 23048
rect 14699 22959 14729 23095
rect 14771 23115 14837 23125
rect 14771 23081 14787 23115
rect 14821 23101 14837 23115
rect 14821 23081 14940 23101
rect 14771 23071 14940 23081
rect 14791 23019 14857 23029
rect 14791 22985 14807 23019
rect 14841 22985 14857 23019
rect 14791 22975 14857 22985
rect 14811 22947 14841 22975
rect 14910 22947 14940 23071
rect 14982 23041 15012 23241
rect 15114 23137 15144 23175
rect 15209 23143 15239 23241
rect 15293 23203 15323 23241
rect 15407 23209 15437 23241
rect 15292 23193 15358 23203
rect 15292 23159 15308 23193
rect 15342 23159 15358 23193
rect 15292 23149 15358 23159
rect 15407 23193 15488 23209
rect 15407 23159 15444 23193
rect 15478 23159 15488 23193
rect 15407 23143 15488 23159
rect 15054 23127 15144 23137
rect 15054 23093 15070 23127
rect 15104 23093 15144 23127
rect 15054 23083 15144 23093
rect 15114 23048 15144 23083
rect 15196 23127 15250 23143
rect 15196 23093 15206 23127
rect 15240 23107 15250 23127
rect 15240 23093 15365 23107
rect 15196 23077 15365 23093
rect 14982 23031 15056 23041
rect 14982 22997 15006 23031
rect 15040 22997 15056 23031
rect 15114 23018 15158 23048
rect 15128 23003 15158 23018
rect 15229 23019 15293 23035
rect 14982 22987 15056 22997
rect 15009 22959 15039 22987
rect 15229 22985 15249 23019
rect 15283 22985 15293 23019
rect 15229 22969 15293 22985
rect 15229 22947 15259 22969
rect 15335 22947 15365 23077
rect 15430 22959 15460 23143
rect 15890 23161 15920 23197
rect 15881 23131 15920 23161
rect 15618 23093 15648 23125
rect 15702 23093 15732 23125
rect 15881 23093 15911 23131
rect 16709 23319 16739 23345
rect 16793 23319 16823 23345
rect 16981 23325 17011 23351
rect 17066 23325 17096 23351
rect 17161 23325 17191 23351
rect 17264 23325 17294 23351
rect 17396 23325 17426 23351
rect 17491 23325 17521 23351
rect 17575 23325 17605 23351
rect 17689 23325 17719 23351
rect 17900 23325 17930 23351
rect 17984 23325 18014 23351
rect 18172 23325 18202 23351
rect 18269 23325 18299 23351
rect 16709 23176 16739 23191
rect 16676 23146 16739 23176
rect 15987 23093 16017 23125
rect 16676 23093 16706 23146
rect 16793 23102 16823 23191
rect 16981 23161 17011 23241
rect 15508 23077 15650 23093
rect 15508 23043 15518 23077
rect 15552 23043 15650 23077
rect 15508 23027 15650 23043
rect 15692 23077 15911 23093
rect 15692 23043 15702 23077
rect 15736 23043 15911 23077
rect 15692 23027 15911 23043
rect 15953 23077 16017 23093
rect 15953 23043 15963 23077
rect 15997 23043 16017 23077
rect 15953 23027 16017 23043
rect 16652 23077 16706 23093
rect 16652 23043 16662 23077
rect 16696 23043 16706 23077
rect 16748 23092 16823 23102
rect 16916 23145 17011 23161
rect 16916 23111 16926 23145
rect 16960 23111 17011 23145
rect 17066 23125 17096 23241
rect 17161 23209 17191 23241
rect 17161 23193 17222 23209
rect 17161 23159 17178 23193
rect 17212 23159 17222 23193
rect 17161 23143 17222 23159
rect 16916 23095 17011 23111
rect 16748 23058 16764 23092
rect 16798 23058 16823 23092
rect 16748 23048 16823 23058
rect 16652 23027 16706 23043
rect 15620 23005 15650 23027
rect 15704 23005 15734 23027
rect 15881 22998 15911 23027
rect 15987 23005 16017 23027
rect 15881 22974 15922 22998
rect 15892 22959 15922 22974
rect 16676 23004 16706 23027
rect 16676 22974 16739 23004
rect 16709 22959 16739 22974
rect 16793 22959 16823 23048
rect 16981 22959 17011 23095
rect 17053 23115 17119 23125
rect 17053 23081 17069 23115
rect 17103 23101 17119 23115
rect 17103 23081 17222 23101
rect 17053 23071 17222 23081
rect 17073 23019 17139 23029
rect 17073 22985 17089 23019
rect 17123 22985 17139 23019
rect 17073 22975 17139 22985
rect 17093 22947 17123 22975
rect 17192 22947 17222 23071
rect 17264 23041 17294 23241
rect 17396 23137 17426 23175
rect 17491 23143 17521 23241
rect 17575 23203 17605 23241
rect 17689 23209 17719 23241
rect 17574 23193 17640 23203
rect 17574 23159 17590 23193
rect 17624 23159 17640 23193
rect 17574 23149 17640 23159
rect 17689 23193 17770 23209
rect 17689 23159 17726 23193
rect 17760 23159 17770 23193
rect 17689 23143 17770 23159
rect 17336 23127 17426 23137
rect 17336 23093 17352 23127
rect 17386 23093 17426 23127
rect 17336 23083 17426 23093
rect 17396 23048 17426 23083
rect 17478 23127 17532 23143
rect 17478 23093 17488 23127
rect 17522 23107 17532 23127
rect 17522 23093 17647 23107
rect 17478 23077 17647 23093
rect 17264 23031 17338 23041
rect 17264 22997 17288 23031
rect 17322 22997 17338 23031
rect 17396 23018 17440 23048
rect 17410 23003 17440 23018
rect 17511 23019 17575 23035
rect 17264 22987 17338 22997
rect 17291 22959 17321 22987
rect 17511 22985 17531 23019
rect 17565 22985 17575 23019
rect 17511 22969 17575 22985
rect 17511 22947 17541 22969
rect 17617 22947 17647 23077
rect 17712 22959 17742 23143
rect 18172 23161 18202 23197
rect 18163 23131 18202 23161
rect 17900 23093 17930 23125
rect 17984 23093 18014 23125
rect 18163 23093 18193 23131
rect 18269 23093 18299 23125
rect 17790 23077 17932 23093
rect 17790 23043 17800 23077
rect 17834 23043 17932 23077
rect 17790 23027 17932 23043
rect 17974 23077 18193 23093
rect 17974 23043 17984 23077
rect 18018 23043 18193 23077
rect 17974 23027 18193 23043
rect 18235 23077 18299 23093
rect 18235 23043 18245 23077
rect 18279 23043 18299 23077
rect 18235 23027 18299 23043
rect 17902 23005 17932 23027
rect 17986 23005 18016 23027
rect 18163 22998 18193 23027
rect 18269 23005 18299 23027
rect 18163 22974 18204 22998
rect 18174 22959 18204 22974
rect 12181 22845 12211 22871
rect 12265 22845 12295 22871
rect 12453 22845 12483 22871
rect 12565 22845 12595 22871
rect 12664 22845 12694 22871
rect 12763 22845 12793 22871
rect 12882 22845 12912 22871
rect 12983 22845 13013 22871
rect 13089 22845 13119 22871
rect 13184 22845 13214 22871
rect 13374 22845 13404 22871
rect 13458 22845 13488 22871
rect 13646 22845 13676 22871
rect 13741 22845 13771 22871
rect 14427 22849 14457 22875
rect 14511 22849 14541 22875
rect 14699 22849 14729 22875
rect 14811 22849 14841 22875
rect 14910 22849 14940 22875
rect 15009 22849 15039 22875
rect 15128 22849 15158 22875
rect 15229 22849 15259 22875
rect 15335 22849 15365 22875
rect 15430 22849 15460 22875
rect 15620 22849 15650 22875
rect 15704 22849 15734 22875
rect 15892 22849 15922 22875
rect 15987 22849 16017 22875
rect 16709 22849 16739 22875
rect 16793 22849 16823 22875
rect 16981 22849 17011 22875
rect 17093 22849 17123 22875
rect 17192 22849 17222 22875
rect 17291 22849 17321 22875
rect 17410 22849 17440 22875
rect 17511 22849 17541 22875
rect 17617 22849 17647 22875
rect 17712 22849 17742 22875
rect 17902 22849 17932 22875
rect 17986 22849 18016 22875
rect 18174 22849 18204 22875
rect 18269 22849 18299 22875
rect 9556 17747 9586 17773
rect 16471 17637 16501 17663
rect 17345 17639 17375 17665
rect 9556 17595 9586 17617
rect 15693 17599 15723 17625
rect 9556 17579 9642 17595
rect 9556 17545 9592 17579
rect 9626 17545 9642 17579
rect 9556 17529 9642 17545
rect 9556 17497 9586 17529
rect 18113 17629 18143 17655
rect 19235 17631 19265 17657
rect 20109 17633 20139 17659
rect 16471 17485 16501 17507
rect 17345 17487 17375 17509
rect 20877 17623 20907 17649
rect 16471 17469 16557 17485
rect 15693 17447 15723 17469
rect 15693 17431 15779 17447
rect 15693 17397 15729 17431
rect 15763 17397 15779 17431
rect 15693 17381 15779 17397
rect 16471 17435 16507 17469
rect 16541 17435 16557 17469
rect 16471 17419 16557 17435
rect 17345 17471 17431 17487
rect 17345 17437 17381 17471
rect 17415 17437 17431 17471
rect 17345 17421 17431 17437
rect 18113 17477 18143 17499
rect 19235 17479 19265 17501
rect 20109 17481 20139 17503
rect 21491 17621 21521 17647
rect 22365 17623 22395 17649
rect 18113 17461 18199 17477
rect 18113 17427 18149 17461
rect 18183 17427 18199 17461
rect 16471 17387 16501 17419
rect 17345 17389 17375 17421
rect 18113 17411 18199 17427
rect 19235 17463 19321 17479
rect 19235 17429 19271 17463
rect 19305 17429 19321 17463
rect 19235 17413 19321 17429
rect 20109 17465 20195 17481
rect 20109 17431 20145 17465
rect 20179 17431 20195 17465
rect 20109 17415 20195 17431
rect 20877 17471 20907 17493
rect 23133 17613 23163 17639
rect 20877 17455 20963 17471
rect 20877 17421 20913 17455
rect 20947 17421 20963 17455
rect 15693 17349 15723 17381
rect 9556 17271 9586 17297
rect 18113 17379 18143 17411
rect 19235 17381 19265 17413
rect 20109 17383 20139 17415
rect 20877 17405 20963 17421
rect 21491 17469 21521 17491
rect 22365 17471 22395 17493
rect 21491 17453 21577 17469
rect 21491 17419 21527 17453
rect 21561 17419 21577 17453
rect 16471 17161 16501 17187
rect 17345 17163 17375 17189
rect 20877 17373 20907 17405
rect 21491 17403 21577 17419
rect 22365 17455 22451 17471
rect 22365 17421 22401 17455
rect 22435 17421 22451 17455
rect 22365 17405 22451 17421
rect 23133 17461 23163 17483
rect 23133 17445 23219 17461
rect 23133 17411 23169 17445
rect 23203 17411 23219 17445
rect 18113 17153 18143 17179
rect 19235 17155 19265 17181
rect 20109 17157 20139 17183
rect 21491 17371 21521 17403
rect 22365 17373 22395 17405
rect 23133 17395 23219 17411
rect 15693 17123 15723 17149
rect 20877 17147 20907 17173
rect 23133 17363 23163 17395
rect 21491 17145 21521 17171
rect 22365 17147 22395 17173
rect 23133 17137 23163 17163
rect 16456 16647 16486 16673
rect 4555 16539 4585 16565
rect 4639 16539 4669 16565
rect 4723 16539 4753 16565
rect 4807 16539 4837 16565
rect 4995 16539 5025 16565
rect 9421 16543 9451 16569
rect 9505 16543 9535 16569
rect 9589 16543 9619 16569
rect 9673 16543 9703 16569
rect 9861 16543 9891 16569
rect 17224 16637 17254 16663
rect 18098 16639 18128 16665
rect 16456 16415 16486 16447
rect 18712 16637 18742 16663
rect 16400 16399 16486 16415
rect 17224 16405 17254 16437
rect 18098 16407 18128 16439
rect 19480 16627 19510 16653
rect 20354 16629 20384 16655
rect 21476 16631 21506 16657
rect 16400 16365 16416 16399
rect 16450 16365 16486 16399
rect 16400 16349 16486 16365
rect 4555 16307 4585 16339
rect 4639 16307 4669 16339
rect 4723 16307 4753 16339
rect 4807 16307 4837 16339
rect 4995 16307 5025 16339
rect 9421 16311 9451 16343
rect 9505 16311 9535 16343
rect 9589 16311 9619 16343
rect 9673 16311 9703 16343
rect 9861 16311 9891 16343
rect 16456 16327 16486 16349
rect 17168 16389 17254 16405
rect 17168 16355 17184 16389
rect 17218 16355 17254 16389
rect 17168 16339 17254 16355
rect 18042 16391 18128 16407
rect 18712 16405 18742 16437
rect 22244 16621 22274 16647
rect 23118 16623 23148 16649
rect 18042 16357 18058 16391
rect 18092 16357 18128 16391
rect 18042 16341 18128 16357
rect 4543 16291 4597 16307
rect 4543 16257 4553 16291
rect 4587 16257 4597 16291
rect 4543 16241 4597 16257
rect 4639 16291 4753 16307
rect 4639 16257 4670 16291
rect 4704 16257 4753 16291
rect 4639 16241 4753 16257
rect 4795 16291 4849 16307
rect 4795 16257 4805 16291
rect 4839 16257 4849 16291
rect 4795 16241 4849 16257
rect 4891 16291 5025 16307
rect 4891 16257 4901 16291
rect 4935 16274 5025 16291
rect 9409 16295 9463 16311
rect 4935 16257 5021 16274
rect 4891 16241 5021 16257
rect 9409 16261 9419 16295
rect 9453 16261 9463 16295
rect 9409 16245 9463 16261
rect 9505 16295 9619 16311
rect 9505 16261 9536 16295
rect 9570 16261 9619 16295
rect 9505 16245 9619 16261
rect 9661 16295 9715 16311
rect 9661 16261 9671 16295
rect 9705 16261 9715 16295
rect 9661 16245 9715 16261
rect 9757 16295 9891 16311
rect 9757 16261 9767 16295
rect 9801 16278 9891 16295
rect 9801 16261 9887 16278
rect 9757 16245 9887 16261
rect 4555 16219 4585 16241
rect 4639 16219 4669 16241
rect 4723 16219 4753 16241
rect 4807 16219 4837 16241
rect 4991 16219 5021 16241
rect 9421 16223 9451 16245
rect 9505 16223 9535 16245
rect 9589 16223 9619 16245
rect 9673 16223 9703 16245
rect 9857 16223 9887 16245
rect 17224 16317 17254 16339
rect 18098 16319 18128 16341
rect 18656 16389 18742 16405
rect 19480 16395 19510 16427
rect 20354 16397 20384 16429
rect 21476 16399 21506 16431
rect 18656 16355 18672 16389
rect 18706 16355 18742 16389
rect 18656 16339 18742 16355
rect 16456 16171 16486 16197
rect 18712 16317 18742 16339
rect 19424 16379 19510 16395
rect 19424 16345 19440 16379
rect 19474 16345 19510 16379
rect 19424 16329 19510 16345
rect 20298 16381 20384 16397
rect 20298 16347 20314 16381
rect 20348 16347 20384 16381
rect 20298 16331 20384 16347
rect 21420 16383 21506 16399
rect 22244 16389 22274 16421
rect 23118 16391 23148 16423
rect 21420 16349 21436 16383
rect 21470 16349 21506 16383
rect 21420 16333 21506 16349
rect 17224 16161 17254 16187
rect 18098 16163 18128 16189
rect 19480 16307 19510 16329
rect 20354 16309 20384 16331
rect 21476 16311 21506 16333
rect 22188 16373 22274 16389
rect 22188 16339 22204 16373
rect 22238 16339 22274 16373
rect 22188 16323 22274 16339
rect 23062 16375 23148 16391
rect 23062 16341 23078 16375
rect 23112 16341 23148 16375
rect 23062 16325 23148 16341
rect 18712 16161 18742 16187
rect 22244 16301 22274 16323
rect 23118 16303 23148 16325
rect 19480 16151 19510 16177
rect 20354 16153 20384 16179
rect 21476 16155 21506 16181
rect 22244 16145 22274 16171
rect 23118 16147 23148 16173
rect 4555 16063 4585 16089
rect 4639 16063 4669 16089
rect 4723 16063 4753 16089
rect 4807 16063 4837 16089
rect 4991 16063 5021 16089
rect 9421 16067 9451 16093
rect 9505 16067 9535 16093
rect 9589 16067 9619 16093
rect 9673 16067 9703 16093
rect 9857 16067 9887 16093
rect 4873 15795 4903 15821
rect 9739 15799 9769 15825
rect 4681 15753 4711 15779
rect 4765 15753 4795 15779
rect 4681 15563 4711 15669
rect 4624 15547 4711 15563
rect 4624 15513 4640 15547
rect 4674 15513 4711 15547
rect 4624 15497 4711 15513
rect 4681 15457 4711 15497
rect 4765 15563 4795 15669
rect 9547 15757 9577 15783
rect 9631 15757 9661 15783
rect 6687 15685 6717 15711
rect 6787 15685 6817 15711
rect 6891 15685 6921 15711
rect 6977 15685 7007 15711
rect 7143 15685 7173 15711
rect 4873 15563 4903 15595
rect 4765 15547 4831 15563
rect 4765 15513 4781 15547
rect 4815 15513 4831 15547
rect 4765 15497 4831 15513
rect 4873 15547 4939 15563
rect 4873 15513 4889 15547
rect 4923 15513 4939 15547
rect 4873 15497 4939 15513
rect 4765 15457 4795 15497
rect 4873 15475 4903 15497
rect 4681 15347 4711 15373
rect 4765 15347 4795 15373
rect 6687 15453 6717 15601
rect 6787 15453 6817 15601
rect 6891 15453 6921 15601
rect 6977 15453 7007 15601
rect 9547 15567 9577 15673
rect 9490 15551 9577 15567
rect 9490 15517 9506 15551
rect 9540 15517 9577 15551
rect 9490 15501 9577 15517
rect 7143 15453 7173 15485
rect 6629 15437 6717 15453
rect 6629 15403 6639 15437
rect 6673 15403 6717 15437
rect 6629 15387 6717 15403
rect 4873 15319 4903 15345
rect 6687 15319 6717 15387
rect 6775 15437 6829 15453
rect 6775 15403 6785 15437
rect 6819 15403 6829 15437
rect 6775 15387 6829 15403
rect 6881 15437 6935 15453
rect 6881 15403 6891 15437
rect 6925 15403 6935 15437
rect 6881 15387 6935 15403
rect 6977 15437 7041 15453
rect 6977 15403 6987 15437
rect 7021 15403 7041 15437
rect 6977 15387 7041 15403
rect 7088 15437 7173 15453
rect 7088 15403 7098 15437
rect 7132 15403 7173 15437
rect 7088 15387 7173 15403
rect 6775 15319 6805 15387
rect 6881 15319 6911 15387
rect 6977 15319 7007 15387
rect 7143 15365 7173 15387
rect 9547 15461 9577 15501
rect 9631 15567 9661 15673
rect 11553 15689 11583 15715
rect 11653 15689 11683 15715
rect 11757 15689 11787 15715
rect 11843 15689 11873 15715
rect 12009 15689 12039 15715
rect 9739 15567 9769 15599
rect 9631 15551 9697 15567
rect 9631 15517 9647 15551
rect 9681 15517 9697 15551
rect 9631 15501 9697 15517
rect 9739 15551 9805 15567
rect 9739 15517 9755 15551
rect 9789 15517 9805 15551
rect 9739 15501 9805 15517
rect 9631 15461 9661 15501
rect 9739 15479 9769 15501
rect 9547 15351 9577 15377
rect 9631 15351 9661 15377
rect 11553 15457 11583 15605
rect 11653 15457 11683 15605
rect 11757 15457 11787 15605
rect 11843 15457 11873 15605
rect 12009 15457 12039 15489
rect 11495 15441 11583 15457
rect 11495 15407 11505 15441
rect 11539 15407 11583 15441
rect 11495 15391 11583 15407
rect 9739 15323 9769 15349
rect 11553 15323 11583 15391
rect 11641 15441 11695 15457
rect 11641 15407 11651 15441
rect 11685 15407 11695 15441
rect 11641 15391 11695 15407
rect 11747 15441 11801 15457
rect 11747 15407 11757 15441
rect 11791 15407 11801 15441
rect 11747 15391 11801 15407
rect 11843 15441 11907 15457
rect 11843 15407 11853 15441
rect 11887 15407 11907 15441
rect 11843 15391 11907 15407
rect 11954 15441 12039 15457
rect 11954 15407 11964 15441
rect 11998 15407 12039 15441
rect 11954 15391 12039 15407
rect 11641 15323 11671 15391
rect 11747 15323 11777 15391
rect 11843 15323 11873 15391
rect 12009 15369 12039 15391
rect 6057 15185 6087 15211
rect 6687 15209 6717 15235
rect 6775 15209 6805 15235
rect 6881 15209 6911 15235
rect 6977 15209 7007 15235
rect 7143 15209 7173 15235
rect 10923 15189 10953 15215
rect 11553 15213 11583 15239
rect 11641 15213 11671 15239
rect 11747 15213 11777 15239
rect 11843 15213 11873 15239
rect 12009 15213 12039 15239
rect 5865 15143 5895 15169
rect 5949 15143 5979 15169
rect 4565 14975 4595 15001
rect 4649 14975 4679 15001
rect 4733 14975 4763 15001
rect 4817 14975 4847 15001
rect 5005 14975 5035 15001
rect 5865 14953 5895 15059
rect 5808 14937 5895 14953
rect 5808 14903 5824 14937
rect 5858 14903 5895 14937
rect 5808 14887 5895 14903
rect 5865 14847 5895 14887
rect 5949 14953 5979 15059
rect 10731 15147 10761 15173
rect 10815 15147 10845 15173
rect 6057 14953 6087 14985
rect 9431 14979 9461 15005
rect 9515 14979 9545 15005
rect 9599 14979 9629 15005
rect 9683 14979 9713 15005
rect 9871 14979 9901 15005
rect 5949 14937 6015 14953
rect 5949 14903 5965 14937
rect 5999 14903 6015 14937
rect 5949 14887 6015 14903
rect 6057 14937 6123 14953
rect 6057 14903 6073 14937
rect 6107 14903 6123 14937
rect 6057 14887 6123 14903
rect 5949 14847 5979 14887
rect 6057 14865 6087 14887
rect 4565 14743 4595 14775
rect 4649 14743 4679 14775
rect 4733 14743 4763 14775
rect 4817 14743 4847 14775
rect 5005 14743 5035 14775
rect 4553 14727 4607 14743
rect 4553 14693 4563 14727
rect 4597 14693 4607 14727
rect 4553 14677 4607 14693
rect 4649 14727 4763 14743
rect 4649 14693 4680 14727
rect 4714 14693 4763 14727
rect 4649 14677 4763 14693
rect 4805 14727 4859 14743
rect 4805 14693 4815 14727
rect 4849 14693 4859 14727
rect 4805 14677 4859 14693
rect 4901 14727 5035 14743
rect 5865 14737 5895 14763
rect 5949 14737 5979 14763
rect 10731 14957 10761 15063
rect 10674 14941 10761 14957
rect 10674 14907 10690 14941
rect 10724 14907 10761 14941
rect 10674 14891 10761 14907
rect 10731 14851 10761 14891
rect 10815 14957 10845 15063
rect 10923 14957 10953 14989
rect 10815 14941 10881 14957
rect 10815 14907 10831 14941
rect 10865 14907 10881 14941
rect 10815 14891 10881 14907
rect 10923 14941 10989 14957
rect 10923 14907 10939 14941
rect 10973 14907 10989 14941
rect 10923 14891 10989 14907
rect 10815 14851 10845 14891
rect 10923 14869 10953 14891
rect 9431 14747 9461 14779
rect 9515 14747 9545 14779
rect 9599 14747 9629 14779
rect 9683 14747 9713 14779
rect 9871 14747 9901 14779
rect 4901 14693 4911 14727
rect 4945 14710 5035 14727
rect 4945 14693 5031 14710
rect 6057 14709 6087 14735
rect 9419 14731 9473 14747
rect 4901 14677 5031 14693
rect 9419 14697 9429 14731
rect 9463 14697 9473 14731
rect 9419 14681 9473 14697
rect 9515 14731 9629 14747
rect 9515 14697 9546 14731
rect 9580 14697 9629 14731
rect 9515 14681 9629 14697
rect 9671 14731 9725 14747
rect 9671 14697 9681 14731
rect 9715 14697 9725 14731
rect 9671 14681 9725 14697
rect 9767 14731 9901 14747
rect 10731 14741 10761 14767
rect 10815 14741 10845 14767
rect 23563 14785 23593 14811
rect 23647 14785 23677 14811
rect 9767 14697 9777 14731
rect 9811 14714 9901 14731
rect 9811 14697 9897 14714
rect 10923 14713 10953 14739
rect 23835 14735 23865 14811
rect 23919 14735 23949 14811
rect 24107 14785 24137 14811
rect 9767 14681 9897 14697
rect 4565 14655 4595 14677
rect 4649 14655 4679 14677
rect 4733 14655 4763 14677
rect 4817 14655 4847 14677
rect 5001 14655 5031 14677
rect 9431 14659 9461 14681
rect 9515 14659 9545 14681
rect 9599 14659 9629 14681
rect 9683 14659 9713 14681
rect 9867 14659 9897 14681
rect 23563 14553 23593 14701
rect 23647 14553 23677 14701
rect 24293 14735 24323 14811
rect 24377 14735 24407 14810
rect 24472 14785 24502 14811
rect 24556 14785 24586 14811
rect 24744 14785 24774 14811
rect 24932 14785 24962 14811
rect 23835 14555 23865 14651
rect 23919 14636 23949 14651
rect 24107 14636 24137 14701
rect 25029 14738 25059 14811
rect 25307 14785 25337 14811
rect 24293 14636 24323 14651
rect 23919 14606 24323 14636
rect 24016 14561 24129 14606
rect 23539 14537 23593 14553
rect 4565 14499 4595 14525
rect 4649 14499 4679 14525
rect 4733 14499 4763 14525
rect 4817 14499 4847 14525
rect 5001 14499 5031 14525
rect 9431 14503 9461 14529
rect 9515 14503 9545 14529
rect 9599 14503 9629 14529
rect 9683 14503 9713 14529
rect 9867 14503 9897 14529
rect 23539 14503 23549 14537
rect 23583 14503 23593 14537
rect 23539 14487 23593 14503
rect 23635 14537 23689 14553
rect 23635 14503 23645 14537
rect 23679 14503 23689 14537
rect 23635 14487 23689 14503
rect 23731 14545 23966 14555
rect 23731 14525 23916 14545
rect 23563 14419 23593 14487
rect 23647 14419 23677 14487
rect 23731 14419 23761 14525
rect 23900 14511 23916 14525
rect 23950 14511 23966 14545
rect 23900 14501 23966 14511
rect 24016 14541 24234 14561
rect 24377 14553 24407 14651
rect 24472 14565 24502 14701
rect 24556 14565 24586 14701
rect 24016 14507 24150 14541
rect 24184 14507 24234 14541
rect 24016 14487 24234 14507
rect 23828 14453 23858 14479
rect 24016 14462 24046 14487
rect 24204 14469 24234 14487
rect 24288 14541 24407 14553
rect 24288 14507 24315 14541
rect 24349 14523 24407 14541
rect 24449 14549 24514 14565
rect 24349 14507 24365 14523
rect 24288 14497 24365 14507
rect 24449 14515 24459 14549
rect 24493 14515 24514 14549
rect 24449 14499 24514 14515
rect 24556 14549 24610 14565
rect 24744 14553 24774 14701
rect 24932 14553 24962 14701
rect 25029 14553 25059 14654
rect 25307 14553 25337 14585
rect 24556 14515 24566 14549
rect 24600 14515 24610 14549
rect 24556 14499 24610 14515
rect 24685 14537 24964 14553
rect 24685 14503 24695 14537
rect 24729 14503 24964 14537
rect 25029 14543 25188 14553
rect 25029 14523 25138 14543
rect 24288 14469 24318 14497
rect 24474 14419 24504 14499
rect 24558 14419 24588 14499
rect 24685 14488 24964 14503
rect 24685 14487 24776 14488
rect 24746 14419 24776 14487
rect 24934 14419 24964 14488
rect 25087 14509 25138 14523
rect 25172 14509 25188 14543
rect 25087 14499 25188 14509
rect 25263 14537 25337 14553
rect 25263 14503 25275 14537
rect 25309 14503 25337 14537
rect 25087 14469 25117 14499
rect 25263 14487 25337 14503
rect 23828 14339 23858 14369
rect 24016 14339 24046 14378
rect 23563 14309 23593 14335
rect 23647 14309 23677 14335
rect 23731 14309 23761 14335
rect 23828 14309 24046 14339
rect 24204 14309 24234 14385
rect 24288 14309 24318 14385
rect 25307 14465 25337 14487
rect 24474 14309 24504 14335
rect 24558 14309 24588 14335
rect 24746 14309 24776 14335
rect 24934 14309 24964 14335
rect 25087 14309 25117 14385
rect 25307 14309 25337 14335
rect 4883 14231 4913 14257
rect 4691 14189 4721 14215
rect 4775 14189 4805 14215
rect 4691 13999 4721 14105
rect 4634 13983 4721 13999
rect 4634 13949 4650 13983
rect 4684 13949 4721 13983
rect 4634 13933 4721 13949
rect 4691 13893 4721 13933
rect 4775 13999 4805 14105
rect 5903 14219 5933 14245
rect 6003 14219 6033 14245
rect 6107 14219 6137 14245
rect 6193 14219 6223 14245
rect 6359 14219 6389 14245
rect 9749 14235 9779 14261
rect 4883 13999 4913 14031
rect 4775 13983 4841 13999
rect 4775 13949 4791 13983
rect 4825 13949 4841 13983
rect 4775 13933 4841 13949
rect 4883 13983 4949 13999
rect 5903 13987 5933 14135
rect 6003 13987 6033 14135
rect 6107 13987 6137 14135
rect 6193 13987 6223 14135
rect 8163 14203 8193 14229
rect 7963 14179 8029 14189
rect 7963 14145 7979 14179
rect 8013 14145 8029 14179
rect 7963 14135 8029 14145
rect 7801 14087 7831 14113
rect 7897 14087 7927 14113
rect 7969 14087 7999 14135
rect 8065 14087 8095 14113
rect 6359 13987 6389 14019
rect 9557 14193 9587 14219
rect 9641 14193 9671 14219
rect 9557 14003 9587 14109
rect 4883 13949 4899 13983
rect 4933 13949 4949 13983
rect 4883 13933 4949 13949
rect 5845 13971 5933 13987
rect 5845 13937 5855 13971
rect 5889 13937 5933 13971
rect 4775 13893 4805 13933
rect 4883 13911 4913 13933
rect 5845 13921 5933 13937
rect 4691 13783 4721 13809
rect 4775 13783 4805 13809
rect 5903 13853 5933 13921
rect 5991 13971 6045 13987
rect 5991 13937 6001 13971
rect 6035 13937 6045 13971
rect 5991 13921 6045 13937
rect 6097 13971 6151 13987
rect 6097 13937 6107 13971
rect 6141 13937 6151 13971
rect 6097 13921 6151 13937
rect 6193 13971 6257 13987
rect 6193 13937 6203 13971
rect 6237 13937 6257 13971
rect 6193 13921 6257 13937
rect 6304 13971 6389 13987
rect 7801 13971 7831 14003
rect 7897 13971 7927 14003
rect 6304 13937 6314 13971
rect 6348 13937 6389 13971
rect 6304 13921 6389 13937
rect 5991 13853 6021 13921
rect 6097 13853 6127 13921
rect 6193 13853 6223 13921
rect 6359 13899 6389 13921
rect 7747 13955 7831 13971
rect 7747 13921 7757 13955
rect 7791 13921 7831 13955
rect 7747 13905 7831 13921
rect 7873 13955 7927 13971
rect 7873 13921 7883 13955
rect 7917 13921 7927 13955
rect 7873 13905 7927 13921
rect 4883 13755 4913 13781
rect 7083 13845 7113 13871
rect 5903 13743 5933 13769
rect 5991 13743 6021 13769
rect 6097 13743 6127 13769
rect 6193 13743 6223 13769
rect 6359 13743 6389 13769
rect 6914 13729 6944 13755
rect 6986 13729 7016 13755
rect 7801 13843 7831 13905
rect 7897 13843 7927 13905
rect 7969 13888 7999 14003
rect 8065 13971 8095 14003
rect 8163 13971 8193 14003
rect 9500 13987 9587 14003
rect 8049 13955 8103 13971
rect 8049 13921 8059 13955
rect 8093 13921 8103 13955
rect 8049 13905 8103 13921
rect 8145 13955 8200 13971
rect 8145 13921 8155 13955
rect 8189 13921 8200 13955
rect 9500 13953 9516 13987
rect 9550 13953 9587 13987
rect 9500 13937 9587 13953
rect 8145 13905 8200 13921
rect 7969 13887 8010 13888
rect 7969 13858 8011 13887
rect 7981 13843 8011 13858
rect 8065 13843 8095 13905
rect 8163 13883 8193 13905
rect 9557 13897 9587 13937
rect 9641 14003 9671 14109
rect 10769 14223 10799 14249
rect 10869 14223 10899 14249
rect 10973 14223 11003 14249
rect 11059 14223 11089 14249
rect 11225 14223 11255 14249
rect 9749 14003 9779 14035
rect 9641 13987 9707 14003
rect 9641 13953 9657 13987
rect 9691 13953 9707 13987
rect 9641 13937 9707 13953
rect 9749 13987 9815 14003
rect 10769 13991 10799 14139
rect 10869 13991 10899 14139
rect 10973 13991 11003 14139
rect 11059 13991 11089 14139
rect 13029 14207 13059 14233
rect 12829 14183 12895 14193
rect 12829 14149 12845 14183
rect 12879 14149 12895 14183
rect 12829 14139 12895 14149
rect 12667 14091 12697 14117
rect 12763 14091 12793 14117
rect 12835 14091 12865 14139
rect 12931 14091 12961 14117
rect 11225 13991 11255 14023
rect 9749 13953 9765 13987
rect 9799 13953 9815 13987
rect 9749 13937 9815 13953
rect 10711 13975 10799 13991
rect 10711 13941 10721 13975
rect 10755 13941 10799 13975
rect 9641 13897 9671 13937
rect 9749 13915 9779 13937
rect 10711 13925 10799 13941
rect 7801 13733 7831 13759
rect 7897 13733 7927 13759
rect 7981 13733 8011 13759
rect 8065 13733 8095 13759
rect 9557 13787 9587 13813
rect 9641 13787 9671 13813
rect 10769 13857 10799 13925
rect 10857 13975 10911 13991
rect 10857 13941 10867 13975
rect 10901 13941 10911 13975
rect 10857 13925 10911 13941
rect 10963 13975 11017 13991
rect 10963 13941 10973 13975
rect 11007 13941 11017 13975
rect 10963 13925 11017 13941
rect 11059 13975 11123 13991
rect 11059 13941 11069 13975
rect 11103 13941 11123 13975
rect 11059 13925 11123 13941
rect 11170 13975 11255 13991
rect 12667 13975 12697 14007
rect 12763 13975 12793 14007
rect 11170 13941 11180 13975
rect 11214 13941 11255 13975
rect 11170 13925 11255 13941
rect 10857 13857 10887 13925
rect 10963 13857 10993 13925
rect 11059 13857 11089 13925
rect 11225 13903 11255 13925
rect 12613 13959 12697 13975
rect 12613 13925 12623 13959
rect 12657 13925 12697 13959
rect 12613 13909 12697 13925
rect 12739 13959 12793 13975
rect 12739 13925 12749 13959
rect 12783 13925 12793 13959
rect 12739 13909 12793 13925
rect 9749 13759 9779 13785
rect 11949 13849 11979 13875
rect 8163 13727 8193 13753
rect 10769 13747 10799 13773
rect 10857 13747 10887 13773
rect 10963 13747 10993 13773
rect 11059 13747 11089 13773
rect 11225 13747 11255 13773
rect 11780 13733 11810 13759
rect 11852 13733 11882 13759
rect 12667 13847 12697 13909
rect 12763 13847 12793 13909
rect 12835 13892 12865 14007
rect 12931 13975 12961 14007
rect 13029 13975 13059 14007
rect 12915 13959 12969 13975
rect 12915 13925 12925 13959
rect 12959 13925 12969 13959
rect 12915 13909 12969 13925
rect 13011 13959 13066 13975
rect 13011 13925 13021 13959
rect 13055 13925 13066 13959
rect 13011 13909 13066 13925
rect 12835 13891 12876 13892
rect 12835 13862 12877 13891
rect 12847 13847 12877 13862
rect 12931 13847 12961 13909
rect 13029 13887 13059 13909
rect 12667 13737 12697 13763
rect 12763 13737 12793 13763
rect 12847 13737 12877 13763
rect 12931 13737 12961 13763
rect 13029 13731 13059 13757
rect 6914 13613 6944 13645
rect 6844 13597 6944 13613
rect 6844 13563 6860 13597
rect 6894 13563 6944 13597
rect 6844 13547 6944 13563
rect 6986 13613 7016 13645
rect 7083 13613 7113 13645
rect 11780 13617 11810 13649
rect 6986 13597 7040 13613
rect 6986 13563 6996 13597
rect 7030 13563 7040 13597
rect 6986 13547 7040 13563
rect 7083 13597 7149 13613
rect 7083 13563 7099 13597
rect 7133 13563 7149 13597
rect 7083 13547 7149 13563
rect 11710 13601 11810 13617
rect 11710 13567 11726 13601
rect 11760 13567 11810 13601
rect 11710 13551 11810 13567
rect 11852 13617 11882 13649
rect 11949 13617 11979 13649
rect 11852 13601 11906 13617
rect 11852 13567 11862 13601
rect 11896 13567 11906 13601
rect 11852 13551 11906 13567
rect 11949 13601 12015 13617
rect 11949 13567 11965 13601
rect 11999 13567 12015 13601
rect 11949 13551 12015 13567
rect 6902 13479 6932 13547
rect 6986 13479 7016 13547
rect 7083 13525 7113 13547
rect 6299 13377 6329 13403
rect 11768 13483 11798 13551
rect 11852 13483 11882 13551
rect 11949 13529 11979 13551
rect 4557 13307 4587 13333
rect 4641 13307 4671 13333
rect 4725 13307 4755 13333
rect 4809 13307 4839 13333
rect 4997 13307 5027 13333
rect 6111 13356 6165 13372
rect 6111 13322 6121 13356
rect 6155 13322 6165 13356
rect 6111 13306 6165 13322
rect 6027 13264 6057 13305
rect 6111 13264 6141 13306
rect 6204 13264 6234 13290
rect 6027 13131 6057 13180
rect 6111 13162 6141 13180
rect 4557 13075 4587 13107
rect 4641 13075 4671 13107
rect 4725 13075 4755 13107
rect 4809 13075 4839 13107
rect 4997 13075 5027 13107
rect 4545 13059 4599 13075
rect 4545 13025 4555 13059
rect 4589 13025 4599 13059
rect 4545 13009 4599 13025
rect 4641 13059 4755 13075
rect 4641 13025 4672 13059
rect 4706 13025 4755 13059
rect 4641 13009 4755 13025
rect 4797 13059 4851 13075
rect 4797 13025 4807 13059
rect 4841 13025 4851 13059
rect 4797 13009 4851 13025
rect 4893 13059 5027 13075
rect 4893 13025 4903 13059
rect 4937 13042 5027 13059
rect 5973 13083 6057 13131
rect 5973 13049 5983 13083
rect 6017 13049 6057 13083
rect 4937 13025 5023 13042
rect 4893 13009 5023 13025
rect 4557 12987 4587 13009
rect 4641 12987 4671 13009
rect 4725 12987 4755 13009
rect 4809 12987 4839 13009
rect 4993 12987 5023 13009
rect 5973 13026 6057 13049
rect 6027 13011 6057 13026
rect 6099 13137 6141 13162
rect 6204 13139 6234 13180
rect 6902 13369 6932 13395
rect 6986 13369 7016 13395
rect 7083 13369 7113 13395
rect 11165 13381 11195 13407
rect 9423 13311 9453 13337
rect 9507 13311 9537 13337
rect 9591 13311 9621 13337
rect 9675 13311 9705 13337
rect 9863 13311 9893 13337
rect 6299 13145 6329 13177
rect 6099 13011 6129 13137
rect 6183 13123 6237 13139
rect 6183 13106 6193 13123
rect 6171 13089 6193 13106
rect 6227 13089 6237 13123
rect 6171 13073 6237 13089
rect 6279 13129 6333 13145
rect 6279 13095 6289 13129
rect 6323 13095 6333 13129
rect 10977 13360 11031 13376
rect 10977 13326 10987 13360
rect 11021 13326 11031 13360
rect 10977 13310 11031 13326
rect 10893 13268 10923 13309
rect 10977 13268 11007 13310
rect 11070 13268 11100 13294
rect 10893 13135 10923 13184
rect 10977 13166 11007 13184
rect 6279 13079 6333 13095
rect 9423 13079 9453 13111
rect 9507 13079 9537 13111
rect 9591 13079 9621 13111
rect 9675 13079 9705 13111
rect 9863 13079 9893 13111
rect 6171 13050 6213 13073
rect 6299 13057 6329 13079
rect 9411 13063 9465 13079
rect 6171 13026 6208 13050
rect 6171 13011 6201 13026
rect 9411 13029 9421 13063
rect 9455 13029 9465 13063
rect 9411 13013 9465 13029
rect 9507 13063 9621 13079
rect 9507 13029 9538 13063
rect 9572 13029 9621 13063
rect 9507 13013 9621 13029
rect 9663 13063 9717 13079
rect 9663 13029 9673 13063
rect 9707 13029 9717 13063
rect 9663 13013 9717 13029
rect 9759 13063 9893 13079
rect 9759 13029 9769 13063
rect 9803 13046 9893 13063
rect 10839 13087 10923 13135
rect 10839 13053 10849 13087
rect 10883 13053 10923 13087
rect 9803 13029 9889 13046
rect 9759 13013 9889 13029
rect 9423 12991 9453 13013
rect 9507 12991 9537 13013
rect 9591 12991 9621 13013
rect 9675 12991 9705 13013
rect 9859 12991 9889 13013
rect 10839 13030 10923 13053
rect 10893 13015 10923 13030
rect 10965 13141 11007 13166
rect 11070 13143 11100 13184
rect 11768 13373 11798 13399
rect 11852 13373 11882 13399
rect 11949 13373 11979 13399
rect 11165 13149 11195 13181
rect 10965 13015 10995 13141
rect 11049 13127 11103 13143
rect 11049 13110 11059 13127
rect 11037 13093 11059 13110
rect 11093 13093 11103 13127
rect 11037 13077 11103 13093
rect 11145 13133 11199 13149
rect 11145 13099 11155 13133
rect 11189 13099 11199 13133
rect 11145 13083 11199 13099
rect 11037 13054 11079 13077
rect 11165 13061 11195 13083
rect 11037 13030 11074 13054
rect 11037 13015 11067 13030
rect 6027 12901 6057 12927
rect 6099 12901 6129 12927
rect 6171 12901 6201 12927
rect 6299 12901 6329 12927
rect 10893 12905 10923 12931
rect 10965 12905 10995 12931
rect 11037 12905 11067 12931
rect 11165 12905 11195 12931
rect 4557 12831 4587 12857
rect 4641 12831 4671 12857
rect 4725 12831 4755 12857
rect 4809 12831 4839 12857
rect 4993 12831 5023 12857
rect 9423 12835 9453 12861
rect 9507 12835 9537 12861
rect 9591 12835 9621 12861
rect 9675 12835 9705 12861
rect 9859 12835 9889 12861
rect 4875 12563 4905 12589
rect 9741 12567 9771 12593
rect 4683 12521 4713 12547
rect 4767 12521 4797 12547
rect 4683 12331 4713 12437
rect 4626 12315 4713 12331
rect 4626 12281 4642 12315
rect 4676 12281 4713 12315
rect 4626 12265 4713 12281
rect 4683 12225 4713 12265
rect 4767 12331 4797 12437
rect 9549 12525 9579 12551
rect 9633 12525 9663 12551
rect 4875 12331 4905 12363
rect 6251 12357 6281 12383
rect 4767 12315 4833 12331
rect 4767 12281 4783 12315
rect 4817 12281 4833 12315
rect 4767 12265 4833 12281
rect 4875 12315 4941 12331
rect 4875 12281 4891 12315
rect 4925 12281 4941 12315
rect 4875 12265 4941 12281
rect 6059 12315 6089 12341
rect 6143 12315 6173 12341
rect 4767 12225 4797 12265
rect 4875 12243 4905 12265
rect 4683 12115 4713 12141
rect 4767 12115 4797 12141
rect 6059 12125 6089 12231
rect 4875 12087 4905 12113
rect 6002 12109 6089 12125
rect 6002 12075 6018 12109
rect 6052 12075 6089 12109
rect 6002 12059 6089 12075
rect 6059 12019 6089 12059
rect 6143 12125 6173 12231
rect 9549 12335 9579 12441
rect 9492 12319 9579 12335
rect 9492 12285 9508 12319
rect 9542 12285 9579 12319
rect 9492 12269 9579 12285
rect 9549 12229 9579 12269
rect 9633 12335 9663 12441
rect 9741 12335 9771 12367
rect 11117 12361 11147 12387
rect 9633 12319 9699 12335
rect 9633 12285 9649 12319
rect 9683 12285 9699 12319
rect 9633 12269 9699 12285
rect 9741 12319 9807 12335
rect 9741 12285 9757 12319
rect 9791 12285 9807 12319
rect 9741 12269 9807 12285
rect 10925 12319 10955 12345
rect 11009 12319 11039 12345
rect 9633 12229 9663 12269
rect 9741 12247 9771 12269
rect 6251 12125 6281 12157
rect 6143 12109 6209 12125
rect 6143 12075 6159 12109
rect 6193 12075 6209 12109
rect 6143 12059 6209 12075
rect 6251 12109 6317 12125
rect 9549 12119 9579 12145
rect 9633 12119 9663 12145
rect 10925 12129 10955 12235
rect 6251 12075 6267 12109
rect 6301 12075 6317 12109
rect 9741 12091 9771 12117
rect 10868 12113 10955 12129
rect 6251 12059 6317 12075
rect 10868 12079 10884 12113
rect 10918 12079 10955 12113
rect 10868 12063 10955 12079
rect 6143 12019 6173 12059
rect 6251 12037 6281 12059
rect 6059 11909 6089 11935
rect 6143 11909 6173 11935
rect 10925 12023 10955 12063
rect 11009 12129 11039 12235
rect 11117 12129 11147 12161
rect 11009 12113 11075 12129
rect 11009 12079 11025 12113
rect 11059 12079 11075 12113
rect 11009 12063 11075 12079
rect 11117 12113 11183 12129
rect 11117 12079 11133 12113
rect 11167 12079 11183 12113
rect 11117 12063 11183 12079
rect 11009 12023 11039 12063
rect 11117 12041 11147 12063
rect 10925 11913 10955 11939
rect 11009 11913 11039 11939
rect 6251 11881 6281 11907
rect 11117 11885 11147 11911
rect 4567 11743 4597 11769
rect 4651 11743 4681 11769
rect 4735 11743 4765 11769
rect 4819 11743 4849 11769
rect 5007 11743 5037 11769
rect 9433 11747 9463 11773
rect 9517 11747 9547 11773
rect 9601 11747 9631 11773
rect 9685 11747 9715 11773
rect 9873 11747 9903 11773
rect 4567 11511 4597 11543
rect 4651 11511 4681 11543
rect 4735 11511 4765 11543
rect 4819 11511 4849 11543
rect 5007 11511 5037 11543
rect 9433 11515 9463 11547
rect 9517 11515 9547 11547
rect 9601 11515 9631 11547
rect 9685 11515 9715 11547
rect 9873 11515 9903 11547
rect 4555 11495 4609 11511
rect 4555 11461 4565 11495
rect 4599 11461 4609 11495
rect 4555 11445 4609 11461
rect 4651 11495 4765 11511
rect 4651 11461 4682 11495
rect 4716 11461 4765 11495
rect 4651 11445 4765 11461
rect 4807 11495 4861 11511
rect 4807 11461 4817 11495
rect 4851 11461 4861 11495
rect 4807 11445 4861 11461
rect 4903 11495 5037 11511
rect 4903 11461 4913 11495
rect 4947 11478 5037 11495
rect 9421 11499 9475 11515
rect 4947 11461 5033 11478
rect 4903 11445 5033 11461
rect 9421 11465 9431 11499
rect 9465 11465 9475 11499
rect 9421 11449 9475 11465
rect 9517 11499 9631 11515
rect 9517 11465 9548 11499
rect 9582 11465 9631 11499
rect 9517 11449 9631 11465
rect 9673 11499 9727 11515
rect 9673 11465 9683 11499
rect 9717 11465 9727 11499
rect 9673 11449 9727 11465
rect 9769 11499 9903 11515
rect 9769 11465 9779 11499
rect 9813 11482 9903 11499
rect 9813 11465 9899 11482
rect 9769 11449 9899 11465
rect 4567 11423 4597 11445
rect 4651 11423 4681 11445
rect 4735 11423 4765 11445
rect 4819 11423 4849 11445
rect 5003 11423 5033 11445
rect 9433 11427 9463 11449
rect 9517 11427 9547 11449
rect 9601 11427 9631 11449
rect 9685 11427 9715 11449
rect 9869 11427 9899 11449
rect 4567 11267 4597 11293
rect 4651 11267 4681 11293
rect 4735 11267 4765 11293
rect 4819 11267 4849 11293
rect 5003 11267 5033 11293
rect 9433 11271 9463 11297
rect 9517 11271 9547 11297
rect 9601 11271 9631 11297
rect 9685 11271 9715 11297
rect 9869 11271 9899 11297
rect 4885 10999 4915 11025
rect 9751 11003 9781 11029
rect 4693 10957 4723 10983
rect 4777 10957 4807 10983
rect 4693 10767 4723 10873
rect 4636 10751 4723 10767
rect 4636 10717 4652 10751
rect 4686 10717 4723 10751
rect 4636 10701 4723 10717
rect 4693 10661 4723 10701
rect 4777 10767 4807 10873
rect 9559 10961 9589 10987
rect 9643 10961 9673 10987
rect 4885 10767 4915 10799
rect 9559 10771 9589 10877
rect 4777 10751 4843 10767
rect 4777 10717 4793 10751
rect 4827 10717 4843 10751
rect 4777 10701 4843 10717
rect 4885 10751 4951 10767
rect 4885 10717 4901 10751
rect 4935 10717 4951 10751
rect 4885 10701 4951 10717
rect 9502 10755 9589 10771
rect 9502 10721 9518 10755
rect 9552 10721 9589 10755
rect 9502 10705 9589 10721
rect 4777 10661 4807 10701
rect 4885 10679 4915 10701
rect 4693 10551 4723 10577
rect 4777 10551 4807 10577
rect 9559 10665 9589 10705
rect 9643 10771 9673 10877
rect 9751 10771 9781 10803
rect 9643 10755 9709 10771
rect 9643 10721 9659 10755
rect 9693 10721 9709 10755
rect 9643 10705 9709 10721
rect 9751 10755 9817 10771
rect 9751 10721 9767 10755
rect 9801 10721 9817 10755
rect 9751 10705 9817 10721
rect 9643 10665 9673 10705
rect 9751 10683 9781 10705
rect 9559 10555 9589 10581
rect 9643 10555 9673 10581
rect 4885 10523 4915 10549
rect 9751 10527 9781 10553
rect 6238 6553 6268 6579
rect 6238 6401 6268 6423
rect 6238 6385 6324 6401
rect 6238 6351 6274 6385
rect 6308 6351 6324 6385
rect 6238 6335 6324 6351
rect 6238 6303 6268 6335
rect 6238 6077 6268 6103
rect 10132 5921 10162 5947
rect 10231 5921 10261 5947
rect 10327 5921 10357 5947
rect 10399 5921 10429 5947
rect 10495 5921 10525 5947
rect 10584 5921 10614 5947
rect 10668 5921 10698 5947
rect 10752 5921 10782 5947
rect 10940 5921 10970 5947
rect 11024 5921 11054 5947
rect 11108 5921 11138 5947
rect 11192 5921 11222 5947
rect 11282 5921 11312 5947
rect 11381 5921 11411 5947
rect 10132 5769 10162 5791
rect 10231 5777 10261 5837
rect 10132 5753 10186 5769
rect 10132 5719 10142 5753
rect 10176 5719 10186 5753
rect 10132 5703 10186 5719
rect 10231 5761 10285 5777
rect 10231 5727 10241 5761
rect 10275 5727 10285 5761
rect 10231 5711 10285 5727
rect 10132 5671 10162 5703
rect 1950 5501 1980 5527
rect 2049 5501 2079 5527
rect 2145 5501 2175 5527
rect 2217 5501 2247 5527
rect 2313 5501 2343 5527
rect 2402 5501 2432 5527
rect 2486 5501 2516 5527
rect 2570 5501 2600 5527
rect 2758 5501 2788 5527
rect 2842 5501 2872 5527
rect 2926 5501 2956 5527
rect 3010 5501 3040 5527
rect 3100 5501 3130 5527
rect 3199 5501 3229 5527
rect 1950 5349 1980 5371
rect 2049 5357 2079 5417
rect 1950 5333 2004 5349
rect 1950 5299 1960 5333
rect 1994 5299 2004 5333
rect 1950 5283 2004 5299
rect 2049 5341 2103 5357
rect 2049 5307 2059 5341
rect 2093 5307 2103 5341
rect 2049 5291 2103 5307
rect 1950 5251 1980 5283
rect 2049 5135 2079 5291
rect 2145 5245 2175 5417
rect 2121 5229 2175 5245
rect 2121 5195 2131 5229
rect 2165 5195 2175 5229
rect 2121 5179 2175 5195
rect 2145 5135 2175 5179
rect 2217 5245 2247 5417
rect 2313 5373 2343 5417
rect 2402 5373 2432 5417
rect 2486 5402 2516 5417
rect 2289 5357 2343 5373
rect 2289 5323 2299 5357
rect 2333 5323 2343 5357
rect 2289 5307 2343 5323
rect 2389 5357 2443 5373
rect 2389 5323 2399 5357
rect 2433 5323 2443 5357
rect 2389 5307 2443 5323
rect 2485 5372 2516 5402
rect 2570 5402 2600 5417
rect 2758 5402 2788 5417
rect 2570 5372 2788 5402
rect 2217 5229 2271 5245
rect 2217 5195 2227 5229
rect 2261 5195 2271 5229
rect 2217 5179 2271 5195
rect 2217 5135 2247 5179
rect 2313 5135 2343 5307
rect 2402 5135 2432 5307
rect 2485 5261 2515 5372
rect 2570 5357 2611 5372
rect 2581 5261 2611 5357
rect 2842 5342 2872 5417
rect 2926 5343 2956 5417
rect 2818 5326 2872 5342
rect 2818 5292 2828 5326
rect 2862 5292 2872 5326
rect 2818 5276 2872 5292
rect 2914 5327 2968 5343
rect 2914 5293 2924 5327
rect 2958 5293 2968 5327
rect 2914 5277 2968 5293
rect 2474 5245 2528 5261
rect 2474 5211 2484 5245
rect 2518 5211 2528 5245
rect 2474 5195 2528 5211
rect 2581 5245 2645 5261
rect 2581 5211 2601 5245
rect 2635 5211 2645 5245
rect 2486 5135 2516 5195
rect 2581 5180 2645 5211
rect 2570 5150 2788 5180
rect 2570 5135 2600 5150
rect 2758 5135 2788 5150
rect 2842 5135 2872 5276
rect 2926 5135 2956 5277
rect 3010 5238 3040 5417
rect 3100 5349 3130 5417
rect 4084 5493 4114 5519
rect 4183 5493 4213 5519
rect 4279 5493 4309 5519
rect 4351 5493 4381 5519
rect 4447 5493 4477 5519
rect 4536 5493 4566 5519
rect 4620 5493 4650 5519
rect 4704 5493 4734 5519
rect 4892 5493 4922 5519
rect 4976 5493 5006 5519
rect 5060 5493 5090 5519
rect 5144 5493 5174 5519
rect 5234 5493 5264 5519
rect 5333 5493 5363 5519
rect 6036 5493 6066 5519
rect 6135 5493 6165 5519
rect 6231 5493 6261 5519
rect 6303 5493 6333 5519
rect 6399 5493 6429 5519
rect 6488 5493 6518 5519
rect 6572 5493 6602 5519
rect 6656 5493 6686 5519
rect 6844 5493 6874 5519
rect 6928 5493 6958 5519
rect 7012 5493 7042 5519
rect 7096 5493 7126 5519
rect 7186 5493 7216 5519
rect 7285 5493 7315 5519
rect 8038 5499 8068 5525
rect 8137 5499 8167 5525
rect 8233 5499 8263 5525
rect 8305 5499 8335 5525
rect 8401 5499 8431 5525
rect 8490 5499 8520 5525
rect 8574 5499 8604 5525
rect 8658 5499 8688 5525
rect 8846 5499 8876 5525
rect 8930 5499 8960 5525
rect 9014 5499 9044 5525
rect 9098 5499 9128 5525
rect 9188 5499 9218 5525
rect 9287 5499 9317 5525
rect 3199 5349 3229 5371
rect 3082 5333 3136 5349
rect 3082 5299 3092 5333
rect 3126 5299 3136 5333
rect 3082 5283 3136 5299
rect 3178 5333 3232 5349
rect 3178 5299 3188 5333
rect 3222 5299 3232 5333
rect 3178 5283 3232 5299
rect 4084 5341 4114 5363
rect 4183 5349 4213 5409
rect 4084 5325 4138 5341
rect 4084 5291 4094 5325
rect 4128 5291 4138 5325
rect 3004 5222 3058 5238
rect 3004 5188 3014 5222
rect 3048 5188 3058 5222
rect 3004 5172 3058 5188
rect 3010 5135 3040 5172
rect 3100 5135 3130 5283
rect 3199 5251 3229 5283
rect 4084 5275 4138 5291
rect 4183 5333 4237 5349
rect 4183 5299 4193 5333
rect 4227 5299 4237 5333
rect 4183 5283 4237 5299
rect 4084 5243 4114 5275
rect 1950 5025 1980 5051
rect 2049 5025 2079 5051
rect 2145 5025 2175 5051
rect 2217 5025 2247 5051
rect 2313 5025 2343 5051
rect 2402 5025 2432 5051
rect 2486 5025 2516 5051
rect 2570 5025 2600 5051
rect 2758 5025 2788 5051
rect 2842 5025 2872 5051
rect 2926 5025 2956 5051
rect 3010 5025 3040 5051
rect 3100 5025 3130 5051
rect 3199 5025 3229 5051
rect 4183 5127 4213 5283
rect 4279 5237 4309 5409
rect 4255 5221 4309 5237
rect 4255 5187 4265 5221
rect 4299 5187 4309 5221
rect 4255 5171 4309 5187
rect 4279 5127 4309 5171
rect 4351 5237 4381 5409
rect 4447 5365 4477 5409
rect 4536 5365 4566 5409
rect 4620 5394 4650 5409
rect 4423 5349 4477 5365
rect 4423 5315 4433 5349
rect 4467 5315 4477 5349
rect 4423 5299 4477 5315
rect 4523 5349 4577 5365
rect 4523 5315 4533 5349
rect 4567 5315 4577 5349
rect 4523 5299 4577 5315
rect 4619 5364 4650 5394
rect 4704 5394 4734 5409
rect 4892 5394 4922 5409
rect 4704 5364 4922 5394
rect 4351 5221 4405 5237
rect 4351 5187 4361 5221
rect 4395 5187 4405 5221
rect 4351 5171 4405 5187
rect 4351 5127 4381 5171
rect 4447 5127 4477 5299
rect 4536 5127 4566 5299
rect 4619 5253 4649 5364
rect 4704 5349 4745 5364
rect 4715 5253 4745 5349
rect 4976 5334 5006 5409
rect 5060 5335 5090 5409
rect 4952 5318 5006 5334
rect 4952 5284 4962 5318
rect 4996 5284 5006 5318
rect 4952 5268 5006 5284
rect 5048 5319 5102 5335
rect 5048 5285 5058 5319
rect 5092 5285 5102 5319
rect 5048 5269 5102 5285
rect 4608 5237 4662 5253
rect 4608 5203 4618 5237
rect 4652 5203 4662 5237
rect 4608 5187 4662 5203
rect 4715 5237 4779 5253
rect 4715 5203 4735 5237
rect 4769 5203 4779 5237
rect 4620 5127 4650 5187
rect 4715 5172 4779 5203
rect 4704 5142 4922 5172
rect 4704 5127 4734 5142
rect 4892 5127 4922 5142
rect 4976 5127 5006 5268
rect 5060 5127 5090 5269
rect 5144 5230 5174 5409
rect 5234 5341 5264 5409
rect 5333 5341 5363 5363
rect 6036 5341 6066 5363
rect 6135 5349 6165 5409
rect 5216 5325 5270 5341
rect 5216 5291 5226 5325
rect 5260 5291 5270 5325
rect 5216 5275 5270 5291
rect 5312 5325 5366 5341
rect 5312 5291 5322 5325
rect 5356 5291 5366 5325
rect 5312 5275 5366 5291
rect 6036 5325 6090 5341
rect 6036 5291 6046 5325
rect 6080 5291 6090 5325
rect 6036 5275 6090 5291
rect 6135 5333 6189 5349
rect 6135 5299 6145 5333
rect 6179 5299 6189 5333
rect 6135 5283 6189 5299
rect 5138 5214 5192 5230
rect 5138 5180 5148 5214
rect 5182 5180 5192 5214
rect 5138 5164 5192 5180
rect 5144 5127 5174 5164
rect 5234 5127 5264 5275
rect 5333 5243 5363 5275
rect 6036 5243 6066 5275
rect 6135 5127 6165 5283
rect 6231 5237 6261 5409
rect 6207 5221 6261 5237
rect 6207 5187 6217 5221
rect 6251 5187 6261 5221
rect 6207 5171 6261 5187
rect 6231 5127 6261 5171
rect 6303 5237 6333 5409
rect 6399 5365 6429 5409
rect 6488 5365 6518 5409
rect 6572 5394 6602 5409
rect 6375 5349 6429 5365
rect 6375 5315 6385 5349
rect 6419 5315 6429 5349
rect 6375 5299 6429 5315
rect 6475 5349 6529 5365
rect 6475 5315 6485 5349
rect 6519 5315 6529 5349
rect 6475 5299 6529 5315
rect 6571 5364 6602 5394
rect 6656 5394 6686 5409
rect 6844 5394 6874 5409
rect 6656 5364 6874 5394
rect 6303 5221 6357 5237
rect 6303 5187 6313 5221
rect 6347 5187 6357 5221
rect 6303 5171 6357 5187
rect 6303 5127 6333 5171
rect 6399 5127 6429 5299
rect 6488 5127 6518 5299
rect 6571 5253 6601 5364
rect 6656 5349 6697 5364
rect 6667 5253 6697 5349
rect 6928 5334 6958 5409
rect 7012 5335 7042 5409
rect 6904 5318 6958 5334
rect 6904 5284 6914 5318
rect 6948 5284 6958 5318
rect 6904 5268 6958 5284
rect 7000 5319 7054 5335
rect 7000 5285 7010 5319
rect 7044 5285 7054 5319
rect 7000 5269 7054 5285
rect 6560 5237 6614 5253
rect 6560 5203 6570 5237
rect 6604 5203 6614 5237
rect 6560 5187 6614 5203
rect 6667 5237 6731 5253
rect 6667 5203 6687 5237
rect 6721 5203 6731 5237
rect 6572 5127 6602 5187
rect 6667 5172 6731 5203
rect 6656 5142 6874 5172
rect 6656 5127 6686 5142
rect 6844 5127 6874 5142
rect 6928 5127 6958 5268
rect 7012 5127 7042 5269
rect 7096 5230 7126 5409
rect 7186 5341 7216 5409
rect 7285 5341 7315 5363
rect 8038 5347 8068 5369
rect 8137 5355 8167 5415
rect 7168 5325 7222 5341
rect 7168 5291 7178 5325
rect 7212 5291 7222 5325
rect 7168 5275 7222 5291
rect 7264 5325 7318 5341
rect 7264 5291 7274 5325
rect 7308 5291 7318 5325
rect 7264 5275 7318 5291
rect 8038 5331 8092 5347
rect 8038 5297 8048 5331
rect 8082 5297 8092 5331
rect 8038 5281 8092 5297
rect 8137 5339 8191 5355
rect 8137 5305 8147 5339
rect 8181 5305 8191 5339
rect 8137 5289 8191 5305
rect 7090 5214 7144 5230
rect 7090 5180 7100 5214
rect 7134 5180 7144 5214
rect 7090 5164 7144 5180
rect 7096 5127 7126 5164
rect 7186 5127 7216 5275
rect 7285 5243 7315 5275
rect 8038 5249 8068 5281
rect 8137 5133 8167 5289
rect 8233 5243 8263 5415
rect 8209 5227 8263 5243
rect 8209 5193 8219 5227
rect 8253 5193 8263 5227
rect 8209 5177 8263 5193
rect 8233 5133 8263 5177
rect 8305 5243 8335 5415
rect 8401 5371 8431 5415
rect 8490 5371 8520 5415
rect 8574 5400 8604 5415
rect 8377 5355 8431 5371
rect 8377 5321 8387 5355
rect 8421 5321 8431 5355
rect 8377 5305 8431 5321
rect 8477 5355 8531 5371
rect 8477 5321 8487 5355
rect 8521 5321 8531 5355
rect 8477 5305 8531 5321
rect 8573 5370 8604 5400
rect 8658 5400 8688 5415
rect 8846 5400 8876 5415
rect 8658 5370 8876 5400
rect 8305 5227 8359 5243
rect 8305 5193 8315 5227
rect 8349 5193 8359 5227
rect 8305 5177 8359 5193
rect 8305 5133 8335 5177
rect 8401 5133 8431 5305
rect 8490 5133 8520 5305
rect 8573 5259 8603 5370
rect 8658 5355 8699 5370
rect 8669 5259 8699 5355
rect 8930 5340 8960 5415
rect 9014 5341 9044 5415
rect 8906 5324 8960 5340
rect 8906 5290 8916 5324
rect 8950 5290 8960 5324
rect 8906 5274 8960 5290
rect 9002 5325 9056 5341
rect 9002 5291 9012 5325
rect 9046 5291 9056 5325
rect 9002 5275 9056 5291
rect 8562 5243 8616 5259
rect 8562 5209 8572 5243
rect 8606 5209 8616 5243
rect 8562 5193 8616 5209
rect 8669 5243 8733 5259
rect 8669 5209 8689 5243
rect 8723 5209 8733 5243
rect 8574 5133 8604 5193
rect 8669 5178 8733 5209
rect 8658 5148 8876 5178
rect 8658 5133 8688 5148
rect 8846 5133 8876 5148
rect 8930 5133 8960 5274
rect 9014 5133 9044 5275
rect 9098 5236 9128 5415
rect 9188 5347 9218 5415
rect 10231 5555 10261 5711
rect 10327 5665 10357 5837
rect 10303 5649 10357 5665
rect 10303 5615 10313 5649
rect 10347 5615 10357 5649
rect 10303 5599 10357 5615
rect 10327 5555 10357 5599
rect 10399 5665 10429 5837
rect 10495 5793 10525 5837
rect 10584 5793 10614 5837
rect 10668 5822 10698 5837
rect 10471 5777 10525 5793
rect 10471 5743 10481 5777
rect 10515 5743 10525 5777
rect 10471 5727 10525 5743
rect 10571 5777 10625 5793
rect 10571 5743 10581 5777
rect 10615 5743 10625 5777
rect 10571 5727 10625 5743
rect 10667 5792 10698 5822
rect 10752 5822 10782 5837
rect 10940 5822 10970 5837
rect 10752 5792 10970 5822
rect 10399 5649 10453 5665
rect 10399 5615 10409 5649
rect 10443 5615 10453 5649
rect 10399 5599 10453 5615
rect 10399 5555 10429 5599
rect 10495 5555 10525 5727
rect 10584 5555 10614 5727
rect 10667 5681 10697 5792
rect 10752 5777 10793 5792
rect 10763 5681 10793 5777
rect 11024 5762 11054 5837
rect 11108 5763 11138 5837
rect 11000 5746 11054 5762
rect 11000 5712 11010 5746
rect 11044 5712 11054 5746
rect 11000 5696 11054 5712
rect 11096 5747 11150 5763
rect 11096 5713 11106 5747
rect 11140 5713 11150 5747
rect 11096 5697 11150 5713
rect 10656 5665 10710 5681
rect 10656 5631 10666 5665
rect 10700 5631 10710 5665
rect 10656 5615 10710 5631
rect 10763 5665 10827 5681
rect 10763 5631 10783 5665
rect 10817 5631 10827 5665
rect 10668 5555 10698 5615
rect 10763 5600 10827 5631
rect 10752 5570 10970 5600
rect 10752 5555 10782 5570
rect 10940 5555 10970 5570
rect 11024 5555 11054 5696
rect 11108 5555 11138 5697
rect 11192 5658 11222 5837
rect 11282 5769 11312 5837
rect 12194 5909 12224 5935
rect 12293 5909 12323 5935
rect 12389 5909 12419 5935
rect 12461 5909 12491 5935
rect 12557 5909 12587 5935
rect 12646 5909 12676 5935
rect 12730 5909 12760 5935
rect 12814 5909 12844 5935
rect 13002 5909 13032 5935
rect 13086 5909 13116 5935
rect 13170 5909 13200 5935
rect 13254 5909 13284 5935
rect 13344 5909 13374 5935
rect 13443 5909 13473 5935
rect 14152 5917 14182 5943
rect 14251 5917 14281 5943
rect 14347 5917 14377 5943
rect 14419 5917 14449 5943
rect 14515 5917 14545 5943
rect 14604 5917 14634 5943
rect 14688 5917 14718 5943
rect 14772 5917 14802 5943
rect 14960 5917 14990 5943
rect 15044 5917 15074 5943
rect 15128 5917 15158 5943
rect 15212 5917 15242 5943
rect 15302 5917 15332 5943
rect 15401 5917 15431 5943
rect 16146 5923 16176 5949
rect 16245 5923 16275 5949
rect 16341 5923 16371 5949
rect 16413 5923 16443 5949
rect 16509 5923 16539 5949
rect 16598 5923 16628 5949
rect 16682 5923 16712 5949
rect 16766 5923 16796 5949
rect 16954 5923 16984 5949
rect 17038 5923 17068 5949
rect 17122 5923 17152 5949
rect 17206 5923 17236 5949
rect 17296 5923 17326 5949
rect 17395 5923 17425 5949
rect 11381 5769 11411 5791
rect 11264 5753 11318 5769
rect 11264 5719 11274 5753
rect 11308 5719 11318 5753
rect 11264 5703 11318 5719
rect 11360 5753 11414 5769
rect 11360 5719 11370 5753
rect 11404 5719 11414 5753
rect 11360 5703 11414 5719
rect 12194 5757 12224 5779
rect 12293 5765 12323 5825
rect 12194 5741 12248 5757
rect 12194 5707 12204 5741
rect 12238 5707 12248 5741
rect 11186 5642 11240 5658
rect 11186 5608 11196 5642
rect 11230 5608 11240 5642
rect 11186 5592 11240 5608
rect 11192 5555 11222 5592
rect 11282 5555 11312 5703
rect 11381 5671 11411 5703
rect 12194 5691 12248 5707
rect 12293 5749 12347 5765
rect 12293 5715 12303 5749
rect 12337 5715 12347 5749
rect 12293 5699 12347 5715
rect 12194 5659 12224 5691
rect 10132 5445 10162 5471
rect 10231 5445 10261 5471
rect 10327 5445 10357 5471
rect 10399 5445 10429 5471
rect 10495 5445 10525 5471
rect 10584 5445 10614 5471
rect 10668 5445 10698 5471
rect 10752 5445 10782 5471
rect 10940 5445 10970 5471
rect 11024 5445 11054 5471
rect 11108 5445 11138 5471
rect 11192 5445 11222 5471
rect 11282 5445 11312 5471
rect 11381 5445 11411 5471
rect 12293 5543 12323 5699
rect 12389 5653 12419 5825
rect 12365 5637 12419 5653
rect 12365 5603 12375 5637
rect 12409 5603 12419 5637
rect 12365 5587 12419 5603
rect 12389 5543 12419 5587
rect 12461 5653 12491 5825
rect 12557 5781 12587 5825
rect 12646 5781 12676 5825
rect 12730 5810 12760 5825
rect 12533 5765 12587 5781
rect 12533 5731 12543 5765
rect 12577 5731 12587 5765
rect 12533 5715 12587 5731
rect 12633 5765 12687 5781
rect 12633 5731 12643 5765
rect 12677 5731 12687 5765
rect 12633 5715 12687 5731
rect 12729 5780 12760 5810
rect 12814 5810 12844 5825
rect 13002 5810 13032 5825
rect 12814 5780 13032 5810
rect 12461 5637 12515 5653
rect 12461 5603 12471 5637
rect 12505 5603 12515 5637
rect 12461 5587 12515 5603
rect 12461 5543 12491 5587
rect 12557 5543 12587 5715
rect 12646 5543 12676 5715
rect 12729 5669 12759 5780
rect 12814 5765 12855 5780
rect 12825 5669 12855 5765
rect 13086 5750 13116 5825
rect 13170 5751 13200 5825
rect 13062 5734 13116 5750
rect 13062 5700 13072 5734
rect 13106 5700 13116 5734
rect 13062 5684 13116 5700
rect 13158 5735 13212 5751
rect 13158 5701 13168 5735
rect 13202 5701 13212 5735
rect 13158 5685 13212 5701
rect 12718 5653 12772 5669
rect 12718 5619 12728 5653
rect 12762 5619 12772 5653
rect 12718 5603 12772 5619
rect 12825 5653 12889 5669
rect 12825 5619 12845 5653
rect 12879 5619 12889 5653
rect 12730 5543 12760 5603
rect 12825 5588 12889 5619
rect 12814 5558 13032 5588
rect 12814 5543 12844 5558
rect 13002 5543 13032 5558
rect 13086 5543 13116 5684
rect 13170 5543 13200 5685
rect 13254 5646 13284 5825
rect 13344 5757 13374 5825
rect 13443 5757 13473 5779
rect 14152 5765 14182 5787
rect 14251 5773 14281 5833
rect 13326 5741 13380 5757
rect 13326 5707 13336 5741
rect 13370 5707 13380 5741
rect 13326 5691 13380 5707
rect 13422 5741 13476 5757
rect 13422 5707 13432 5741
rect 13466 5707 13476 5741
rect 13422 5691 13476 5707
rect 14152 5749 14206 5765
rect 14152 5715 14162 5749
rect 14196 5715 14206 5749
rect 14152 5699 14206 5715
rect 14251 5757 14305 5773
rect 14251 5723 14261 5757
rect 14295 5723 14305 5757
rect 14251 5707 14305 5723
rect 13248 5630 13302 5646
rect 13248 5596 13258 5630
rect 13292 5596 13302 5630
rect 13248 5580 13302 5596
rect 13254 5543 13284 5580
rect 13344 5543 13374 5691
rect 13443 5659 13473 5691
rect 14152 5667 14182 5699
rect 14251 5551 14281 5707
rect 14347 5661 14377 5833
rect 14323 5645 14377 5661
rect 14323 5611 14333 5645
rect 14367 5611 14377 5645
rect 14323 5595 14377 5611
rect 14347 5551 14377 5595
rect 14419 5661 14449 5833
rect 14515 5789 14545 5833
rect 14604 5789 14634 5833
rect 14688 5818 14718 5833
rect 14491 5773 14545 5789
rect 14491 5739 14501 5773
rect 14535 5739 14545 5773
rect 14491 5723 14545 5739
rect 14591 5773 14645 5789
rect 14591 5739 14601 5773
rect 14635 5739 14645 5773
rect 14591 5723 14645 5739
rect 14687 5788 14718 5818
rect 14772 5818 14802 5833
rect 14960 5818 14990 5833
rect 14772 5788 14990 5818
rect 14419 5645 14473 5661
rect 14419 5611 14429 5645
rect 14463 5611 14473 5645
rect 14419 5595 14473 5611
rect 14419 5551 14449 5595
rect 14515 5551 14545 5723
rect 14604 5551 14634 5723
rect 14687 5677 14717 5788
rect 14772 5773 14813 5788
rect 14783 5677 14813 5773
rect 15044 5758 15074 5833
rect 15128 5759 15158 5833
rect 15020 5742 15074 5758
rect 15020 5708 15030 5742
rect 15064 5708 15074 5742
rect 15020 5692 15074 5708
rect 15116 5743 15170 5759
rect 15116 5709 15126 5743
rect 15160 5709 15170 5743
rect 15116 5693 15170 5709
rect 14676 5661 14730 5677
rect 14676 5627 14686 5661
rect 14720 5627 14730 5661
rect 14676 5611 14730 5627
rect 14783 5661 14847 5677
rect 14783 5627 14803 5661
rect 14837 5627 14847 5661
rect 14688 5551 14718 5611
rect 14783 5596 14847 5627
rect 14772 5566 14990 5596
rect 14772 5551 14802 5566
rect 14960 5551 14990 5566
rect 15044 5551 15074 5692
rect 15128 5551 15158 5693
rect 15212 5654 15242 5833
rect 15302 5765 15332 5833
rect 15401 5765 15431 5787
rect 16146 5771 16176 5793
rect 16245 5779 16275 5839
rect 15284 5749 15338 5765
rect 15284 5715 15294 5749
rect 15328 5715 15338 5749
rect 15284 5699 15338 5715
rect 15380 5749 15434 5765
rect 15380 5715 15390 5749
rect 15424 5715 15434 5749
rect 15380 5699 15434 5715
rect 16146 5755 16200 5771
rect 16146 5721 16156 5755
rect 16190 5721 16200 5755
rect 16146 5705 16200 5721
rect 16245 5763 16299 5779
rect 16245 5729 16255 5763
rect 16289 5729 16299 5763
rect 16245 5713 16299 5729
rect 15206 5638 15260 5654
rect 15206 5604 15216 5638
rect 15250 5604 15260 5638
rect 15206 5588 15260 5604
rect 15212 5551 15242 5588
rect 15302 5551 15332 5699
rect 15401 5667 15431 5699
rect 16146 5673 16176 5705
rect 16245 5557 16275 5713
rect 16341 5667 16371 5839
rect 16317 5651 16371 5667
rect 16317 5617 16327 5651
rect 16361 5617 16371 5651
rect 16317 5601 16371 5617
rect 16341 5557 16371 5601
rect 16413 5667 16443 5839
rect 16509 5795 16539 5839
rect 16598 5795 16628 5839
rect 16682 5824 16712 5839
rect 16485 5779 16539 5795
rect 16485 5745 16495 5779
rect 16529 5745 16539 5779
rect 16485 5729 16539 5745
rect 16585 5779 16639 5795
rect 16585 5745 16595 5779
rect 16629 5745 16639 5779
rect 16585 5729 16639 5745
rect 16681 5794 16712 5824
rect 16766 5824 16796 5839
rect 16954 5824 16984 5839
rect 16766 5794 16984 5824
rect 16413 5651 16467 5667
rect 16413 5617 16423 5651
rect 16457 5617 16467 5651
rect 16413 5601 16467 5617
rect 16413 5557 16443 5601
rect 16509 5557 16539 5729
rect 16598 5557 16628 5729
rect 16681 5683 16711 5794
rect 16766 5779 16807 5794
rect 16777 5683 16807 5779
rect 17038 5764 17068 5839
rect 17122 5765 17152 5839
rect 17014 5748 17068 5764
rect 17014 5714 17024 5748
rect 17058 5714 17068 5748
rect 17014 5698 17068 5714
rect 17110 5749 17164 5765
rect 17110 5715 17120 5749
rect 17154 5715 17164 5749
rect 17110 5699 17164 5715
rect 16670 5667 16724 5683
rect 16670 5633 16680 5667
rect 16714 5633 16724 5667
rect 16670 5617 16724 5633
rect 16777 5667 16841 5683
rect 16777 5633 16797 5667
rect 16831 5633 16841 5667
rect 16682 5557 16712 5617
rect 16777 5602 16841 5633
rect 16766 5572 16984 5602
rect 16766 5557 16796 5572
rect 16954 5557 16984 5572
rect 17038 5557 17068 5698
rect 17122 5557 17152 5699
rect 17206 5660 17236 5839
rect 17296 5771 17326 5839
rect 17395 5771 17425 5793
rect 17278 5755 17332 5771
rect 17278 5721 17288 5755
rect 17322 5721 17332 5755
rect 17278 5705 17332 5721
rect 17374 5755 17428 5771
rect 17374 5721 17384 5755
rect 17418 5721 17428 5755
rect 17374 5705 17428 5721
rect 17200 5644 17254 5660
rect 17200 5610 17210 5644
rect 17244 5610 17254 5644
rect 17200 5594 17254 5610
rect 17206 5557 17236 5594
rect 17296 5557 17326 5705
rect 17395 5673 17425 5705
rect 12194 5433 12224 5459
rect 12293 5433 12323 5459
rect 12389 5433 12419 5459
rect 12461 5433 12491 5459
rect 12557 5433 12587 5459
rect 12646 5433 12676 5459
rect 12730 5433 12760 5459
rect 12814 5433 12844 5459
rect 13002 5433 13032 5459
rect 13086 5433 13116 5459
rect 13170 5433 13200 5459
rect 13254 5433 13284 5459
rect 13344 5433 13374 5459
rect 13443 5433 13473 5459
rect 14152 5441 14182 5467
rect 14251 5441 14281 5467
rect 14347 5441 14377 5467
rect 14419 5441 14449 5467
rect 14515 5441 14545 5467
rect 14604 5441 14634 5467
rect 14688 5441 14718 5467
rect 14772 5441 14802 5467
rect 14960 5441 14990 5467
rect 15044 5441 15074 5467
rect 15128 5441 15158 5467
rect 15212 5441 15242 5467
rect 15302 5441 15332 5467
rect 15401 5441 15431 5467
rect 16146 5447 16176 5473
rect 16245 5447 16275 5473
rect 16341 5447 16371 5473
rect 16413 5447 16443 5473
rect 16509 5447 16539 5473
rect 16598 5447 16628 5473
rect 16682 5447 16712 5473
rect 16766 5447 16796 5473
rect 16954 5447 16984 5473
rect 17038 5447 17068 5473
rect 17122 5447 17152 5473
rect 17206 5447 17236 5473
rect 17296 5447 17326 5473
rect 17395 5447 17425 5473
rect 9287 5347 9317 5369
rect 18427 5349 18457 5375
rect 18595 5349 18625 5375
rect 18691 5349 18721 5375
rect 18816 5349 18846 5375
rect 18912 5349 18942 5375
rect 19021 5349 19051 5375
rect 9170 5331 9224 5347
rect 9170 5297 9180 5331
rect 9214 5297 9224 5331
rect 9170 5281 9224 5297
rect 9266 5331 9320 5347
rect 9266 5297 9276 5331
rect 9310 5297 9320 5331
rect 9266 5281 9320 5297
rect 9092 5220 9146 5236
rect 9092 5186 9102 5220
rect 9136 5186 9146 5220
rect 9092 5170 9146 5186
rect 9098 5133 9128 5170
rect 9188 5133 9218 5281
rect 9287 5249 9317 5281
rect 18427 5120 18457 5265
rect 18595 5227 18625 5265
rect 18691 5233 18721 5265
rect 18816 5233 18846 5265
rect 18499 5217 18625 5227
rect 18499 5183 18515 5217
rect 18549 5197 18625 5217
rect 18667 5217 18721 5233
rect 18549 5183 18565 5197
rect 18499 5173 18565 5183
rect 18667 5183 18677 5217
rect 18711 5183 18721 5217
rect 18427 5104 18481 5120
rect 4084 5017 4114 5043
rect 4183 5017 4213 5043
rect 4279 5017 4309 5043
rect 4351 5017 4381 5043
rect 4447 5017 4477 5043
rect 4536 5017 4566 5043
rect 4620 5017 4650 5043
rect 4704 5017 4734 5043
rect 4892 5017 4922 5043
rect 4976 5017 5006 5043
rect 5060 5017 5090 5043
rect 5144 5017 5174 5043
rect 5234 5017 5264 5043
rect 5333 5017 5363 5043
rect 6036 5017 6066 5043
rect 6135 5017 6165 5043
rect 6231 5017 6261 5043
rect 6303 5017 6333 5043
rect 6399 5017 6429 5043
rect 6488 5017 6518 5043
rect 6572 5017 6602 5043
rect 6656 5017 6686 5043
rect 6844 5017 6874 5043
rect 6928 5017 6958 5043
rect 7012 5017 7042 5043
rect 7096 5017 7126 5043
rect 7186 5017 7216 5043
rect 7285 5017 7315 5043
rect 8038 5023 8068 5049
rect 8137 5023 8167 5049
rect 8233 5023 8263 5049
rect 8305 5023 8335 5049
rect 8401 5023 8431 5049
rect 8490 5023 8520 5049
rect 8574 5023 8604 5049
rect 8658 5023 8688 5049
rect 8846 5023 8876 5049
rect 8930 5023 8960 5049
rect 9014 5023 9044 5049
rect 9098 5023 9128 5049
rect 9188 5023 9218 5049
rect 9287 5023 9317 5049
rect 10160 5047 10190 5073
rect 10259 5047 10289 5073
rect 10355 5047 10385 5073
rect 10427 5047 10457 5073
rect 10523 5047 10553 5073
rect 10612 5047 10642 5073
rect 10696 5047 10726 5073
rect 10780 5047 10810 5073
rect 10968 5047 10998 5073
rect 11052 5047 11082 5073
rect 11136 5047 11166 5073
rect 11220 5047 11250 5073
rect 11310 5047 11340 5073
rect 11409 5047 11439 5073
rect 18427 5070 18437 5104
rect 18471 5070 18481 5104
rect 18427 5054 18481 5070
rect 10160 4895 10190 4917
rect 10259 4903 10289 4963
rect 10160 4879 10214 4895
rect 10160 4845 10170 4879
rect 10204 4845 10214 4879
rect 10160 4829 10214 4845
rect 10259 4887 10313 4903
rect 10259 4853 10269 4887
rect 10303 4853 10313 4887
rect 10259 4837 10313 4853
rect 10160 4797 10190 4829
rect 10259 4681 10289 4837
rect 10355 4791 10385 4963
rect 10331 4775 10385 4791
rect 10331 4741 10341 4775
rect 10375 4741 10385 4775
rect 10331 4725 10385 4741
rect 10355 4681 10385 4725
rect 10427 4791 10457 4963
rect 10523 4919 10553 4963
rect 10612 4919 10642 4963
rect 10696 4948 10726 4963
rect 10499 4903 10553 4919
rect 10499 4869 10509 4903
rect 10543 4869 10553 4903
rect 10499 4853 10553 4869
rect 10599 4903 10653 4919
rect 10599 4869 10609 4903
rect 10643 4869 10653 4903
rect 10599 4853 10653 4869
rect 10695 4918 10726 4948
rect 10780 4948 10810 4963
rect 10968 4948 10998 4963
rect 10780 4918 10998 4948
rect 10427 4775 10481 4791
rect 10427 4741 10437 4775
rect 10471 4741 10481 4775
rect 10427 4725 10481 4741
rect 10427 4681 10457 4725
rect 10523 4681 10553 4853
rect 10612 4681 10642 4853
rect 10695 4807 10725 4918
rect 10780 4903 10821 4918
rect 10791 4807 10821 4903
rect 11052 4888 11082 4963
rect 11136 4889 11166 4963
rect 11028 4872 11082 4888
rect 11028 4838 11038 4872
rect 11072 4838 11082 4872
rect 11028 4822 11082 4838
rect 11124 4873 11178 4889
rect 11124 4839 11134 4873
rect 11168 4839 11178 4873
rect 11124 4823 11178 4839
rect 10684 4791 10738 4807
rect 10684 4757 10694 4791
rect 10728 4757 10738 4791
rect 10684 4741 10738 4757
rect 10791 4791 10855 4807
rect 10791 4757 10811 4791
rect 10845 4757 10855 4791
rect 10696 4681 10726 4741
rect 10791 4726 10855 4757
rect 10780 4696 10998 4726
rect 10780 4681 10810 4696
rect 10968 4681 10998 4696
rect 11052 4681 11082 4822
rect 11136 4681 11166 4823
rect 11220 4784 11250 4963
rect 11310 4895 11340 4963
rect 12430 5003 12460 5029
rect 12529 5003 12559 5029
rect 12625 5003 12655 5029
rect 12697 5003 12727 5029
rect 12793 5003 12823 5029
rect 12882 5003 12912 5029
rect 12966 5003 12996 5029
rect 13050 5003 13080 5029
rect 13238 5003 13268 5029
rect 13322 5003 13352 5029
rect 13406 5003 13436 5029
rect 13490 5003 13520 5029
rect 13580 5003 13610 5029
rect 13679 5003 13709 5029
rect 11409 4895 11439 4917
rect 11292 4879 11346 4895
rect 11292 4845 11302 4879
rect 11336 4845 11346 4879
rect 11292 4829 11346 4845
rect 11388 4879 11442 4895
rect 11388 4845 11398 4879
rect 11432 4845 11442 4879
rect 11388 4829 11442 4845
rect 12430 4851 12460 4873
rect 12529 4859 12559 4919
rect 12430 4835 12484 4851
rect 11214 4768 11268 4784
rect 11214 4734 11224 4768
rect 11258 4734 11268 4768
rect 11214 4718 11268 4734
rect 11220 4681 11250 4718
rect 11310 4681 11340 4829
rect 11409 4797 11439 4829
rect 12430 4801 12440 4835
rect 12474 4801 12484 4835
rect 12430 4785 12484 4801
rect 12529 4843 12583 4859
rect 12529 4809 12539 4843
rect 12573 4809 12583 4843
rect 12529 4793 12583 4809
rect 12430 4753 12460 4785
rect 10160 4571 10190 4597
rect 10259 4571 10289 4597
rect 10355 4571 10385 4597
rect 10427 4571 10457 4597
rect 10523 4571 10553 4597
rect 10612 4571 10642 4597
rect 10696 4571 10726 4597
rect 10780 4571 10810 4597
rect 10968 4571 10998 4597
rect 11052 4571 11082 4597
rect 11136 4571 11166 4597
rect 11220 4571 11250 4597
rect 11310 4571 11340 4597
rect 11409 4571 11439 4597
rect 12529 4637 12559 4793
rect 12625 4747 12655 4919
rect 12601 4731 12655 4747
rect 12601 4697 12611 4731
rect 12645 4697 12655 4731
rect 12601 4681 12655 4697
rect 12625 4637 12655 4681
rect 12697 4747 12727 4919
rect 12793 4875 12823 4919
rect 12882 4875 12912 4919
rect 12966 4904 12996 4919
rect 12769 4859 12823 4875
rect 12769 4825 12779 4859
rect 12813 4825 12823 4859
rect 12769 4809 12823 4825
rect 12869 4859 12923 4875
rect 12869 4825 12879 4859
rect 12913 4825 12923 4859
rect 12869 4809 12923 4825
rect 12965 4874 12996 4904
rect 13050 4904 13080 4919
rect 13238 4904 13268 4919
rect 13050 4874 13268 4904
rect 12697 4731 12751 4747
rect 12697 4697 12707 4731
rect 12741 4697 12751 4731
rect 12697 4681 12751 4697
rect 12697 4637 12727 4681
rect 12793 4637 12823 4809
rect 12882 4637 12912 4809
rect 12965 4763 12995 4874
rect 13050 4859 13091 4874
rect 13061 4763 13091 4859
rect 13322 4844 13352 4919
rect 13406 4845 13436 4919
rect 13298 4828 13352 4844
rect 13298 4794 13308 4828
rect 13342 4794 13352 4828
rect 13298 4778 13352 4794
rect 13394 4829 13448 4845
rect 13394 4795 13404 4829
rect 13438 4795 13448 4829
rect 13394 4779 13448 4795
rect 12954 4747 13008 4763
rect 12954 4713 12964 4747
rect 12998 4713 13008 4747
rect 12954 4697 13008 4713
rect 13061 4747 13125 4763
rect 13061 4713 13081 4747
rect 13115 4713 13125 4747
rect 12966 4637 12996 4697
rect 13061 4682 13125 4713
rect 13050 4652 13268 4682
rect 13050 4637 13080 4652
rect 13238 4637 13268 4652
rect 13322 4637 13352 4778
rect 13406 4637 13436 4779
rect 13490 4740 13520 4919
rect 13580 4851 13610 4919
rect 14432 4997 14462 5023
rect 14531 4997 14561 5023
rect 14627 4997 14657 5023
rect 14699 4997 14729 5023
rect 14795 4997 14825 5023
rect 14884 4997 14914 5023
rect 14968 4997 14998 5023
rect 15052 4997 15082 5023
rect 15240 4997 15270 5023
rect 15324 4997 15354 5023
rect 15408 4997 15438 5023
rect 15492 4997 15522 5023
rect 15582 4997 15612 5023
rect 15681 4997 15711 5023
rect 18427 5022 18457 5054
rect 18523 5022 18553 5173
rect 18667 5167 18721 5183
rect 18763 5217 18846 5233
rect 18763 5183 18773 5217
rect 18807 5183 18846 5217
rect 18912 5197 18942 5265
rect 19021 5197 19051 5219
rect 18763 5167 18846 5183
rect 18904 5181 18958 5197
rect 18595 5104 18649 5120
rect 18595 5070 18605 5104
rect 18639 5070 18649 5104
rect 18595 5054 18649 5070
rect 18691 5067 18721 5167
rect 18904 5147 18914 5181
rect 18948 5147 18958 5181
rect 18904 5131 18958 5147
rect 19000 5181 19054 5197
rect 19000 5147 19010 5181
rect 19044 5147 19054 5181
rect 19000 5131 19054 5147
rect 18595 5022 18625 5054
rect 18691 5037 18839 5067
rect 18809 5022 18839 5037
rect 18912 5022 18942 5131
rect 19021 5099 19051 5131
rect 13679 4851 13709 4873
rect 13562 4835 13616 4851
rect 13562 4801 13572 4835
rect 13606 4801 13616 4835
rect 13562 4785 13616 4801
rect 13658 4835 13712 4851
rect 13658 4801 13668 4835
rect 13702 4801 13712 4835
rect 13658 4785 13712 4801
rect 14432 4845 14462 4867
rect 14531 4853 14561 4913
rect 14432 4829 14486 4845
rect 14432 4795 14442 4829
rect 14476 4795 14486 4829
rect 13484 4724 13538 4740
rect 13484 4690 13494 4724
rect 13528 4690 13538 4724
rect 13484 4674 13538 4690
rect 13490 4637 13520 4674
rect 13580 4637 13610 4785
rect 13679 4753 13709 4785
rect 14432 4779 14486 4795
rect 14531 4837 14585 4853
rect 14531 4803 14541 4837
rect 14575 4803 14585 4837
rect 14531 4787 14585 4803
rect 14432 4747 14462 4779
rect 12430 4527 12460 4553
rect 12529 4527 12559 4553
rect 12625 4527 12655 4553
rect 12697 4527 12727 4553
rect 12793 4527 12823 4553
rect 12882 4527 12912 4553
rect 12966 4527 12996 4553
rect 13050 4527 13080 4553
rect 13238 4527 13268 4553
rect 13322 4527 13352 4553
rect 13406 4527 13436 4553
rect 13490 4527 13520 4553
rect 13580 4527 13610 4553
rect 13679 4527 13709 4553
rect 14531 4631 14561 4787
rect 14627 4741 14657 4913
rect 14603 4725 14657 4741
rect 14603 4691 14613 4725
rect 14647 4691 14657 4725
rect 14603 4675 14657 4691
rect 14627 4631 14657 4675
rect 14699 4741 14729 4913
rect 14795 4869 14825 4913
rect 14884 4869 14914 4913
rect 14968 4898 14998 4913
rect 14771 4853 14825 4869
rect 14771 4819 14781 4853
rect 14815 4819 14825 4853
rect 14771 4803 14825 4819
rect 14871 4853 14925 4869
rect 14871 4819 14881 4853
rect 14915 4819 14925 4853
rect 14871 4803 14925 4819
rect 14967 4868 14998 4898
rect 15052 4898 15082 4913
rect 15240 4898 15270 4913
rect 15052 4868 15270 4898
rect 14699 4725 14753 4741
rect 14699 4691 14709 4725
rect 14743 4691 14753 4725
rect 14699 4675 14753 4691
rect 14699 4631 14729 4675
rect 14795 4631 14825 4803
rect 14884 4631 14914 4803
rect 14967 4757 14997 4868
rect 15052 4853 15093 4868
rect 15063 4757 15093 4853
rect 15324 4838 15354 4913
rect 15408 4839 15438 4913
rect 15300 4822 15354 4838
rect 15300 4788 15310 4822
rect 15344 4788 15354 4822
rect 15300 4772 15354 4788
rect 15396 4823 15450 4839
rect 15396 4789 15406 4823
rect 15440 4789 15450 4823
rect 15396 4773 15450 4789
rect 14956 4741 15010 4757
rect 14956 4707 14966 4741
rect 15000 4707 15010 4741
rect 14956 4691 15010 4707
rect 15063 4741 15127 4757
rect 15063 4707 15083 4741
rect 15117 4707 15127 4741
rect 14968 4631 14998 4691
rect 15063 4676 15127 4707
rect 15052 4646 15270 4676
rect 15052 4631 15082 4646
rect 15240 4631 15270 4646
rect 15324 4631 15354 4772
rect 15408 4631 15438 4773
rect 15492 4734 15522 4913
rect 15582 4845 15612 4913
rect 16454 4979 16484 5005
rect 16553 4979 16583 5005
rect 16649 4979 16679 5005
rect 16721 4979 16751 5005
rect 16817 4979 16847 5005
rect 16906 4979 16936 5005
rect 16990 4979 17020 5005
rect 17074 4979 17104 5005
rect 17262 4979 17292 5005
rect 17346 4979 17376 5005
rect 17430 4979 17460 5005
rect 17514 4979 17544 5005
rect 17604 4979 17634 5005
rect 17703 4979 17733 5005
rect 15681 4845 15711 4867
rect 15564 4829 15618 4845
rect 15564 4795 15574 4829
rect 15608 4795 15618 4829
rect 15564 4779 15618 4795
rect 15660 4829 15714 4845
rect 15660 4795 15670 4829
rect 15704 4795 15714 4829
rect 15660 4779 15714 4795
rect 16454 4827 16484 4849
rect 16553 4835 16583 4895
rect 16454 4811 16508 4827
rect 15486 4718 15540 4734
rect 15486 4684 15496 4718
rect 15530 4684 15540 4718
rect 15486 4668 15540 4684
rect 15492 4631 15522 4668
rect 15582 4631 15612 4779
rect 15681 4747 15711 4779
rect 16454 4777 16464 4811
rect 16498 4777 16508 4811
rect 16454 4761 16508 4777
rect 16553 4819 16607 4835
rect 16553 4785 16563 4819
rect 16597 4785 16607 4819
rect 16553 4769 16607 4785
rect 16454 4729 16484 4761
rect 14432 4521 14462 4547
rect 14531 4521 14561 4547
rect 14627 4521 14657 4547
rect 14699 4521 14729 4547
rect 14795 4521 14825 4547
rect 14884 4521 14914 4547
rect 14968 4521 14998 4547
rect 15052 4521 15082 4547
rect 15240 4521 15270 4547
rect 15324 4521 15354 4547
rect 15408 4521 15438 4547
rect 15492 4521 15522 4547
rect 15582 4521 15612 4547
rect 15681 4521 15711 4547
rect 16553 4613 16583 4769
rect 16649 4723 16679 4895
rect 16625 4707 16679 4723
rect 16625 4673 16635 4707
rect 16669 4673 16679 4707
rect 16625 4657 16679 4673
rect 16649 4613 16679 4657
rect 16721 4723 16751 4895
rect 16817 4851 16847 4895
rect 16906 4851 16936 4895
rect 16990 4880 17020 4895
rect 16793 4835 16847 4851
rect 16793 4801 16803 4835
rect 16837 4801 16847 4835
rect 16793 4785 16847 4801
rect 16893 4835 16947 4851
rect 16893 4801 16903 4835
rect 16937 4801 16947 4835
rect 16893 4785 16947 4801
rect 16989 4850 17020 4880
rect 17074 4880 17104 4895
rect 17262 4880 17292 4895
rect 17074 4850 17292 4880
rect 16721 4707 16775 4723
rect 16721 4673 16731 4707
rect 16765 4673 16775 4707
rect 16721 4657 16775 4673
rect 16721 4613 16751 4657
rect 16817 4613 16847 4785
rect 16906 4613 16936 4785
rect 16989 4739 17019 4850
rect 17074 4835 17115 4850
rect 17085 4739 17115 4835
rect 17346 4820 17376 4895
rect 17430 4821 17460 4895
rect 17322 4804 17376 4820
rect 17322 4770 17332 4804
rect 17366 4770 17376 4804
rect 17322 4754 17376 4770
rect 17418 4805 17472 4821
rect 17418 4771 17428 4805
rect 17462 4771 17472 4805
rect 17418 4755 17472 4771
rect 16978 4723 17032 4739
rect 16978 4689 16988 4723
rect 17022 4689 17032 4723
rect 16978 4673 17032 4689
rect 17085 4723 17149 4739
rect 17085 4689 17105 4723
rect 17139 4689 17149 4723
rect 16990 4613 17020 4673
rect 17085 4658 17149 4689
rect 17074 4628 17292 4658
rect 17074 4613 17104 4628
rect 17262 4613 17292 4628
rect 17346 4613 17376 4754
rect 17430 4613 17460 4755
rect 17514 4716 17544 4895
rect 17604 4827 17634 4895
rect 18427 4912 18457 4938
rect 18523 4912 18553 4938
rect 18595 4912 18625 4938
rect 18809 4912 18839 4938
rect 18912 4912 18942 4938
rect 19021 4873 19051 4899
rect 17703 4827 17733 4849
rect 17586 4811 17640 4827
rect 17586 4777 17596 4811
rect 17630 4777 17640 4811
rect 17586 4761 17640 4777
rect 17682 4811 17736 4827
rect 17682 4777 17692 4811
rect 17726 4777 17736 4811
rect 17682 4761 17736 4777
rect 17508 4700 17562 4716
rect 17508 4666 17518 4700
rect 17552 4666 17562 4700
rect 17508 4650 17562 4666
rect 17514 4613 17544 4650
rect 17604 4613 17634 4761
rect 17703 4729 17733 4761
rect 16454 4503 16484 4529
rect 16553 4503 16583 4529
rect 16649 4503 16679 4529
rect 16721 4503 16751 4529
rect 16817 4503 16847 4529
rect 16906 4503 16936 4529
rect 16990 4503 17020 4529
rect 17074 4503 17104 4529
rect 17262 4503 17292 4529
rect 17346 4503 17376 4529
rect 17430 4503 17460 4529
rect 17514 4503 17544 4529
rect 17604 4503 17634 4529
rect 17703 4503 17733 4529
rect 6208 3293 6238 3319
rect 6208 3141 6238 3163
rect 6208 3125 6294 3141
rect 6208 3091 6244 3125
rect 6278 3091 6294 3125
rect 6208 3075 6294 3091
rect 6208 3043 6238 3075
rect 6208 2817 6238 2843
rect 1920 2241 1950 2267
rect 2019 2241 2049 2267
rect 2115 2241 2145 2267
rect 2187 2241 2217 2267
rect 2283 2241 2313 2267
rect 2372 2241 2402 2267
rect 2456 2241 2486 2267
rect 2540 2241 2570 2267
rect 2728 2241 2758 2267
rect 2812 2241 2842 2267
rect 2896 2241 2926 2267
rect 2980 2241 3010 2267
rect 3070 2241 3100 2267
rect 3169 2241 3199 2267
rect 1920 2089 1950 2111
rect 2019 2097 2049 2157
rect 1920 2073 1974 2089
rect 1920 2039 1930 2073
rect 1964 2039 1974 2073
rect 1920 2023 1974 2039
rect 2019 2081 2073 2097
rect 2019 2047 2029 2081
rect 2063 2047 2073 2081
rect 2019 2031 2073 2047
rect 1920 1991 1950 2023
rect 2019 1875 2049 2031
rect 2115 1985 2145 2157
rect 2091 1969 2145 1985
rect 2091 1935 2101 1969
rect 2135 1935 2145 1969
rect 2091 1919 2145 1935
rect 2115 1875 2145 1919
rect 2187 1985 2217 2157
rect 2283 2113 2313 2157
rect 2372 2113 2402 2157
rect 2456 2142 2486 2157
rect 2259 2097 2313 2113
rect 2259 2063 2269 2097
rect 2303 2063 2313 2097
rect 2259 2047 2313 2063
rect 2359 2097 2413 2113
rect 2359 2063 2369 2097
rect 2403 2063 2413 2097
rect 2359 2047 2413 2063
rect 2455 2112 2486 2142
rect 2540 2142 2570 2157
rect 2728 2142 2758 2157
rect 2540 2112 2758 2142
rect 2187 1969 2241 1985
rect 2187 1935 2197 1969
rect 2231 1935 2241 1969
rect 2187 1919 2241 1935
rect 2187 1875 2217 1919
rect 2283 1875 2313 2047
rect 2372 1875 2402 2047
rect 2455 2001 2485 2112
rect 2540 2097 2581 2112
rect 2551 2001 2581 2097
rect 2812 2082 2842 2157
rect 2896 2083 2926 2157
rect 2788 2066 2842 2082
rect 2788 2032 2798 2066
rect 2832 2032 2842 2066
rect 2788 2016 2842 2032
rect 2884 2067 2938 2083
rect 2884 2033 2894 2067
rect 2928 2033 2938 2067
rect 2884 2017 2938 2033
rect 2444 1985 2498 2001
rect 2444 1951 2454 1985
rect 2488 1951 2498 1985
rect 2444 1935 2498 1951
rect 2551 1985 2615 2001
rect 2551 1951 2571 1985
rect 2605 1951 2615 1985
rect 2456 1875 2486 1935
rect 2551 1920 2615 1951
rect 2540 1890 2758 1920
rect 2540 1875 2570 1890
rect 2728 1875 2758 1890
rect 2812 1875 2842 2016
rect 2896 1875 2926 2017
rect 2980 1978 3010 2157
rect 3070 2089 3100 2157
rect 3990 2237 4020 2263
rect 4089 2237 4119 2263
rect 4185 2237 4215 2263
rect 4257 2237 4287 2263
rect 4353 2237 4383 2263
rect 4442 2237 4472 2263
rect 4526 2237 4556 2263
rect 4610 2237 4640 2263
rect 4798 2237 4828 2263
rect 4882 2237 4912 2263
rect 4966 2237 4996 2263
rect 5050 2237 5080 2263
rect 5140 2237 5170 2263
rect 5239 2237 5269 2263
rect 5942 2237 5972 2263
rect 6041 2237 6071 2263
rect 6137 2237 6167 2263
rect 6209 2237 6239 2263
rect 6305 2237 6335 2263
rect 6394 2237 6424 2263
rect 6478 2237 6508 2263
rect 6562 2237 6592 2263
rect 6750 2237 6780 2263
rect 6834 2237 6864 2263
rect 6918 2237 6948 2263
rect 7002 2237 7032 2263
rect 7092 2237 7122 2263
rect 7191 2237 7221 2263
rect 7944 2243 7974 2269
rect 8043 2243 8073 2269
rect 8139 2243 8169 2269
rect 8211 2243 8241 2269
rect 8307 2243 8337 2269
rect 8396 2243 8426 2269
rect 8480 2243 8510 2269
rect 8564 2243 8594 2269
rect 8752 2243 8782 2269
rect 8836 2243 8866 2269
rect 8920 2243 8950 2269
rect 9004 2243 9034 2269
rect 9094 2243 9124 2269
rect 9193 2243 9223 2269
rect 9896 2243 9926 2269
rect 9995 2243 10025 2269
rect 10091 2243 10121 2269
rect 10163 2243 10193 2269
rect 10259 2243 10289 2269
rect 10348 2243 10378 2269
rect 10432 2243 10462 2269
rect 10516 2243 10546 2269
rect 10704 2243 10734 2269
rect 10788 2243 10818 2269
rect 10872 2243 10902 2269
rect 10956 2243 10986 2269
rect 11046 2243 11076 2269
rect 11145 2243 11175 2269
rect 11888 2243 11918 2269
rect 11987 2243 12017 2269
rect 12083 2243 12113 2269
rect 12155 2243 12185 2269
rect 12251 2243 12281 2269
rect 12340 2243 12370 2269
rect 12424 2243 12454 2269
rect 12508 2243 12538 2269
rect 12696 2243 12726 2269
rect 12780 2243 12810 2269
rect 12864 2243 12894 2269
rect 12948 2243 12978 2269
rect 13038 2243 13068 2269
rect 13137 2243 13167 2269
rect 13840 2243 13870 2269
rect 13939 2243 13969 2269
rect 14035 2243 14065 2269
rect 14107 2243 14137 2269
rect 14203 2243 14233 2269
rect 14292 2243 14322 2269
rect 14376 2243 14406 2269
rect 14460 2243 14490 2269
rect 14648 2243 14678 2269
rect 14732 2243 14762 2269
rect 14816 2243 14846 2269
rect 14900 2243 14930 2269
rect 14990 2243 15020 2269
rect 15089 2243 15119 2269
rect 15904 2243 15934 2269
rect 16003 2243 16033 2269
rect 16099 2243 16129 2269
rect 16171 2243 16201 2269
rect 16267 2243 16297 2269
rect 16356 2243 16386 2269
rect 16440 2243 16470 2269
rect 16524 2243 16554 2269
rect 16712 2243 16742 2269
rect 16796 2243 16826 2269
rect 16880 2243 16910 2269
rect 16964 2243 16994 2269
rect 17054 2243 17084 2269
rect 17153 2243 17183 2269
rect 3169 2089 3199 2111
rect 3052 2073 3106 2089
rect 3052 2039 3062 2073
rect 3096 2039 3106 2073
rect 3052 2023 3106 2039
rect 3148 2073 3202 2089
rect 3148 2039 3158 2073
rect 3192 2039 3202 2073
rect 3148 2023 3202 2039
rect 3990 2085 4020 2107
rect 4089 2093 4119 2153
rect 3990 2069 4044 2085
rect 3990 2035 4000 2069
rect 4034 2035 4044 2069
rect 2974 1962 3028 1978
rect 2974 1928 2984 1962
rect 3018 1928 3028 1962
rect 2974 1912 3028 1928
rect 2980 1875 3010 1912
rect 3070 1875 3100 2023
rect 3169 1991 3199 2023
rect 3990 2019 4044 2035
rect 4089 2077 4143 2093
rect 4089 2043 4099 2077
rect 4133 2043 4143 2077
rect 4089 2027 4143 2043
rect 3990 1987 4020 2019
rect 1920 1765 1950 1791
rect 2019 1765 2049 1791
rect 2115 1765 2145 1791
rect 2187 1765 2217 1791
rect 2283 1765 2313 1791
rect 2372 1765 2402 1791
rect 2456 1765 2486 1791
rect 2540 1765 2570 1791
rect 2728 1765 2758 1791
rect 2812 1765 2842 1791
rect 2896 1765 2926 1791
rect 2980 1765 3010 1791
rect 3070 1765 3100 1791
rect 3169 1765 3199 1791
rect 4089 1871 4119 2027
rect 4185 1981 4215 2153
rect 4161 1965 4215 1981
rect 4161 1931 4171 1965
rect 4205 1931 4215 1965
rect 4161 1915 4215 1931
rect 4185 1871 4215 1915
rect 4257 1981 4287 2153
rect 4353 2109 4383 2153
rect 4442 2109 4472 2153
rect 4526 2138 4556 2153
rect 4329 2093 4383 2109
rect 4329 2059 4339 2093
rect 4373 2059 4383 2093
rect 4329 2043 4383 2059
rect 4429 2093 4483 2109
rect 4429 2059 4439 2093
rect 4473 2059 4483 2093
rect 4429 2043 4483 2059
rect 4525 2108 4556 2138
rect 4610 2138 4640 2153
rect 4798 2138 4828 2153
rect 4610 2108 4828 2138
rect 4257 1965 4311 1981
rect 4257 1931 4267 1965
rect 4301 1931 4311 1965
rect 4257 1915 4311 1931
rect 4257 1871 4287 1915
rect 4353 1871 4383 2043
rect 4442 1871 4472 2043
rect 4525 1997 4555 2108
rect 4610 2093 4651 2108
rect 4621 1997 4651 2093
rect 4882 2078 4912 2153
rect 4966 2079 4996 2153
rect 4858 2062 4912 2078
rect 4858 2028 4868 2062
rect 4902 2028 4912 2062
rect 4858 2012 4912 2028
rect 4954 2063 5008 2079
rect 4954 2029 4964 2063
rect 4998 2029 5008 2063
rect 4954 2013 5008 2029
rect 4514 1981 4568 1997
rect 4514 1947 4524 1981
rect 4558 1947 4568 1981
rect 4514 1931 4568 1947
rect 4621 1981 4685 1997
rect 4621 1947 4641 1981
rect 4675 1947 4685 1981
rect 4526 1871 4556 1931
rect 4621 1916 4685 1947
rect 4610 1886 4828 1916
rect 4610 1871 4640 1886
rect 4798 1871 4828 1886
rect 4882 1871 4912 2012
rect 4966 1871 4996 2013
rect 5050 1974 5080 2153
rect 5140 2085 5170 2153
rect 5239 2085 5269 2107
rect 5942 2085 5972 2107
rect 6041 2093 6071 2153
rect 5122 2069 5176 2085
rect 5122 2035 5132 2069
rect 5166 2035 5176 2069
rect 5122 2019 5176 2035
rect 5218 2069 5272 2085
rect 5218 2035 5228 2069
rect 5262 2035 5272 2069
rect 5218 2019 5272 2035
rect 5942 2069 5996 2085
rect 5942 2035 5952 2069
rect 5986 2035 5996 2069
rect 5942 2019 5996 2035
rect 6041 2077 6095 2093
rect 6041 2043 6051 2077
rect 6085 2043 6095 2077
rect 6041 2027 6095 2043
rect 5044 1958 5098 1974
rect 5044 1924 5054 1958
rect 5088 1924 5098 1958
rect 5044 1908 5098 1924
rect 5050 1871 5080 1908
rect 5140 1871 5170 2019
rect 5239 1987 5269 2019
rect 5942 1987 5972 2019
rect 6041 1871 6071 2027
rect 6137 1981 6167 2153
rect 6113 1965 6167 1981
rect 6113 1931 6123 1965
rect 6157 1931 6167 1965
rect 6113 1915 6167 1931
rect 6137 1871 6167 1915
rect 6209 1981 6239 2153
rect 6305 2109 6335 2153
rect 6394 2109 6424 2153
rect 6478 2138 6508 2153
rect 6281 2093 6335 2109
rect 6281 2059 6291 2093
rect 6325 2059 6335 2093
rect 6281 2043 6335 2059
rect 6381 2093 6435 2109
rect 6381 2059 6391 2093
rect 6425 2059 6435 2093
rect 6381 2043 6435 2059
rect 6477 2108 6508 2138
rect 6562 2138 6592 2153
rect 6750 2138 6780 2153
rect 6562 2108 6780 2138
rect 6209 1965 6263 1981
rect 6209 1931 6219 1965
rect 6253 1931 6263 1965
rect 6209 1915 6263 1931
rect 6209 1871 6239 1915
rect 6305 1871 6335 2043
rect 6394 1871 6424 2043
rect 6477 1997 6507 2108
rect 6562 2093 6603 2108
rect 6573 1997 6603 2093
rect 6834 2078 6864 2153
rect 6918 2079 6948 2153
rect 6810 2062 6864 2078
rect 6810 2028 6820 2062
rect 6854 2028 6864 2062
rect 6810 2012 6864 2028
rect 6906 2063 6960 2079
rect 6906 2029 6916 2063
rect 6950 2029 6960 2063
rect 6906 2013 6960 2029
rect 6466 1981 6520 1997
rect 6466 1947 6476 1981
rect 6510 1947 6520 1981
rect 6466 1931 6520 1947
rect 6573 1981 6637 1997
rect 6573 1947 6593 1981
rect 6627 1947 6637 1981
rect 6478 1871 6508 1931
rect 6573 1916 6637 1947
rect 6562 1886 6780 1916
rect 6562 1871 6592 1886
rect 6750 1871 6780 1886
rect 6834 1871 6864 2012
rect 6918 1871 6948 2013
rect 7002 1974 7032 2153
rect 7092 2085 7122 2153
rect 7191 2085 7221 2107
rect 7944 2091 7974 2113
rect 8043 2099 8073 2159
rect 7074 2069 7128 2085
rect 7074 2035 7084 2069
rect 7118 2035 7128 2069
rect 7074 2019 7128 2035
rect 7170 2069 7224 2085
rect 7170 2035 7180 2069
rect 7214 2035 7224 2069
rect 7170 2019 7224 2035
rect 7944 2075 7998 2091
rect 7944 2041 7954 2075
rect 7988 2041 7998 2075
rect 7944 2025 7998 2041
rect 8043 2083 8097 2099
rect 8043 2049 8053 2083
rect 8087 2049 8097 2083
rect 8043 2033 8097 2049
rect 6996 1958 7050 1974
rect 6996 1924 7006 1958
rect 7040 1924 7050 1958
rect 6996 1908 7050 1924
rect 7002 1871 7032 1908
rect 7092 1871 7122 2019
rect 7191 1987 7221 2019
rect 7944 1993 7974 2025
rect 8043 1877 8073 2033
rect 8139 1987 8169 2159
rect 8115 1971 8169 1987
rect 8115 1937 8125 1971
rect 8159 1937 8169 1971
rect 8115 1921 8169 1937
rect 8139 1877 8169 1921
rect 8211 1987 8241 2159
rect 8307 2115 8337 2159
rect 8396 2115 8426 2159
rect 8480 2144 8510 2159
rect 8283 2099 8337 2115
rect 8283 2065 8293 2099
rect 8327 2065 8337 2099
rect 8283 2049 8337 2065
rect 8383 2099 8437 2115
rect 8383 2065 8393 2099
rect 8427 2065 8437 2099
rect 8383 2049 8437 2065
rect 8479 2114 8510 2144
rect 8564 2144 8594 2159
rect 8752 2144 8782 2159
rect 8564 2114 8782 2144
rect 8211 1971 8265 1987
rect 8211 1937 8221 1971
rect 8255 1937 8265 1971
rect 8211 1921 8265 1937
rect 8211 1877 8241 1921
rect 8307 1877 8337 2049
rect 8396 1877 8426 2049
rect 8479 2003 8509 2114
rect 8564 2099 8605 2114
rect 8575 2003 8605 2099
rect 8836 2084 8866 2159
rect 8920 2085 8950 2159
rect 8812 2068 8866 2084
rect 8812 2034 8822 2068
rect 8856 2034 8866 2068
rect 8812 2018 8866 2034
rect 8908 2069 8962 2085
rect 8908 2035 8918 2069
rect 8952 2035 8962 2069
rect 8908 2019 8962 2035
rect 8468 1987 8522 2003
rect 8468 1953 8478 1987
rect 8512 1953 8522 1987
rect 8468 1937 8522 1953
rect 8575 1987 8639 2003
rect 8575 1953 8595 1987
rect 8629 1953 8639 1987
rect 8480 1877 8510 1937
rect 8575 1922 8639 1953
rect 8564 1892 8782 1922
rect 8564 1877 8594 1892
rect 8752 1877 8782 1892
rect 8836 1877 8866 2018
rect 8920 1877 8950 2019
rect 9004 1980 9034 2159
rect 9094 2091 9124 2159
rect 9193 2091 9223 2113
rect 9896 2091 9926 2113
rect 9995 2099 10025 2159
rect 9076 2075 9130 2091
rect 9076 2041 9086 2075
rect 9120 2041 9130 2075
rect 9076 2025 9130 2041
rect 9172 2075 9226 2091
rect 9172 2041 9182 2075
rect 9216 2041 9226 2075
rect 9172 2025 9226 2041
rect 9896 2075 9950 2091
rect 9896 2041 9906 2075
rect 9940 2041 9950 2075
rect 9896 2025 9950 2041
rect 9995 2083 10049 2099
rect 9995 2049 10005 2083
rect 10039 2049 10049 2083
rect 9995 2033 10049 2049
rect 8998 1964 9052 1980
rect 8998 1930 9008 1964
rect 9042 1930 9052 1964
rect 8998 1914 9052 1930
rect 9004 1877 9034 1914
rect 9094 1877 9124 2025
rect 9193 1993 9223 2025
rect 9896 1993 9926 2025
rect 9995 1877 10025 2033
rect 10091 1987 10121 2159
rect 10067 1971 10121 1987
rect 10067 1937 10077 1971
rect 10111 1937 10121 1971
rect 10067 1921 10121 1937
rect 10091 1877 10121 1921
rect 10163 1987 10193 2159
rect 10259 2115 10289 2159
rect 10348 2115 10378 2159
rect 10432 2144 10462 2159
rect 10235 2099 10289 2115
rect 10235 2065 10245 2099
rect 10279 2065 10289 2099
rect 10235 2049 10289 2065
rect 10335 2099 10389 2115
rect 10335 2065 10345 2099
rect 10379 2065 10389 2099
rect 10335 2049 10389 2065
rect 10431 2114 10462 2144
rect 10516 2144 10546 2159
rect 10704 2144 10734 2159
rect 10516 2114 10734 2144
rect 10163 1971 10217 1987
rect 10163 1937 10173 1971
rect 10207 1937 10217 1971
rect 10163 1921 10217 1937
rect 10163 1877 10193 1921
rect 10259 1877 10289 2049
rect 10348 1877 10378 2049
rect 10431 2003 10461 2114
rect 10516 2099 10557 2114
rect 10527 2003 10557 2099
rect 10788 2084 10818 2159
rect 10872 2085 10902 2159
rect 10764 2068 10818 2084
rect 10764 2034 10774 2068
rect 10808 2034 10818 2068
rect 10764 2018 10818 2034
rect 10860 2069 10914 2085
rect 10860 2035 10870 2069
rect 10904 2035 10914 2069
rect 10860 2019 10914 2035
rect 10420 1987 10474 2003
rect 10420 1953 10430 1987
rect 10464 1953 10474 1987
rect 10420 1937 10474 1953
rect 10527 1987 10591 2003
rect 10527 1953 10547 1987
rect 10581 1953 10591 1987
rect 10432 1877 10462 1937
rect 10527 1922 10591 1953
rect 10516 1892 10734 1922
rect 10516 1877 10546 1892
rect 10704 1877 10734 1892
rect 10788 1877 10818 2018
rect 10872 1877 10902 2019
rect 10956 1980 10986 2159
rect 11046 2091 11076 2159
rect 11145 2091 11175 2113
rect 11888 2091 11918 2113
rect 11987 2099 12017 2159
rect 11028 2075 11082 2091
rect 11028 2041 11038 2075
rect 11072 2041 11082 2075
rect 11028 2025 11082 2041
rect 11124 2075 11178 2091
rect 11124 2041 11134 2075
rect 11168 2041 11178 2075
rect 11124 2025 11178 2041
rect 11888 2075 11942 2091
rect 11888 2041 11898 2075
rect 11932 2041 11942 2075
rect 11888 2025 11942 2041
rect 11987 2083 12041 2099
rect 11987 2049 11997 2083
rect 12031 2049 12041 2083
rect 11987 2033 12041 2049
rect 10950 1964 11004 1980
rect 10950 1930 10960 1964
rect 10994 1930 11004 1964
rect 10950 1914 11004 1930
rect 10956 1877 10986 1914
rect 11046 1877 11076 2025
rect 11145 1993 11175 2025
rect 11888 1993 11918 2025
rect 11987 1877 12017 2033
rect 12083 1987 12113 2159
rect 12059 1971 12113 1987
rect 12059 1937 12069 1971
rect 12103 1937 12113 1971
rect 12059 1921 12113 1937
rect 12083 1877 12113 1921
rect 12155 1987 12185 2159
rect 12251 2115 12281 2159
rect 12340 2115 12370 2159
rect 12424 2144 12454 2159
rect 12227 2099 12281 2115
rect 12227 2065 12237 2099
rect 12271 2065 12281 2099
rect 12227 2049 12281 2065
rect 12327 2099 12381 2115
rect 12327 2065 12337 2099
rect 12371 2065 12381 2099
rect 12327 2049 12381 2065
rect 12423 2114 12454 2144
rect 12508 2144 12538 2159
rect 12696 2144 12726 2159
rect 12508 2114 12726 2144
rect 12155 1971 12209 1987
rect 12155 1937 12165 1971
rect 12199 1937 12209 1971
rect 12155 1921 12209 1937
rect 12155 1877 12185 1921
rect 12251 1877 12281 2049
rect 12340 1877 12370 2049
rect 12423 2003 12453 2114
rect 12508 2099 12549 2114
rect 12519 2003 12549 2099
rect 12780 2084 12810 2159
rect 12864 2085 12894 2159
rect 12756 2068 12810 2084
rect 12756 2034 12766 2068
rect 12800 2034 12810 2068
rect 12756 2018 12810 2034
rect 12852 2069 12906 2085
rect 12852 2035 12862 2069
rect 12896 2035 12906 2069
rect 12852 2019 12906 2035
rect 12412 1987 12466 2003
rect 12412 1953 12422 1987
rect 12456 1953 12466 1987
rect 12412 1937 12466 1953
rect 12519 1987 12583 2003
rect 12519 1953 12539 1987
rect 12573 1953 12583 1987
rect 12424 1877 12454 1937
rect 12519 1922 12583 1953
rect 12508 1892 12726 1922
rect 12508 1877 12538 1892
rect 12696 1877 12726 1892
rect 12780 1877 12810 2018
rect 12864 1877 12894 2019
rect 12948 1980 12978 2159
rect 13038 2091 13068 2159
rect 13137 2091 13167 2113
rect 13840 2091 13870 2113
rect 13939 2099 13969 2159
rect 13020 2075 13074 2091
rect 13020 2041 13030 2075
rect 13064 2041 13074 2075
rect 13020 2025 13074 2041
rect 13116 2075 13170 2091
rect 13116 2041 13126 2075
rect 13160 2041 13170 2075
rect 13116 2025 13170 2041
rect 13840 2075 13894 2091
rect 13840 2041 13850 2075
rect 13884 2041 13894 2075
rect 13840 2025 13894 2041
rect 13939 2083 13993 2099
rect 13939 2049 13949 2083
rect 13983 2049 13993 2083
rect 13939 2033 13993 2049
rect 12942 1964 12996 1980
rect 12942 1930 12952 1964
rect 12986 1930 12996 1964
rect 12942 1914 12996 1930
rect 12948 1877 12978 1914
rect 13038 1877 13068 2025
rect 13137 1993 13167 2025
rect 13840 1993 13870 2025
rect 13939 1877 13969 2033
rect 14035 1987 14065 2159
rect 14011 1971 14065 1987
rect 14011 1937 14021 1971
rect 14055 1937 14065 1971
rect 14011 1921 14065 1937
rect 14035 1877 14065 1921
rect 14107 1987 14137 2159
rect 14203 2115 14233 2159
rect 14292 2115 14322 2159
rect 14376 2144 14406 2159
rect 14179 2099 14233 2115
rect 14179 2065 14189 2099
rect 14223 2065 14233 2099
rect 14179 2049 14233 2065
rect 14279 2099 14333 2115
rect 14279 2065 14289 2099
rect 14323 2065 14333 2099
rect 14279 2049 14333 2065
rect 14375 2114 14406 2144
rect 14460 2144 14490 2159
rect 14648 2144 14678 2159
rect 14460 2114 14678 2144
rect 14107 1971 14161 1987
rect 14107 1937 14117 1971
rect 14151 1937 14161 1971
rect 14107 1921 14161 1937
rect 14107 1877 14137 1921
rect 14203 1877 14233 2049
rect 14292 1877 14322 2049
rect 14375 2003 14405 2114
rect 14460 2099 14501 2114
rect 14471 2003 14501 2099
rect 14732 2084 14762 2159
rect 14816 2085 14846 2159
rect 14708 2068 14762 2084
rect 14708 2034 14718 2068
rect 14752 2034 14762 2068
rect 14708 2018 14762 2034
rect 14804 2069 14858 2085
rect 14804 2035 14814 2069
rect 14848 2035 14858 2069
rect 14804 2019 14858 2035
rect 14364 1987 14418 2003
rect 14364 1953 14374 1987
rect 14408 1953 14418 1987
rect 14364 1937 14418 1953
rect 14471 1987 14535 2003
rect 14471 1953 14491 1987
rect 14525 1953 14535 1987
rect 14376 1877 14406 1937
rect 14471 1922 14535 1953
rect 14460 1892 14678 1922
rect 14460 1877 14490 1892
rect 14648 1877 14678 1892
rect 14732 1877 14762 2018
rect 14816 1877 14846 2019
rect 14900 1980 14930 2159
rect 14990 2091 15020 2159
rect 15089 2091 15119 2113
rect 15904 2091 15934 2113
rect 16003 2099 16033 2159
rect 14972 2075 15026 2091
rect 14972 2041 14982 2075
rect 15016 2041 15026 2075
rect 14972 2025 15026 2041
rect 15068 2075 15122 2091
rect 15068 2041 15078 2075
rect 15112 2041 15122 2075
rect 15068 2025 15122 2041
rect 15904 2075 15958 2091
rect 15904 2041 15914 2075
rect 15948 2041 15958 2075
rect 15904 2025 15958 2041
rect 16003 2083 16057 2099
rect 16003 2049 16013 2083
rect 16047 2049 16057 2083
rect 16003 2033 16057 2049
rect 14894 1964 14948 1980
rect 14894 1930 14904 1964
rect 14938 1930 14948 1964
rect 14894 1914 14948 1930
rect 14900 1877 14930 1914
rect 14990 1877 15020 2025
rect 15089 1993 15119 2025
rect 15904 1993 15934 2025
rect 16003 1877 16033 2033
rect 16099 1987 16129 2159
rect 16075 1971 16129 1987
rect 16075 1937 16085 1971
rect 16119 1937 16129 1971
rect 16075 1921 16129 1937
rect 16099 1877 16129 1921
rect 16171 1987 16201 2159
rect 16267 2115 16297 2159
rect 16356 2115 16386 2159
rect 16440 2144 16470 2159
rect 16243 2099 16297 2115
rect 16243 2065 16253 2099
rect 16287 2065 16297 2099
rect 16243 2049 16297 2065
rect 16343 2099 16397 2115
rect 16343 2065 16353 2099
rect 16387 2065 16397 2099
rect 16343 2049 16397 2065
rect 16439 2114 16470 2144
rect 16524 2144 16554 2159
rect 16712 2144 16742 2159
rect 16524 2114 16742 2144
rect 16171 1971 16225 1987
rect 16171 1937 16181 1971
rect 16215 1937 16225 1971
rect 16171 1921 16225 1937
rect 16171 1877 16201 1921
rect 16267 1877 16297 2049
rect 16356 1877 16386 2049
rect 16439 2003 16469 2114
rect 16524 2099 16565 2114
rect 16535 2003 16565 2099
rect 16796 2084 16826 2159
rect 16880 2085 16910 2159
rect 16772 2068 16826 2084
rect 16772 2034 16782 2068
rect 16816 2034 16826 2068
rect 16772 2018 16826 2034
rect 16868 2069 16922 2085
rect 16868 2035 16878 2069
rect 16912 2035 16922 2069
rect 16868 2019 16922 2035
rect 16428 1987 16482 2003
rect 16428 1953 16438 1987
rect 16472 1953 16482 1987
rect 16428 1937 16482 1953
rect 16535 1987 16599 2003
rect 16535 1953 16555 1987
rect 16589 1953 16599 1987
rect 16440 1877 16470 1937
rect 16535 1922 16599 1953
rect 16524 1892 16742 1922
rect 16524 1877 16554 1892
rect 16712 1877 16742 1892
rect 16796 1877 16826 2018
rect 16880 1877 16910 2019
rect 16964 1980 16994 2159
rect 17054 2091 17084 2159
rect 17153 2091 17183 2113
rect 17036 2075 17090 2091
rect 17036 2041 17046 2075
rect 17080 2041 17090 2075
rect 17036 2025 17090 2041
rect 17132 2075 17186 2091
rect 17132 2041 17142 2075
rect 17176 2041 17186 2075
rect 17132 2025 17186 2041
rect 16958 1964 17012 1980
rect 16958 1930 16968 1964
rect 17002 1930 17012 1964
rect 16958 1914 17012 1930
rect 16964 1877 16994 1914
rect 17054 1877 17084 2025
rect 17153 1993 17183 2025
rect 3990 1761 4020 1787
rect 4089 1761 4119 1787
rect 4185 1761 4215 1787
rect 4257 1761 4287 1787
rect 4353 1761 4383 1787
rect 4442 1761 4472 1787
rect 4526 1761 4556 1787
rect 4610 1761 4640 1787
rect 4798 1761 4828 1787
rect 4882 1761 4912 1787
rect 4966 1761 4996 1787
rect 5050 1761 5080 1787
rect 5140 1761 5170 1787
rect 5239 1761 5269 1787
rect 5942 1761 5972 1787
rect 6041 1761 6071 1787
rect 6137 1761 6167 1787
rect 6209 1761 6239 1787
rect 6305 1761 6335 1787
rect 6394 1761 6424 1787
rect 6478 1761 6508 1787
rect 6562 1761 6592 1787
rect 6750 1761 6780 1787
rect 6834 1761 6864 1787
rect 6918 1761 6948 1787
rect 7002 1761 7032 1787
rect 7092 1761 7122 1787
rect 7191 1761 7221 1787
rect 7944 1767 7974 1793
rect 8043 1767 8073 1793
rect 8139 1767 8169 1793
rect 8211 1767 8241 1793
rect 8307 1767 8337 1793
rect 8396 1767 8426 1793
rect 8480 1767 8510 1793
rect 8564 1767 8594 1793
rect 8752 1767 8782 1793
rect 8836 1767 8866 1793
rect 8920 1767 8950 1793
rect 9004 1767 9034 1793
rect 9094 1767 9124 1793
rect 9193 1767 9223 1793
rect 9896 1767 9926 1793
rect 9995 1767 10025 1793
rect 10091 1767 10121 1793
rect 10163 1767 10193 1793
rect 10259 1767 10289 1793
rect 10348 1767 10378 1793
rect 10432 1767 10462 1793
rect 10516 1767 10546 1793
rect 10704 1767 10734 1793
rect 10788 1767 10818 1793
rect 10872 1767 10902 1793
rect 10956 1767 10986 1793
rect 11046 1767 11076 1793
rect 11145 1767 11175 1793
rect 11888 1767 11918 1793
rect 11987 1767 12017 1793
rect 12083 1767 12113 1793
rect 12155 1767 12185 1793
rect 12251 1767 12281 1793
rect 12340 1767 12370 1793
rect 12424 1767 12454 1793
rect 12508 1767 12538 1793
rect 12696 1767 12726 1793
rect 12780 1767 12810 1793
rect 12864 1767 12894 1793
rect 12948 1767 12978 1793
rect 13038 1767 13068 1793
rect 13137 1767 13167 1793
rect 13840 1767 13870 1793
rect 13939 1767 13969 1793
rect 14035 1767 14065 1793
rect 14107 1767 14137 1793
rect 14203 1767 14233 1793
rect 14292 1767 14322 1793
rect 14376 1767 14406 1793
rect 14460 1767 14490 1793
rect 14648 1767 14678 1793
rect 14732 1767 14762 1793
rect 14816 1767 14846 1793
rect 14900 1767 14930 1793
rect 14990 1767 15020 1793
rect 15089 1767 15119 1793
rect 15904 1767 15934 1793
rect 16003 1767 16033 1793
rect 16099 1767 16129 1793
rect 16171 1767 16201 1793
rect 16267 1767 16297 1793
rect 16356 1767 16386 1793
rect 16440 1767 16470 1793
rect 16524 1767 16554 1793
rect 16712 1767 16742 1793
rect 16796 1767 16826 1793
rect 16880 1767 16910 1793
rect 16964 1767 16994 1793
rect 17054 1767 17084 1793
rect 17153 1767 17183 1793
<< polycont >>
rect 18891 43003 18925 43037
rect 18891 42836 18925 42870
rect 18891 42668 18925 42702
rect 18891 42501 18925 42535
rect 18891 42332 18925 42366
rect 18891 42164 18925 42198
rect 18891 41990 18925 42024
rect 18875 41228 18909 41262
rect 18875 41144 18909 41178
rect 18875 41060 18909 41094
rect 18875 40976 18909 41010
rect 18875 40892 18909 40926
rect 18875 40808 18909 40842
rect 18875 40724 18909 40758
rect 18875 40640 18909 40674
rect 18875 40556 18909 40590
rect 18875 40472 18909 40506
rect 18875 40388 18909 40422
rect 18883 39464 18917 39498
rect 18883 39380 18917 39414
rect 18883 39296 18917 39330
rect 18883 39212 18917 39246
rect 18883 39128 18917 39162
rect 18883 39044 18917 39078
rect 18883 38960 18917 38994
rect 18897 38203 18931 38237
rect 18897 38119 18931 38153
rect 18897 38035 18931 38069
rect 18897 37767 18931 37801
rect 18909 37061 18943 37095
rect 18909 36977 18943 37011
rect 18909 36893 18943 36927
rect 18909 36801 18943 36835
rect 18917 36097 18951 36131
rect 18941 34815 18975 34849
rect 18941 34554 18975 34588
rect 18941 34370 18975 34404
rect 18825 34296 18859 34330
rect 18825 34160 18859 34194
rect 18891 34058 18925 34092
rect 18999 34101 19033 34135
rect 18891 33922 18925 33956
rect 18987 33858 19021 33892
rect 18825 33748 18859 33782
rect 18903 33639 18937 33673
rect 18999 33659 19033 33693
rect 18873 33496 18907 33530
rect 18926 33334 18960 33368
rect 18941 33232 18975 33266
rect 18941 32533 18975 32567
rect 18941 32272 18975 32306
rect 18941 32088 18975 32122
rect 18825 32014 18859 32048
rect 18825 31878 18859 31912
rect 18891 31776 18925 31810
rect 18999 31819 19033 31853
rect 18891 31640 18925 31674
rect 18987 31576 19021 31610
rect 18825 31466 18859 31500
rect 18903 31357 18937 31391
rect 18999 31377 19033 31411
rect 18873 31214 18907 31248
rect 18926 31052 18960 31086
rect 18941 30950 18975 30984
rect 18945 30287 18979 30321
rect 18945 30026 18979 30060
rect 18945 29842 18979 29876
rect 18829 29768 18863 29802
rect 18829 29632 18863 29666
rect 18895 29530 18929 29564
rect 19003 29573 19037 29607
rect 18895 29394 18929 29428
rect 18991 29330 19025 29364
rect 18829 29220 18863 29254
rect 18907 29111 18941 29145
rect 19003 29131 19037 29165
rect 18877 28968 18911 29002
rect 18930 28806 18964 28840
rect 18945 28704 18979 28738
rect 18937 28101 18971 28135
rect 18937 27840 18971 27874
rect 18937 27656 18971 27690
rect 18821 27582 18855 27616
rect 18821 27446 18855 27480
rect 18887 27344 18921 27378
rect 18995 27387 19029 27421
rect 18887 27208 18921 27242
rect 18983 27144 19017 27178
rect 18821 27034 18855 27068
rect 18899 26925 18933 26959
rect 18995 26945 19029 26979
rect 18869 26782 18903 26816
rect 18922 26620 18956 26654
rect 18937 26518 18971 26552
rect 18941 25855 18975 25889
rect 18941 25594 18975 25628
rect 18941 25410 18975 25444
rect 18825 25336 18859 25370
rect 18825 25200 18859 25234
rect 18891 25098 18925 25132
rect 18999 25141 19033 25175
rect 18891 24962 18925 24996
rect 18987 24898 19021 24932
rect 18825 24788 18859 24822
rect 18903 24679 18937 24713
rect 18999 24699 19033 24733
rect 18873 24536 18907 24570
rect 18926 24374 18960 24408
rect 18941 24272 18975 24306
rect 7702 23043 7736 23077
rect 7966 23111 8000 23145
rect 8218 23159 8252 23193
rect 7804 23058 7838 23092
rect 8109 23081 8143 23115
rect 8129 22985 8163 23019
rect 8630 23159 8664 23193
rect 8766 23159 8800 23193
rect 8392 23093 8426 23127
rect 8528 23093 8562 23127
rect 8328 22997 8362 23031
rect 8571 22985 8605 23019
rect 8840 23043 8874 23077
rect 9024 23043 9058 23077
rect 9285 23043 9319 23077
rect 9948 23047 9982 23081
rect 10212 23115 10246 23149
rect 10464 23163 10498 23197
rect 10050 23062 10084 23096
rect 10355 23085 10389 23119
rect 10375 22989 10409 23023
rect 10876 23163 10910 23197
rect 11012 23163 11046 23197
rect 10638 23097 10672 23131
rect 10774 23097 10808 23131
rect 10574 23001 10608 23035
rect 10817 22989 10851 23023
rect 11086 23047 11120 23081
rect 11270 23047 11304 23081
rect 11531 23047 11565 23081
rect 12134 23039 12168 23073
rect 12398 23107 12432 23141
rect 12650 23155 12684 23189
rect 12236 23054 12270 23088
rect 12541 23077 12575 23111
rect 12561 22981 12595 23015
rect 13062 23155 13096 23189
rect 13198 23155 13232 23189
rect 12824 23089 12858 23123
rect 12960 23089 12994 23123
rect 12760 22993 12794 23027
rect 13003 22981 13037 23015
rect 13272 23039 13306 23073
rect 13456 23039 13490 23073
rect 13717 23039 13751 23073
rect 14380 23043 14414 23077
rect 14644 23111 14678 23145
rect 14896 23159 14930 23193
rect 14482 23058 14516 23092
rect 14787 23081 14821 23115
rect 14807 22985 14841 23019
rect 15308 23159 15342 23193
rect 15444 23159 15478 23193
rect 15070 23093 15104 23127
rect 15206 23093 15240 23127
rect 15006 22997 15040 23031
rect 15249 22985 15283 23019
rect 15518 23043 15552 23077
rect 15702 23043 15736 23077
rect 15963 23043 15997 23077
rect 16662 23043 16696 23077
rect 16926 23111 16960 23145
rect 17178 23159 17212 23193
rect 16764 23058 16798 23092
rect 17069 23081 17103 23115
rect 17089 22985 17123 23019
rect 17590 23159 17624 23193
rect 17726 23159 17760 23193
rect 17352 23093 17386 23127
rect 17488 23093 17522 23127
rect 17288 22997 17322 23031
rect 17531 22985 17565 23019
rect 17800 23043 17834 23077
rect 17984 23043 18018 23077
rect 18245 23043 18279 23077
rect 9592 17545 9626 17579
rect 15729 17397 15763 17431
rect 16507 17435 16541 17469
rect 17381 17437 17415 17471
rect 18149 17427 18183 17461
rect 19271 17429 19305 17463
rect 20145 17431 20179 17465
rect 20913 17421 20947 17455
rect 21527 17419 21561 17453
rect 22401 17421 22435 17455
rect 23169 17411 23203 17445
rect 16416 16365 16450 16399
rect 17184 16355 17218 16389
rect 18058 16357 18092 16391
rect 4553 16257 4587 16291
rect 4670 16257 4704 16291
rect 4805 16257 4839 16291
rect 4901 16257 4935 16291
rect 9419 16261 9453 16295
rect 9536 16261 9570 16295
rect 9671 16261 9705 16295
rect 9767 16261 9801 16295
rect 18672 16355 18706 16389
rect 19440 16345 19474 16379
rect 20314 16347 20348 16381
rect 21436 16349 21470 16383
rect 22204 16339 22238 16373
rect 23078 16341 23112 16375
rect 4640 15513 4674 15547
rect 4781 15513 4815 15547
rect 4889 15513 4923 15547
rect 9506 15517 9540 15551
rect 6639 15403 6673 15437
rect 6785 15403 6819 15437
rect 6891 15403 6925 15437
rect 6987 15403 7021 15437
rect 7098 15403 7132 15437
rect 9647 15517 9681 15551
rect 9755 15517 9789 15551
rect 11505 15407 11539 15441
rect 11651 15407 11685 15441
rect 11757 15407 11791 15441
rect 11853 15407 11887 15441
rect 11964 15407 11998 15441
rect 5824 14903 5858 14937
rect 5965 14903 5999 14937
rect 6073 14903 6107 14937
rect 4563 14693 4597 14727
rect 4680 14693 4714 14727
rect 4815 14693 4849 14727
rect 10690 14907 10724 14941
rect 10831 14907 10865 14941
rect 10939 14907 10973 14941
rect 4911 14693 4945 14727
rect 9429 14697 9463 14731
rect 9546 14697 9580 14731
rect 9681 14697 9715 14731
rect 9777 14697 9811 14731
rect 23549 14503 23583 14537
rect 23645 14503 23679 14537
rect 23916 14511 23950 14545
rect 24150 14507 24184 14541
rect 24315 14507 24349 14541
rect 24459 14515 24493 14549
rect 24566 14515 24600 14549
rect 24695 14503 24729 14537
rect 25138 14509 25172 14543
rect 25275 14503 25309 14537
rect 4650 13949 4684 13983
rect 4791 13949 4825 13983
rect 7979 14145 8013 14179
rect 4899 13949 4933 13983
rect 5855 13937 5889 13971
rect 6001 13937 6035 13971
rect 6107 13937 6141 13971
rect 6203 13937 6237 13971
rect 6314 13937 6348 13971
rect 7757 13921 7791 13955
rect 7883 13921 7917 13955
rect 8059 13921 8093 13955
rect 8155 13921 8189 13955
rect 9516 13953 9550 13987
rect 9657 13953 9691 13987
rect 12845 14149 12879 14183
rect 9765 13953 9799 13987
rect 10721 13941 10755 13975
rect 10867 13941 10901 13975
rect 10973 13941 11007 13975
rect 11069 13941 11103 13975
rect 11180 13941 11214 13975
rect 12623 13925 12657 13959
rect 12749 13925 12783 13959
rect 12925 13925 12959 13959
rect 13021 13925 13055 13959
rect 6860 13563 6894 13597
rect 6996 13563 7030 13597
rect 7099 13563 7133 13597
rect 11726 13567 11760 13601
rect 11862 13567 11896 13601
rect 11965 13567 11999 13601
rect 6121 13322 6155 13356
rect 4555 13025 4589 13059
rect 4672 13025 4706 13059
rect 4807 13025 4841 13059
rect 4903 13025 4937 13059
rect 5983 13049 6017 13083
rect 6193 13089 6227 13123
rect 6289 13095 6323 13129
rect 10987 13326 11021 13360
rect 9421 13029 9455 13063
rect 9538 13029 9572 13063
rect 9673 13029 9707 13063
rect 9769 13029 9803 13063
rect 10849 13053 10883 13087
rect 11059 13093 11093 13127
rect 11155 13099 11189 13133
rect 4642 12281 4676 12315
rect 4783 12281 4817 12315
rect 4891 12281 4925 12315
rect 6018 12075 6052 12109
rect 9508 12285 9542 12319
rect 9649 12285 9683 12319
rect 9757 12285 9791 12319
rect 6159 12075 6193 12109
rect 6267 12075 6301 12109
rect 10884 12079 10918 12113
rect 11025 12079 11059 12113
rect 11133 12079 11167 12113
rect 4565 11461 4599 11495
rect 4682 11461 4716 11495
rect 4817 11461 4851 11495
rect 4913 11461 4947 11495
rect 9431 11465 9465 11499
rect 9548 11465 9582 11499
rect 9683 11465 9717 11499
rect 9779 11465 9813 11499
rect 4652 10717 4686 10751
rect 4793 10717 4827 10751
rect 4901 10717 4935 10751
rect 9518 10721 9552 10755
rect 9659 10721 9693 10755
rect 9767 10721 9801 10755
rect 6274 6351 6308 6385
rect 10142 5719 10176 5753
rect 10241 5727 10275 5761
rect 1960 5299 1994 5333
rect 2059 5307 2093 5341
rect 2131 5195 2165 5229
rect 2299 5323 2333 5357
rect 2399 5323 2433 5357
rect 2227 5195 2261 5229
rect 2828 5292 2862 5326
rect 2924 5293 2958 5327
rect 2484 5211 2518 5245
rect 2601 5211 2635 5245
rect 3092 5299 3126 5333
rect 3188 5299 3222 5333
rect 4094 5291 4128 5325
rect 3014 5188 3048 5222
rect 4193 5299 4227 5333
rect 4265 5187 4299 5221
rect 4433 5315 4467 5349
rect 4533 5315 4567 5349
rect 4361 5187 4395 5221
rect 4962 5284 4996 5318
rect 5058 5285 5092 5319
rect 4618 5203 4652 5237
rect 4735 5203 4769 5237
rect 5226 5291 5260 5325
rect 5322 5291 5356 5325
rect 6046 5291 6080 5325
rect 6145 5299 6179 5333
rect 5148 5180 5182 5214
rect 6217 5187 6251 5221
rect 6385 5315 6419 5349
rect 6485 5315 6519 5349
rect 6313 5187 6347 5221
rect 6914 5284 6948 5318
rect 7010 5285 7044 5319
rect 6570 5203 6604 5237
rect 6687 5203 6721 5237
rect 7178 5291 7212 5325
rect 7274 5291 7308 5325
rect 8048 5297 8082 5331
rect 8147 5305 8181 5339
rect 7100 5180 7134 5214
rect 8219 5193 8253 5227
rect 8387 5321 8421 5355
rect 8487 5321 8521 5355
rect 8315 5193 8349 5227
rect 8916 5290 8950 5324
rect 9012 5291 9046 5325
rect 8572 5209 8606 5243
rect 8689 5209 8723 5243
rect 10313 5615 10347 5649
rect 10481 5743 10515 5777
rect 10581 5743 10615 5777
rect 10409 5615 10443 5649
rect 11010 5712 11044 5746
rect 11106 5713 11140 5747
rect 10666 5631 10700 5665
rect 10783 5631 10817 5665
rect 11274 5719 11308 5753
rect 11370 5719 11404 5753
rect 12204 5707 12238 5741
rect 11196 5608 11230 5642
rect 12303 5715 12337 5749
rect 12375 5603 12409 5637
rect 12543 5731 12577 5765
rect 12643 5731 12677 5765
rect 12471 5603 12505 5637
rect 13072 5700 13106 5734
rect 13168 5701 13202 5735
rect 12728 5619 12762 5653
rect 12845 5619 12879 5653
rect 13336 5707 13370 5741
rect 13432 5707 13466 5741
rect 14162 5715 14196 5749
rect 14261 5723 14295 5757
rect 13258 5596 13292 5630
rect 14333 5611 14367 5645
rect 14501 5739 14535 5773
rect 14601 5739 14635 5773
rect 14429 5611 14463 5645
rect 15030 5708 15064 5742
rect 15126 5709 15160 5743
rect 14686 5627 14720 5661
rect 14803 5627 14837 5661
rect 15294 5715 15328 5749
rect 15390 5715 15424 5749
rect 16156 5721 16190 5755
rect 16255 5729 16289 5763
rect 15216 5604 15250 5638
rect 16327 5617 16361 5651
rect 16495 5745 16529 5779
rect 16595 5745 16629 5779
rect 16423 5617 16457 5651
rect 17024 5714 17058 5748
rect 17120 5715 17154 5749
rect 16680 5633 16714 5667
rect 16797 5633 16831 5667
rect 17288 5721 17322 5755
rect 17384 5721 17418 5755
rect 17210 5610 17244 5644
rect 9180 5297 9214 5331
rect 9276 5297 9310 5331
rect 9102 5186 9136 5220
rect 18515 5183 18549 5217
rect 18677 5183 18711 5217
rect 18437 5070 18471 5104
rect 10170 4845 10204 4879
rect 10269 4853 10303 4887
rect 10341 4741 10375 4775
rect 10509 4869 10543 4903
rect 10609 4869 10643 4903
rect 10437 4741 10471 4775
rect 11038 4838 11072 4872
rect 11134 4839 11168 4873
rect 10694 4757 10728 4791
rect 10811 4757 10845 4791
rect 11302 4845 11336 4879
rect 11398 4845 11432 4879
rect 11224 4734 11258 4768
rect 12440 4801 12474 4835
rect 12539 4809 12573 4843
rect 12611 4697 12645 4731
rect 12779 4825 12813 4859
rect 12879 4825 12913 4859
rect 12707 4697 12741 4731
rect 13308 4794 13342 4828
rect 13404 4795 13438 4829
rect 12964 4713 12998 4747
rect 13081 4713 13115 4747
rect 18773 5183 18807 5217
rect 18605 5070 18639 5104
rect 18914 5147 18948 5181
rect 19010 5147 19044 5181
rect 13572 4801 13606 4835
rect 13668 4801 13702 4835
rect 14442 4795 14476 4829
rect 13494 4690 13528 4724
rect 14541 4803 14575 4837
rect 14613 4691 14647 4725
rect 14781 4819 14815 4853
rect 14881 4819 14915 4853
rect 14709 4691 14743 4725
rect 15310 4788 15344 4822
rect 15406 4789 15440 4823
rect 14966 4707 15000 4741
rect 15083 4707 15117 4741
rect 15574 4795 15608 4829
rect 15670 4795 15704 4829
rect 15496 4684 15530 4718
rect 16464 4777 16498 4811
rect 16563 4785 16597 4819
rect 16635 4673 16669 4707
rect 16803 4801 16837 4835
rect 16903 4801 16937 4835
rect 16731 4673 16765 4707
rect 17332 4770 17366 4804
rect 17428 4771 17462 4805
rect 16988 4689 17022 4723
rect 17105 4689 17139 4723
rect 17596 4777 17630 4811
rect 17692 4777 17726 4811
rect 17518 4666 17552 4700
rect 6244 3091 6278 3125
rect 1930 2039 1964 2073
rect 2029 2047 2063 2081
rect 2101 1935 2135 1969
rect 2269 2063 2303 2097
rect 2369 2063 2403 2097
rect 2197 1935 2231 1969
rect 2798 2032 2832 2066
rect 2894 2033 2928 2067
rect 2454 1951 2488 1985
rect 2571 1951 2605 1985
rect 3062 2039 3096 2073
rect 3158 2039 3192 2073
rect 4000 2035 4034 2069
rect 2984 1928 3018 1962
rect 4099 2043 4133 2077
rect 4171 1931 4205 1965
rect 4339 2059 4373 2093
rect 4439 2059 4473 2093
rect 4267 1931 4301 1965
rect 4868 2028 4902 2062
rect 4964 2029 4998 2063
rect 4524 1947 4558 1981
rect 4641 1947 4675 1981
rect 5132 2035 5166 2069
rect 5228 2035 5262 2069
rect 5952 2035 5986 2069
rect 6051 2043 6085 2077
rect 5054 1924 5088 1958
rect 6123 1931 6157 1965
rect 6291 2059 6325 2093
rect 6391 2059 6425 2093
rect 6219 1931 6253 1965
rect 6820 2028 6854 2062
rect 6916 2029 6950 2063
rect 6476 1947 6510 1981
rect 6593 1947 6627 1981
rect 7084 2035 7118 2069
rect 7180 2035 7214 2069
rect 7954 2041 7988 2075
rect 8053 2049 8087 2083
rect 7006 1924 7040 1958
rect 8125 1937 8159 1971
rect 8293 2065 8327 2099
rect 8393 2065 8427 2099
rect 8221 1937 8255 1971
rect 8822 2034 8856 2068
rect 8918 2035 8952 2069
rect 8478 1953 8512 1987
rect 8595 1953 8629 1987
rect 9086 2041 9120 2075
rect 9182 2041 9216 2075
rect 9906 2041 9940 2075
rect 10005 2049 10039 2083
rect 9008 1930 9042 1964
rect 10077 1937 10111 1971
rect 10245 2065 10279 2099
rect 10345 2065 10379 2099
rect 10173 1937 10207 1971
rect 10774 2034 10808 2068
rect 10870 2035 10904 2069
rect 10430 1953 10464 1987
rect 10547 1953 10581 1987
rect 11038 2041 11072 2075
rect 11134 2041 11168 2075
rect 11898 2041 11932 2075
rect 11997 2049 12031 2083
rect 10960 1930 10994 1964
rect 12069 1937 12103 1971
rect 12237 2065 12271 2099
rect 12337 2065 12371 2099
rect 12165 1937 12199 1971
rect 12766 2034 12800 2068
rect 12862 2035 12896 2069
rect 12422 1953 12456 1987
rect 12539 1953 12573 1987
rect 13030 2041 13064 2075
rect 13126 2041 13160 2075
rect 13850 2041 13884 2075
rect 13949 2049 13983 2083
rect 12952 1930 12986 1964
rect 14021 1937 14055 1971
rect 14189 2065 14223 2099
rect 14289 2065 14323 2099
rect 14117 1937 14151 1971
rect 14718 2034 14752 2068
rect 14814 2035 14848 2069
rect 14374 1953 14408 1987
rect 14491 1953 14525 1987
rect 14982 2041 15016 2075
rect 15078 2041 15112 2075
rect 15914 2041 15948 2075
rect 16013 2049 16047 2083
rect 14904 1930 14938 1964
rect 16085 1937 16119 1971
rect 16253 2065 16287 2099
rect 16353 2065 16387 2099
rect 16181 1937 16215 1971
rect 16782 2034 16816 2068
rect 16878 2035 16912 2069
rect 16438 1953 16472 1987
rect 16555 1953 16589 1987
rect 17046 2041 17080 2075
rect 17142 2041 17176 2075
rect 16968 1930 17002 1964
<< locali >>
rect 18579 43493 18613 43510
rect 19123 43493 19157 43510
rect 18579 43481 18846 43493
rect 18613 43447 18684 43481
rect 18718 43447 18777 43481
rect 18811 43447 18846 43481
rect 18579 43435 18846 43447
rect 18978 43481 19157 43493
rect 18978 43447 18995 43481
rect 19029 43447 19123 43481
rect 18978 43435 19157 43447
rect 18579 43391 18613 43435
rect 19123 43391 19157 43435
rect 18613 43374 18773 43382
rect 18613 43357 18655 43374
rect 18579 43340 18655 43357
rect 18689 43340 18723 43374
rect 18757 43340 18773 43374
rect 18963 43374 19123 43382
rect 18963 43340 18979 43374
rect 19013 43340 19047 43374
rect 19081 43357 19123 43374
rect 19081 43340 19157 43357
rect 18579 43299 18613 43340
rect 18579 43207 18613 43265
rect 18647 43294 19089 43306
rect 18647 43290 18882 43294
rect 18647 43256 18655 43290
rect 18689 43256 18723 43290
rect 18757 43256 18793 43290
rect 18827 43258 18882 43290
rect 18916 43290 19089 43294
rect 18916 43258 18979 43290
rect 18827 43256 18979 43258
rect 19013 43256 19047 43290
rect 19081 43256 19089 43290
rect 18647 43240 19089 43256
rect 19123 43299 19157 43340
rect 18613 43173 18655 43206
rect 18579 43172 18655 43173
rect 18689 43172 18723 43206
rect 18757 43172 18773 43206
rect 18579 43115 18613 43172
rect 18807 43138 18841 43240
rect 18579 43038 18613 43081
rect 18647 43122 18841 43138
rect 18647 43088 18655 43122
rect 18689 43088 18723 43122
rect 18757 43088 18793 43122
rect 18827 43088 18841 43122
rect 18647 43072 18841 43088
rect 18579 43023 18655 43038
rect 18613 43004 18655 43023
rect 18689 43004 18723 43038
rect 18757 43004 18773 43038
rect 18579 42931 18613 42989
rect 18807 42970 18841 43072
rect 18959 43138 18997 43240
rect 19123 43207 19157 43265
rect 19031 43172 19047 43206
rect 19081 43173 19123 43206
rect 19081 43172 19157 43173
rect 18959 43122 19089 43138
rect 18959 43088 18979 43122
rect 19013 43088 19047 43122
rect 19081 43088 19089 43122
rect 18959 43072 19089 43088
rect 19123 43115 19157 43172
rect 18647 42954 18841 42970
rect 18647 42920 18655 42954
rect 18689 42920 18723 42954
rect 18757 42920 18793 42954
rect 18827 42920 18841 42954
rect 18647 42904 18841 42920
rect 18579 42870 18613 42897
rect 18579 42839 18655 42870
rect 18613 42836 18655 42839
rect 18689 42836 18723 42870
rect 18757 42836 18773 42870
rect 18579 42747 18613 42805
rect 18807 42802 18841 42904
rect 18647 42786 18841 42802
rect 18647 42752 18655 42786
rect 18689 42752 18723 42786
rect 18757 42752 18793 42786
rect 18827 42752 18841 42786
rect 18647 42736 18841 42752
rect 18579 42702 18613 42713
rect 18579 42668 18655 42702
rect 18689 42668 18723 42702
rect 18757 42668 18773 42702
rect 18579 42655 18613 42668
rect 18807 42634 18841 42736
rect 18579 42563 18613 42621
rect 18647 42618 18841 42634
rect 18647 42584 18655 42618
rect 18689 42584 18723 42618
rect 18757 42584 18793 42618
rect 18827 42584 18841 42618
rect 18647 42568 18841 42584
rect 18613 42529 18655 42534
rect 18579 42500 18655 42529
rect 18689 42500 18723 42534
rect 18757 42500 18773 42534
rect 18579 42471 18613 42500
rect 18807 42466 18841 42568
rect 18579 42379 18613 42437
rect 18647 42450 18841 42466
rect 18647 42416 18655 42450
rect 18689 42416 18723 42450
rect 18757 42416 18793 42450
rect 18827 42416 18841 42450
rect 18647 42400 18841 42416
rect 18613 42345 18655 42366
rect 18579 42332 18655 42345
rect 18689 42332 18723 42366
rect 18757 42332 18773 42366
rect 18579 42287 18613 42332
rect 18807 42298 18841 42400
rect 18579 42198 18613 42253
rect 18647 42282 18841 42298
rect 18647 42248 18655 42282
rect 18689 42248 18723 42282
rect 18757 42248 18793 42282
rect 18827 42248 18841 42282
rect 18647 42232 18841 42248
rect 18579 42195 18655 42198
rect 18613 42164 18655 42195
rect 18689 42164 18723 42198
rect 18757 42164 18773 42198
rect 18579 42103 18613 42161
rect 18807 42130 18841 42232
rect 18579 42030 18613 42069
rect 18647 42114 18841 42130
rect 18647 42080 18655 42114
rect 18689 42080 18723 42114
rect 18757 42080 18793 42114
rect 18827 42080 18841 42114
rect 18647 42064 18841 42080
rect 18877 43037 18925 43053
rect 18877 43003 18891 43037
rect 18877 42870 18925 43003
rect 18877 42836 18891 42870
rect 18877 42702 18925 42836
rect 18877 42668 18891 42702
rect 18877 42535 18925 42668
rect 18877 42501 18891 42535
rect 18877 42366 18925 42501
rect 18877 42332 18891 42366
rect 18877 42198 18925 42332
rect 18877 42164 18891 42198
rect 18579 42011 18655 42030
rect 18613 41996 18655 42011
rect 18689 41996 18723 42030
rect 18757 41996 18793 42030
rect 18827 41996 18843 42030
rect 18613 41988 18843 41996
rect 18877 42024 18925 42164
rect 18959 42970 18997 43072
rect 19123 43038 19157 43081
rect 19031 43004 19047 43038
rect 19081 43023 19157 43038
rect 19081 43004 19123 43023
rect 18959 42954 19089 42970
rect 18959 42920 18979 42954
rect 19013 42920 19047 42954
rect 19081 42920 19089 42954
rect 18959 42904 19089 42920
rect 19123 42931 19157 42989
rect 18959 42802 18997 42904
rect 19123 42870 19157 42897
rect 19031 42836 19047 42870
rect 19081 42839 19157 42870
rect 19081 42836 19123 42839
rect 18959 42786 19089 42802
rect 18959 42752 18979 42786
rect 19013 42752 19047 42786
rect 19081 42752 19089 42786
rect 18959 42736 19089 42752
rect 19123 42747 19157 42805
rect 18959 42634 18997 42736
rect 19123 42702 19157 42713
rect 19031 42668 19047 42702
rect 19081 42668 19157 42702
rect 19123 42655 19157 42668
rect 18959 42618 19089 42634
rect 18959 42584 18979 42618
rect 19013 42584 19047 42618
rect 19081 42584 19089 42618
rect 18959 42568 19089 42584
rect 18959 42466 18997 42568
rect 19123 42563 19157 42621
rect 19031 42500 19047 42534
rect 19081 42529 19123 42534
rect 19081 42500 19157 42529
rect 19123 42471 19157 42500
rect 18959 42450 19089 42466
rect 18959 42416 18979 42450
rect 19013 42416 19047 42450
rect 19081 42416 19089 42450
rect 18959 42400 19089 42416
rect 18959 42298 18997 42400
rect 19123 42379 19157 42437
rect 19031 42332 19047 42366
rect 19081 42345 19123 42366
rect 19081 42332 19157 42345
rect 18959 42282 19089 42298
rect 18959 42248 18979 42282
rect 19013 42248 19047 42282
rect 19081 42248 19089 42282
rect 18959 42232 19089 42248
rect 19123 42287 19157 42332
rect 18959 42130 18997 42232
rect 19123 42198 19157 42253
rect 19031 42164 19047 42198
rect 19081 42195 19157 42198
rect 19081 42164 19123 42195
rect 18959 42114 19089 42130
rect 18959 42080 18979 42114
rect 19013 42080 19047 42114
rect 19081 42080 19089 42114
rect 18959 42064 19089 42080
rect 19123 42103 19157 42161
rect 19123 42030 19157 42069
rect 18877 41990 18886 42024
rect 18579 41948 18613 41977
rect 18877 41965 18925 41990
rect 18963 41996 18979 42030
rect 19013 41996 19047 42030
rect 19081 42011 19157 42030
rect 19081 41996 19123 42011
rect 18963 41984 19123 41996
rect 19123 41948 19157 41977
rect 18563 41507 18597 41524
rect 19107 41507 19141 41524
rect 18563 41495 18830 41507
rect 18597 41461 18668 41495
rect 18702 41461 18761 41495
rect 18795 41461 18830 41495
rect 18563 41449 18830 41461
rect 18962 41495 19141 41507
rect 18962 41461 18979 41495
rect 19013 41461 19107 41495
rect 18962 41449 19141 41461
rect 18563 41415 18597 41449
rect 19107 41415 19141 41449
rect 18563 41403 18757 41415
rect 18597 41397 18757 41403
rect 18597 41369 18639 41397
rect 18563 41363 18639 41369
rect 18673 41363 18707 41397
rect 18741 41363 18757 41397
rect 18563 41347 18757 41363
rect 18791 41398 18981 41415
rect 18791 41364 18868 41398
rect 18902 41364 18981 41398
rect 18563 41311 18597 41347
rect 18791 41345 18981 41364
rect 19015 41403 19141 41415
rect 19015 41397 19107 41403
rect 19015 41363 19031 41397
rect 19065 41369 19107 41397
rect 19065 41363 19141 41369
rect 19015 41347 19141 41363
rect 18791 41278 18825 41345
rect 18563 41219 18597 41277
rect 18631 41262 18825 41278
rect 18631 41228 18639 41262
rect 18673 41228 18707 41262
rect 18741 41228 18775 41262
rect 18809 41228 18825 41262
rect 18631 41212 18825 41228
rect 18563 41178 18597 41185
rect 18563 41144 18639 41178
rect 18673 41144 18707 41178
rect 18741 41144 18757 41178
rect 18563 41127 18597 41144
rect 18791 41110 18825 41212
rect 18563 41035 18597 41093
rect 18631 41094 18825 41110
rect 18631 41060 18639 41094
rect 18673 41060 18707 41094
rect 18741 41060 18775 41094
rect 18809 41060 18825 41094
rect 18631 41044 18825 41060
rect 18597 41001 18639 41010
rect 18563 40976 18639 41001
rect 18673 40976 18707 41010
rect 18741 40976 18757 41010
rect 18563 40943 18597 40976
rect 18791 40942 18825 41044
rect 18563 40851 18597 40909
rect 18631 40926 18825 40942
rect 18631 40892 18639 40926
rect 18673 40892 18707 40926
rect 18741 40892 18775 40926
rect 18809 40892 18825 40926
rect 18631 40876 18825 40892
rect 18597 40817 18639 40842
rect 18563 40808 18639 40817
rect 18673 40808 18707 40842
rect 18741 40808 18757 40842
rect 18563 40759 18597 40808
rect 18791 40774 18825 40876
rect 18563 40674 18597 40725
rect 18631 40758 18825 40774
rect 18631 40724 18639 40758
rect 18673 40724 18707 40758
rect 18741 40724 18775 40758
rect 18809 40724 18825 40758
rect 18631 40708 18825 40724
rect 18563 40667 18639 40674
rect 18597 40640 18639 40667
rect 18673 40640 18707 40674
rect 18741 40640 18757 40674
rect 18563 40575 18597 40633
rect 18791 40606 18825 40708
rect 18563 40506 18597 40541
rect 18631 40590 18825 40606
rect 18631 40556 18639 40590
rect 18673 40556 18707 40590
rect 18741 40556 18775 40590
rect 18809 40556 18825 40590
rect 18631 40540 18825 40556
rect 18563 40483 18639 40506
rect 18597 40472 18639 40483
rect 18673 40472 18707 40506
rect 18741 40472 18757 40506
rect 18563 40391 18597 40449
rect 18791 40438 18825 40540
rect 18631 40422 18825 40438
rect 18631 40388 18639 40422
rect 18673 40388 18707 40422
rect 18741 40388 18775 40422
rect 18809 40388 18825 40422
rect 18631 40372 18825 40388
rect 18859 41262 18909 41290
rect 18859 41228 18875 41262
rect 18859 41178 18909 41228
rect 18859 41144 18875 41178
rect 18859 41094 18909 41144
rect 18859 41060 18875 41094
rect 18859 41010 18909 41060
rect 18859 40976 18875 41010
rect 18859 40926 18909 40976
rect 18859 40892 18875 40926
rect 18859 40842 18909 40892
rect 18859 40808 18875 40842
rect 18859 40758 18909 40808
rect 18859 40724 18875 40758
rect 18859 40674 18909 40724
rect 18859 40640 18875 40674
rect 18859 40590 18909 40640
rect 18859 40556 18875 40590
rect 18859 40506 18909 40556
rect 18859 40472 18875 40506
rect 18859 40468 18909 40472
rect 18859 40434 18870 40468
rect 18904 40434 18909 40468
rect 18859 40422 18909 40434
rect 18859 40388 18875 40422
rect 18859 40372 18909 40388
rect 18943 41278 18981 41345
rect 19107 41311 19141 41347
rect 18943 41262 19073 41278
rect 18943 41228 18963 41262
rect 18997 41228 19031 41262
rect 19065 41228 19073 41262
rect 18943 41212 19073 41228
rect 19107 41219 19141 41277
rect 18943 41110 18981 41212
rect 19107 41178 19141 41185
rect 19015 41144 19031 41178
rect 19065 41144 19141 41178
rect 19107 41127 19141 41144
rect 18943 41094 19073 41110
rect 18943 41060 18963 41094
rect 18997 41060 19031 41094
rect 19065 41060 19073 41094
rect 18943 41044 19073 41060
rect 18943 40942 18981 41044
rect 19107 41035 19141 41093
rect 19015 40976 19031 41010
rect 19065 41001 19107 41010
rect 19065 40976 19141 41001
rect 19107 40943 19141 40976
rect 18943 40926 19073 40942
rect 18943 40892 18963 40926
rect 18997 40892 19031 40926
rect 19065 40892 19073 40926
rect 18943 40876 19073 40892
rect 18943 40774 18981 40876
rect 19107 40851 19141 40909
rect 19015 40808 19031 40842
rect 19065 40817 19107 40842
rect 19065 40808 19141 40817
rect 18943 40758 19073 40774
rect 18943 40724 18963 40758
rect 18997 40724 19031 40758
rect 19065 40724 19073 40758
rect 18943 40708 19073 40724
rect 19107 40759 19141 40808
rect 18943 40606 18981 40708
rect 19107 40674 19141 40725
rect 19015 40640 19031 40674
rect 19065 40667 19141 40674
rect 19065 40640 19107 40667
rect 18943 40590 19073 40606
rect 18943 40556 18963 40590
rect 18997 40556 19031 40590
rect 19065 40556 19073 40590
rect 18943 40540 19073 40556
rect 19107 40575 19141 40633
rect 18943 40438 18981 40540
rect 19107 40506 19141 40541
rect 19015 40472 19031 40506
rect 19065 40483 19141 40506
rect 19065 40472 19107 40483
rect 18943 40422 19073 40438
rect 18943 40388 18963 40422
rect 18997 40388 19031 40422
rect 19065 40388 19073 40422
rect 18943 40372 19073 40388
rect 19107 40391 19141 40449
rect 18563 40338 18597 40357
rect 18791 40338 18825 40372
rect 18943 40338 18981 40372
rect 19107 40338 19141 40357
rect 18563 40304 18639 40338
rect 18673 40304 18707 40338
rect 18741 40304 18757 40338
rect 18563 40299 18757 40304
rect 18597 40287 18757 40299
rect 18563 40236 18597 40265
rect 18791 40253 18981 40338
rect 19015 40304 19031 40338
rect 19065 40304 19141 40338
rect 19015 40299 19141 40304
rect 19015 40287 19107 40299
rect 19107 40236 19141 40265
rect 18571 39711 18605 39728
rect 19115 39711 19149 39728
rect 18571 39699 18838 39711
rect 18605 39665 18676 39699
rect 18710 39665 18769 39699
rect 18803 39665 18838 39699
rect 18571 39653 18838 39665
rect 18970 39699 19149 39711
rect 18970 39665 18987 39699
rect 19021 39665 19115 39699
rect 18970 39653 19149 39665
rect 18571 39608 18605 39653
rect 18571 39607 18765 39608
rect 18605 39582 18765 39607
rect 18605 39573 18647 39582
rect 18571 39548 18647 39573
rect 18681 39548 18715 39582
rect 18749 39548 18765 39582
rect 18799 39606 18989 39619
rect 19115 39609 19149 39653
rect 18799 39570 18862 39606
rect 18896 39570 18989 39606
rect 18799 39555 18989 39570
rect 18571 39515 18605 39548
rect 18799 39514 18833 39555
rect 18571 39423 18605 39481
rect 18639 39498 18833 39514
rect 18639 39464 18647 39498
rect 18681 39464 18715 39498
rect 18749 39464 18783 39498
rect 18817 39464 18833 39498
rect 18639 39448 18833 39464
rect 18605 39389 18647 39414
rect 18571 39380 18647 39389
rect 18681 39380 18715 39414
rect 18749 39380 18765 39414
rect 18571 39331 18605 39380
rect 18799 39346 18833 39448
rect 18571 39246 18605 39297
rect 18639 39330 18833 39346
rect 18639 39296 18647 39330
rect 18681 39296 18715 39330
rect 18749 39296 18783 39330
rect 18817 39296 18833 39330
rect 18639 39280 18833 39296
rect 18571 39239 18647 39246
rect 18605 39212 18647 39239
rect 18681 39212 18715 39246
rect 18749 39212 18765 39246
rect 18571 39147 18605 39205
rect 18799 39178 18833 39280
rect 18571 39078 18605 39113
rect 18639 39162 18833 39178
rect 18639 39128 18647 39162
rect 18681 39128 18715 39162
rect 18749 39128 18783 39162
rect 18817 39128 18833 39162
rect 18639 39112 18833 39128
rect 18571 39055 18647 39078
rect 18605 39044 18647 39055
rect 18681 39044 18715 39078
rect 18749 39044 18765 39078
rect 18571 38963 18605 39021
rect 18799 39010 18833 39112
rect 18639 38994 18833 39010
rect 18639 38960 18647 38994
rect 18681 38960 18715 38994
rect 18749 38960 18783 38994
rect 18817 38960 18833 38994
rect 18639 38944 18833 38960
rect 18867 39498 18917 39515
rect 18867 39464 18883 39498
rect 18867 39414 18917 39464
rect 18867 39380 18883 39414
rect 18867 39330 18917 39380
rect 18867 39296 18883 39330
rect 18867 39246 18917 39296
rect 18867 39212 18883 39246
rect 18867 39162 18917 39212
rect 18867 39128 18883 39162
rect 18867 39090 18917 39128
rect 18867 39056 18876 39090
rect 18910 39078 18917 39090
rect 18867 39044 18883 39056
rect 18867 38994 18917 39044
rect 18867 38960 18883 38994
rect 18867 38944 18917 38960
rect 18951 39514 18989 39555
rect 19023 39607 19149 39609
rect 19023 39582 19115 39607
rect 19023 39548 19039 39582
rect 19073 39573 19115 39582
rect 19073 39548 19149 39573
rect 19115 39515 19149 39548
rect 18951 39498 19081 39514
rect 18951 39464 18971 39498
rect 19005 39464 19039 39498
rect 19073 39464 19081 39498
rect 18951 39448 19081 39464
rect 18951 39346 18989 39448
rect 19115 39423 19149 39481
rect 19023 39380 19039 39414
rect 19073 39389 19115 39414
rect 19073 39380 19149 39389
rect 18951 39330 19081 39346
rect 18951 39296 18971 39330
rect 19005 39296 19039 39330
rect 19073 39296 19081 39330
rect 18951 39280 19081 39296
rect 19115 39331 19149 39380
rect 18951 39178 18989 39280
rect 19115 39246 19149 39297
rect 19023 39212 19039 39246
rect 19073 39239 19149 39246
rect 19073 39212 19115 39239
rect 18951 39162 19081 39178
rect 18951 39128 18971 39162
rect 19005 39128 19039 39162
rect 19073 39128 19081 39162
rect 18951 39112 19081 39128
rect 19115 39147 19149 39205
rect 18951 39010 18989 39112
rect 19115 39078 19149 39113
rect 19023 39044 19039 39078
rect 19073 39055 19149 39078
rect 19073 39044 19115 39055
rect 18951 38994 19081 39010
rect 18951 38960 18971 38994
rect 19005 38960 19039 38994
rect 19073 38960 19081 38994
rect 18951 38944 19081 38960
rect 19115 38963 19149 39021
rect 18571 38910 18605 38929
rect 18571 38876 18647 38910
rect 18681 38876 18715 38910
rect 18749 38876 18765 38910
rect 18571 38871 18765 38876
rect 18605 38859 18765 38871
rect 18799 38894 18833 38944
rect 18951 38894 18989 38944
rect 19115 38910 19149 38929
rect 18571 38808 18605 38837
rect 18799 38825 18989 38894
rect 19023 38876 19039 38910
rect 19073 38876 19149 38910
rect 19023 38871 19149 38876
rect 19023 38859 19115 38871
rect 19115 38808 19149 38837
rect 18585 38449 18619 38466
rect 19129 38449 19163 38466
rect 18585 38437 18852 38449
rect 18619 38403 18690 38437
rect 18724 38403 18783 38437
rect 18817 38403 18852 38437
rect 18585 38391 18852 38403
rect 18984 38437 19163 38449
rect 18984 38403 19001 38437
rect 19035 38403 19129 38437
rect 18984 38391 19163 38403
rect 18585 38345 18619 38391
rect 18809 38340 19001 38357
rect 18619 38311 18661 38337
rect 18585 38303 18661 38311
rect 18695 38303 18711 38337
rect 18809 38306 18886 38340
rect 18920 38306 19001 38340
rect 19129 38345 19163 38391
rect 18585 38253 18619 38303
rect 18809 38287 19001 38306
rect 19036 38303 19052 38337
rect 19086 38311 19129 38337
rect 19086 38303 19163 38311
rect 19036 38287 19163 38303
rect 18809 38269 18847 38287
rect 18585 38169 18619 38219
rect 18653 38253 18847 38269
rect 18965 38253 19001 38287
rect 19129 38253 19163 38287
rect 18653 38219 18661 38253
rect 18695 38219 18729 38253
rect 18763 38219 18797 38253
rect 18831 38219 18847 38253
rect 18653 38203 18847 38219
rect 18585 38161 18661 38169
rect 18619 38135 18661 38161
rect 18695 38135 18729 38169
rect 18763 38135 18779 38169
rect 18585 38069 18619 38127
rect 18813 38101 18847 38203
rect 18653 38085 18847 38101
rect 18653 38051 18661 38085
rect 18695 38051 18729 38085
rect 18763 38051 18797 38085
rect 18831 38051 18847 38085
rect 18653 38035 18847 38051
rect 18585 38001 18619 38035
rect 18585 37977 18661 38001
rect 18619 37967 18661 37977
rect 18695 37967 18729 38001
rect 18763 37967 18779 38001
rect 18585 37885 18619 37943
rect 18813 37933 18847 38035
rect 18653 37917 18847 37933
rect 18653 37883 18661 37917
rect 18695 37883 18729 37917
rect 18763 37883 18797 37917
rect 18831 37883 18847 37917
rect 18653 37867 18847 37883
rect 18881 38237 18931 38253
rect 18881 38203 18897 38237
rect 18881 38153 18931 38203
rect 18881 38119 18897 38153
rect 18881 38069 18931 38119
rect 18881 38035 18897 38069
rect 18585 37815 18619 37851
rect 18585 37799 18847 37815
rect 18585 37793 18661 37799
rect 18619 37765 18661 37793
rect 18695 37765 18729 37799
rect 18763 37765 18797 37799
rect 18831 37765 18847 37799
rect 18619 37759 18847 37765
rect 18585 37756 18847 37759
rect 18881 37801 18931 38035
rect 18965 38219 19045 38253
rect 19079 38219 19095 38253
rect 18965 38085 19001 38219
rect 19129 38169 19163 38219
rect 19037 38135 19053 38169
rect 19087 38161 19163 38169
rect 19087 38135 19129 38161
rect 18965 38051 19045 38085
rect 19079 38051 19095 38085
rect 19129 38069 19163 38127
rect 18965 37917 19001 38051
rect 19129 38001 19163 38035
rect 19037 37967 19053 38001
rect 19087 37977 19163 38001
rect 19087 37967 19129 37977
rect 18965 37883 19045 37917
rect 19079 37883 19095 37917
rect 19129 37885 19163 37943
rect 19129 37809 19163 37851
rect 18881 37794 18897 37801
rect 18881 37760 18888 37794
rect 18922 37760 18931 37767
rect 18585 37730 18619 37756
rect 18881 37751 18931 37760
rect 19037 37775 19053 37809
rect 19087 37793 19163 37809
rect 19087 37775 19129 37793
rect 19037 37759 19129 37775
rect 19037 37756 19163 37759
rect 19129 37730 19163 37756
rect 18597 37295 18631 37312
rect 19141 37295 19175 37312
rect 18597 37283 18864 37295
rect 18631 37249 18702 37283
rect 18736 37249 18795 37283
rect 18829 37249 18864 37283
rect 18597 37237 18864 37249
rect 18996 37283 19175 37295
rect 18996 37249 19013 37283
rect 19047 37249 19141 37283
rect 18996 37237 19175 37249
rect 18597 37195 18631 37237
rect 18821 37192 19013 37198
rect 19141 37195 19175 37237
rect 18631 37179 18723 37187
rect 18631 37161 18673 37179
rect 18597 37145 18673 37161
rect 18707 37145 18723 37179
rect 18821 37158 18892 37192
rect 18926 37158 19013 37192
rect 18821 37145 19013 37158
rect 19048 37179 19141 37195
rect 19048 37145 19064 37179
rect 19098 37161 19141 37179
rect 19098 37145 19175 37161
rect 18597 37103 18631 37145
rect 18821 37111 18859 37145
rect 18977 37111 19013 37145
rect 18597 37011 18631 37069
rect 18665 37095 18859 37111
rect 18665 37061 18673 37095
rect 18707 37061 18741 37095
rect 18775 37061 18809 37095
rect 18843 37061 18859 37095
rect 18665 37045 18859 37061
rect 18631 36977 18673 37011
rect 18707 36977 18741 37011
rect 18775 36977 18791 37011
rect 18597 36919 18631 36977
rect 18825 36943 18859 37045
rect 18597 36843 18631 36885
rect 18665 36927 18859 36943
rect 18665 36893 18673 36927
rect 18707 36893 18741 36927
rect 18775 36893 18809 36927
rect 18843 36893 18859 36927
rect 18665 36877 18859 36893
rect 18893 37095 18943 37111
rect 18893 37061 18909 37095
rect 18893 37011 18943 37061
rect 18893 36977 18909 37011
rect 18893 36927 18943 36977
rect 18893 36920 18909 36927
rect 18893 36884 18900 36920
rect 18934 36884 18943 36893
rect 18597 36827 18673 36843
rect 18631 36809 18673 36827
rect 18707 36809 18741 36843
rect 18775 36809 18809 36843
rect 18843 36809 18859 36843
rect 18631 36793 18859 36809
rect 18597 36790 18859 36793
rect 18893 36835 18943 36884
rect 18977 37095 19107 37111
rect 18977 37061 19057 37095
rect 19091 37061 19107 37095
rect 18977 37045 19107 37061
rect 19141 37103 19175 37145
rect 18977 36943 19013 37045
rect 19141 37011 19175 37069
rect 19049 36977 19065 37011
rect 19099 36977 19141 37011
rect 18977 36927 19107 36943
rect 18977 36893 19057 36927
rect 19091 36893 19107 36927
rect 18977 36877 19107 36893
rect 19141 36919 19175 36977
rect 19141 36843 19175 36885
rect 18893 36801 18909 36835
rect 18597 36764 18631 36790
rect 18893 36785 18943 36801
rect 19049 36809 19065 36843
rect 19099 36827 19175 36843
rect 19099 36809 19141 36827
rect 19049 36793 19141 36809
rect 19049 36790 19175 36793
rect 19141 36764 19175 36790
rect 18605 36411 18639 36428
rect 19149 36411 19183 36428
rect 18605 36399 18872 36411
rect 18639 36365 18710 36399
rect 18744 36365 18803 36399
rect 18837 36365 18872 36399
rect 18605 36353 18872 36365
rect 19004 36399 19183 36411
rect 19004 36365 19021 36399
rect 19055 36365 19149 36399
rect 19004 36353 19183 36365
rect 18605 36307 18639 36353
rect 19149 36307 19183 36353
rect 18639 36299 18867 36307
rect 18639 36273 18681 36299
rect 18605 36265 18681 36273
rect 18715 36265 18749 36299
rect 18783 36265 18817 36299
rect 18851 36265 18867 36299
rect 18985 36299 19149 36307
rect 18985 36265 19001 36299
rect 19035 36265 19073 36299
rect 19107 36273 19149 36299
rect 19107 36265 19183 36273
rect 18605 36215 18639 36265
rect 18605 36131 18639 36181
rect 18673 36226 19115 36231
rect 18673 36215 18904 36226
rect 18673 36181 18681 36215
rect 18715 36181 18749 36215
rect 18783 36181 18817 36215
rect 18851 36190 18904 36215
rect 18940 36215 19115 36226
rect 18940 36190 19001 36215
rect 18851 36181 19001 36190
rect 19035 36181 19073 36215
rect 19107 36181 19115 36215
rect 18673 36165 18869 36181
rect 18989 36165 19115 36181
rect 19149 36215 19183 36265
rect 18901 36131 18951 36147
rect 19149 36131 19183 36181
rect 18605 36123 18681 36131
rect 18639 36097 18681 36123
rect 18715 36097 18749 36131
rect 18783 36097 18817 36131
rect 18851 36097 18867 36131
rect 18639 36089 18867 36097
rect 18605 36085 18867 36089
rect 18901 36130 18917 36131
rect 18901 36094 18904 36130
rect 18948 36094 18951 36097
rect 18605 36060 18639 36085
rect 18901 36081 18951 36094
rect 18985 36097 19001 36131
rect 19035 36097 19073 36131
rect 19107 36123 19183 36131
rect 19107 36097 19149 36123
rect 18985 36089 19149 36097
rect 18985 36085 19183 36089
rect 19149 36060 19183 36085
rect 18629 35023 18663 35040
rect 19173 35023 19207 35040
rect 18629 35011 18896 35023
rect 18663 34977 18734 35011
rect 18768 34977 18827 35011
rect 18861 34977 18896 35011
rect 18629 34965 18896 34977
rect 19028 35011 19207 35023
rect 19028 34977 19045 35011
rect 19079 34977 19173 35011
rect 19028 34965 19207 34977
rect 18629 34919 18663 34965
rect 18629 34829 18663 34885
rect 18697 34914 19139 34930
rect 18697 34913 18836 34914
rect 18870 34913 19139 34914
rect 18697 34879 18705 34913
rect 18739 34879 18776 34913
rect 18810 34880 18836 34913
rect 18881 34883 19059 34913
rect 18810 34879 18847 34880
rect 18881 34879 18894 34883
rect 19008 34879 19059 34883
rect 19093 34879 19139 34913
rect 19173 34919 19207 34965
rect 18697 34863 18894 34879
rect 18629 34827 18705 34829
rect 18663 34795 18705 34827
rect 18739 34795 18773 34829
rect 18807 34795 18841 34829
rect 18875 34795 18891 34829
rect 18663 34793 18891 34795
rect 18629 34786 18891 34793
rect 18925 34815 18941 34849
rect 18975 34815 18991 34849
rect 19173 34845 19207 34885
rect 18629 34735 18663 34786
rect 18925 34748 18991 34815
rect 19081 34829 19207 34845
rect 19081 34795 19097 34829
rect 19131 34827 19207 34829
rect 19131 34795 19173 34827
rect 19081 34793 19173 34795
rect 19081 34781 19207 34793
rect 18629 34643 18663 34701
rect 18701 34734 18991 34748
rect 19173 34735 19207 34781
rect 18701 34732 19071 34734
rect 18701 34698 18705 34732
rect 18739 34698 18773 34732
rect 18807 34700 19071 34732
rect 19105 34700 19121 34734
rect 18807 34698 19121 34700
rect 18701 34694 19121 34698
rect 18701 34682 18847 34694
rect 19067 34684 19121 34694
rect 18875 34646 19042 34660
rect 18875 34644 19129 34646
rect 18629 34551 18663 34609
rect 18706 34634 19129 34644
rect 18706 34630 19058 34634
rect 19092 34630 19129 34634
rect 18706 34628 19026 34630
rect 18706 34594 18711 34628
rect 18745 34594 18779 34628
rect 18813 34594 18847 34628
rect 18881 34622 19026 34628
rect 18881 34613 18901 34622
rect 18881 34594 18891 34613
rect 19017 34611 19026 34622
rect 18706 34578 18891 34594
rect 19025 34596 19026 34611
rect 19092 34600 19094 34630
rect 19060 34596 19094 34600
rect 19128 34596 19129 34630
rect 18925 34554 18941 34588
rect 18975 34554 18991 34588
rect 19025 34580 19129 34596
rect 19173 34643 19207 34701
rect 18663 34517 18735 34544
rect 18629 34510 18735 34517
rect 18769 34510 18815 34544
rect 18849 34510 18865 34544
rect 18629 34459 18663 34510
rect 18925 34478 18991 34554
rect 19173 34551 19207 34609
rect 19051 34512 19067 34546
rect 19101 34517 19173 34546
rect 19101 34512 19207 34517
rect 18925 34476 19130 34478
rect 18629 34367 18663 34425
rect 18697 34462 19130 34476
rect 18697 34458 19028 34462
rect 18697 34424 18705 34458
rect 18739 34424 18776 34458
rect 18810 34424 18847 34458
rect 18881 34438 19028 34458
rect 18881 34424 18884 34438
rect 18697 34408 18884 34424
rect 19025 34428 19028 34438
rect 19062 34428 19096 34462
rect 19025 34412 19130 34428
rect 19173 34459 19207 34512
rect 18663 34334 18763 34361
rect 18663 34333 18713 34334
rect 18629 34300 18713 34333
rect 18747 34300 18763 34334
rect 18629 34298 18763 34300
rect 18809 34330 18884 34408
rect 18629 34275 18663 34298
rect 18809 34296 18825 34330
rect 18859 34296 18884 34330
rect 18925 34370 18941 34404
rect 18975 34370 18991 34404
rect 18925 34262 18991 34370
rect 19173 34367 19207 34425
rect 19067 34356 19173 34359
rect 19067 34322 19083 34356
rect 19117 34333 19173 34356
rect 19117 34322 19207 34333
rect 19067 34317 19207 34322
rect 19173 34275 19207 34317
rect 18629 34183 18663 34241
rect 18629 34091 18663 34149
rect 18723 34228 19117 34262
rect 18723 34135 18757 34228
rect 18791 34160 18825 34194
rect 18859 34181 19049 34194
rect 18859 34160 18867 34181
rect 18791 34147 18867 34160
rect 18901 34147 19049 34181
rect 18791 34135 19049 34147
rect 18791 34130 18999 34135
rect 18983 34101 18999 34130
rect 19033 34101 19049 34135
rect 19083 34158 19117 34228
rect 19083 34105 19117 34124
rect 19173 34183 19207 34241
rect 18723 34085 18757 34101
rect 18797 34094 18941 34096
rect 18797 34060 18799 34094
rect 18833 34092 18941 34094
rect 18833 34060 18891 34092
rect 18797 34058 18891 34060
rect 18925 34058 18941 34092
rect 19173 34091 19207 34149
rect 18629 33999 18663 34057
rect 19083 34055 19117 34071
rect 18697 34006 18713 34040
rect 18747 34024 18763 34040
rect 18747 34021 19083 34024
rect 18747 34006 19117 34021
rect 18697 33990 19117 34006
rect 19173 33999 19207 34057
rect 18629 33956 18663 33965
rect 18629 33922 18705 33956
rect 18739 33922 18773 33956
rect 18807 33922 18823 33956
rect 18875 33922 18891 33956
rect 18925 33922 18941 33956
rect 18629 33907 18663 33922
rect 18875 33888 18927 33922
rect 18977 33898 19037 33990
rect 19173 33954 19207 33965
rect 18629 33815 18663 33873
rect 18629 33723 18663 33781
rect 18629 33631 18663 33689
rect 18718 33854 18927 33888
rect 18971 33892 19037 33898
rect 18971 33858 18987 33892
rect 19021 33858 19037 33892
rect 19073 33936 19207 33954
rect 19073 33902 19089 33936
rect 19123 33907 19207 33936
rect 19123 33902 19173 33907
rect 19073 33880 19173 33902
rect 18718 33717 18752 33854
rect 18786 33782 18859 33820
rect 18893 33816 18927 33854
rect 18893 33782 19117 33816
rect 18786 33780 18825 33782
rect 18786 33746 18799 33780
rect 18833 33746 19043 33748
rect 18786 33714 19043 33746
rect 18718 33667 18752 33683
rect 18999 33693 19043 33714
rect 18846 33677 18965 33680
rect 18846 33643 18867 33677
rect 18901 33673 18965 33677
rect 18901 33643 18903 33673
rect 18846 33639 18903 33643
rect 18937 33639 18965 33673
rect 19033 33659 19043 33693
rect 19083 33737 19117 33782
rect 19083 33681 19117 33703
rect 19173 33815 19207 33873
rect 19173 33723 19207 33781
rect 18999 33643 19043 33659
rect 18846 33632 18965 33639
rect 19083 33626 19117 33642
rect 18629 33541 18663 33597
rect 18697 33591 18713 33625
rect 18747 33598 18808 33625
rect 19029 33598 19083 33609
rect 18747 33592 19083 33598
rect 18747 33591 19117 33592
rect 18697 33575 19117 33591
rect 19173 33631 19207 33689
rect 18782 33564 19055 33575
rect 19173 33541 19207 33597
rect 18629 33539 18705 33541
rect 18663 33507 18705 33539
rect 18739 33507 18755 33541
rect 18663 33505 18755 33507
rect 18629 33488 18755 33505
rect 18857 33496 18873 33530
rect 18907 33524 19047 33530
rect 18907 33496 18988 33524
rect 18629 33447 18663 33488
rect 18857 33484 18988 33496
rect 19028 33484 19047 33524
rect 19081 33507 19097 33541
rect 19131 33539 19207 33541
rect 19131 33507 19173 33539
rect 19081 33505 19173 33507
rect 19081 33491 19207 33505
rect 18857 33474 19047 33484
rect 19173 33447 19207 33491
rect 18629 33369 18663 33413
rect 18697 33439 19121 33440
rect 18697 33437 18867 33439
rect 18697 33403 18713 33437
rect 18747 33403 18781 33437
rect 18815 33405 18867 33437
rect 18901 33437 19121 33439
rect 18901 33405 19071 33437
rect 18815 33403 19071 33405
rect 19105 33403 19121 33437
rect 19173 33369 19207 33413
rect 18629 33355 18763 33369
rect 18663 33353 18763 33355
rect 18663 33321 18729 33353
rect 18629 33319 18729 33321
rect 18629 33303 18763 33319
rect 18797 33360 18926 33368
rect 18797 33326 18799 33360
rect 18833 33334 18926 33360
rect 18960 33334 19063 33368
rect 18833 33326 19063 33334
rect 18797 33322 19063 33326
rect 18629 33263 18663 33303
rect 18797 33269 18831 33322
rect 18697 33235 18713 33269
rect 18747 33235 18781 33269
rect 18815 33235 18831 33269
rect 18865 33266 18995 33288
rect 18629 33200 18663 33229
rect 18865 33232 18940 33266
rect 18976 33232 18995 33266
rect 19029 33269 19063 33322
rect 19097 33355 19207 33369
rect 19097 33353 19173 33355
rect 19131 33321 19173 33353
rect 19131 33319 19207 33321
rect 19097 33303 19207 33319
rect 19029 33235 19071 33269
rect 19105 33235 19121 33269
rect 19173 33263 19207 33303
rect 18865 33218 18995 33232
rect 19173 33200 19207 33229
rect 18629 32741 18663 32758
rect 19173 32741 19207 32758
rect 18629 32729 18896 32741
rect 18663 32695 18734 32729
rect 18768 32695 18827 32729
rect 18861 32695 18896 32729
rect 18629 32683 18896 32695
rect 19028 32729 19207 32741
rect 19028 32695 19045 32729
rect 19079 32695 19173 32729
rect 19028 32683 19207 32695
rect 18629 32637 18663 32683
rect 18629 32547 18663 32603
rect 18697 32632 19139 32648
rect 18697 32631 18836 32632
rect 18870 32631 19139 32632
rect 18697 32597 18705 32631
rect 18739 32597 18776 32631
rect 18810 32598 18836 32631
rect 18881 32601 19059 32631
rect 18810 32597 18847 32598
rect 18881 32597 18894 32601
rect 19008 32597 19059 32601
rect 19093 32597 19139 32631
rect 19173 32637 19207 32683
rect 18697 32581 18894 32597
rect 18629 32545 18705 32547
rect 18663 32513 18705 32545
rect 18739 32513 18773 32547
rect 18807 32513 18841 32547
rect 18875 32513 18891 32547
rect 18663 32511 18891 32513
rect 18629 32504 18891 32511
rect 18925 32533 18941 32567
rect 18975 32533 18991 32567
rect 19173 32563 19207 32603
rect 18629 32453 18663 32504
rect 18925 32466 18991 32533
rect 19081 32547 19207 32563
rect 19081 32513 19097 32547
rect 19131 32545 19207 32547
rect 19131 32513 19173 32545
rect 19081 32511 19173 32513
rect 19081 32499 19207 32511
rect 18629 32361 18663 32419
rect 18701 32452 18991 32466
rect 19173 32453 19207 32499
rect 18701 32450 19071 32452
rect 18701 32416 18705 32450
rect 18739 32416 18773 32450
rect 18807 32418 19071 32450
rect 19105 32418 19121 32452
rect 18807 32416 19121 32418
rect 18701 32412 19121 32416
rect 18701 32400 18847 32412
rect 19067 32402 19121 32412
rect 18875 32364 19042 32378
rect 18875 32362 19129 32364
rect 18629 32269 18663 32327
rect 18706 32352 19129 32362
rect 18706 32348 19058 32352
rect 19092 32348 19129 32352
rect 18706 32346 19026 32348
rect 18706 32312 18711 32346
rect 18745 32312 18779 32346
rect 18813 32312 18847 32346
rect 18881 32340 19026 32346
rect 18881 32331 18901 32340
rect 18881 32312 18891 32331
rect 19017 32329 19026 32340
rect 18706 32296 18891 32312
rect 19025 32314 19026 32329
rect 19092 32318 19094 32348
rect 19060 32314 19094 32318
rect 19128 32314 19129 32348
rect 18925 32272 18941 32306
rect 18975 32272 18991 32306
rect 19025 32298 19129 32314
rect 19173 32361 19207 32419
rect 18663 32235 18735 32262
rect 18629 32228 18735 32235
rect 18769 32228 18815 32262
rect 18849 32228 18865 32262
rect 18629 32177 18663 32228
rect 18925 32196 18991 32272
rect 19173 32269 19207 32327
rect 19051 32230 19067 32264
rect 19101 32235 19173 32264
rect 19101 32230 19207 32235
rect 18925 32194 19130 32196
rect 18629 32085 18663 32143
rect 18697 32180 19130 32194
rect 18697 32176 19028 32180
rect 18697 32142 18705 32176
rect 18739 32142 18776 32176
rect 18810 32142 18847 32176
rect 18881 32156 19028 32176
rect 18881 32142 18884 32156
rect 18697 32126 18884 32142
rect 19025 32146 19028 32156
rect 19062 32146 19096 32180
rect 19025 32130 19130 32146
rect 19173 32177 19207 32230
rect 18663 32052 18763 32079
rect 18663 32051 18713 32052
rect 18629 32018 18713 32051
rect 18747 32018 18763 32052
rect 18629 32016 18763 32018
rect 18809 32048 18884 32126
rect 18629 31993 18663 32016
rect 18809 32014 18825 32048
rect 18859 32014 18884 32048
rect 18925 32088 18941 32122
rect 18975 32088 18991 32122
rect 18925 31980 18991 32088
rect 19173 32085 19207 32143
rect 19067 32074 19173 32077
rect 19067 32040 19083 32074
rect 19117 32051 19173 32074
rect 19117 32040 19207 32051
rect 19067 32035 19207 32040
rect 19173 31993 19207 32035
rect 18629 31901 18663 31959
rect 18629 31809 18663 31867
rect 18723 31946 19117 31980
rect 18723 31853 18757 31946
rect 18791 31878 18825 31912
rect 18859 31899 19049 31912
rect 18859 31878 18867 31899
rect 18791 31865 18867 31878
rect 18901 31865 19049 31899
rect 18791 31853 19049 31865
rect 18791 31848 18999 31853
rect 18983 31819 18999 31848
rect 19033 31819 19049 31853
rect 19083 31876 19117 31946
rect 19083 31823 19117 31842
rect 19173 31901 19207 31959
rect 18723 31803 18757 31819
rect 18797 31812 18941 31814
rect 18797 31778 18799 31812
rect 18833 31810 18941 31812
rect 18833 31778 18891 31810
rect 18797 31776 18891 31778
rect 18925 31776 18941 31810
rect 19173 31809 19207 31867
rect 18629 31717 18663 31775
rect 19083 31773 19117 31789
rect 18697 31724 18713 31758
rect 18747 31742 18763 31758
rect 18747 31739 19083 31742
rect 18747 31724 19117 31739
rect 18697 31708 19117 31724
rect 19173 31717 19207 31775
rect 18629 31674 18663 31683
rect 18629 31640 18705 31674
rect 18739 31640 18773 31674
rect 18807 31640 18823 31674
rect 18875 31640 18891 31674
rect 18925 31640 18941 31674
rect 18629 31625 18663 31640
rect 18875 31606 18927 31640
rect 18977 31616 19037 31708
rect 19173 31672 19207 31683
rect 18629 31533 18663 31591
rect 18629 31441 18663 31499
rect 18629 31349 18663 31407
rect 18718 31572 18927 31606
rect 18971 31610 19037 31616
rect 18971 31576 18987 31610
rect 19021 31576 19037 31610
rect 19073 31654 19207 31672
rect 19073 31620 19089 31654
rect 19123 31625 19207 31654
rect 19123 31620 19173 31625
rect 19073 31598 19173 31620
rect 18718 31435 18752 31572
rect 18786 31500 18859 31538
rect 18893 31534 18927 31572
rect 18893 31500 19117 31534
rect 18786 31498 18825 31500
rect 18786 31464 18799 31498
rect 18833 31464 19043 31466
rect 18786 31432 19043 31464
rect 18718 31385 18752 31401
rect 18999 31411 19043 31432
rect 18846 31395 18965 31398
rect 18846 31361 18867 31395
rect 18901 31391 18965 31395
rect 18901 31361 18903 31391
rect 18846 31357 18903 31361
rect 18937 31357 18965 31391
rect 19033 31377 19043 31411
rect 19083 31455 19117 31500
rect 19083 31399 19117 31421
rect 19173 31533 19207 31591
rect 19173 31441 19207 31499
rect 18999 31361 19043 31377
rect 18846 31350 18965 31357
rect 19083 31344 19117 31360
rect 18629 31259 18663 31315
rect 18697 31309 18713 31343
rect 18747 31316 18808 31343
rect 19029 31316 19083 31327
rect 18747 31310 19083 31316
rect 18747 31309 19117 31310
rect 18697 31293 19117 31309
rect 19173 31349 19207 31407
rect 18782 31282 19055 31293
rect 19173 31259 19207 31315
rect 18629 31257 18705 31259
rect 18663 31225 18705 31257
rect 18739 31225 18755 31259
rect 18663 31223 18755 31225
rect 18629 31206 18755 31223
rect 18857 31214 18873 31248
rect 18907 31242 19047 31248
rect 18907 31214 18988 31242
rect 18629 31165 18663 31206
rect 18857 31202 18988 31214
rect 19028 31202 19047 31242
rect 19081 31225 19097 31259
rect 19131 31257 19207 31259
rect 19131 31225 19173 31257
rect 19081 31223 19173 31225
rect 19081 31209 19207 31223
rect 18857 31192 19047 31202
rect 19173 31165 19207 31209
rect 18629 31087 18663 31131
rect 18697 31157 19121 31158
rect 18697 31155 18867 31157
rect 18697 31121 18713 31155
rect 18747 31121 18781 31155
rect 18815 31123 18867 31155
rect 18901 31155 19121 31157
rect 18901 31123 19071 31155
rect 18815 31121 19071 31123
rect 19105 31121 19121 31155
rect 19173 31087 19207 31131
rect 18629 31073 18763 31087
rect 18663 31071 18763 31073
rect 18663 31039 18729 31071
rect 18629 31037 18729 31039
rect 18629 31021 18763 31037
rect 18797 31078 18926 31086
rect 18797 31044 18799 31078
rect 18833 31052 18926 31078
rect 18960 31052 19063 31086
rect 18833 31044 19063 31052
rect 18797 31040 19063 31044
rect 18629 30981 18663 31021
rect 18797 30987 18831 31040
rect 18697 30953 18713 30987
rect 18747 30953 18781 30987
rect 18815 30953 18831 30987
rect 18865 30984 18995 31006
rect 18629 30918 18663 30947
rect 18865 30950 18940 30984
rect 18976 30950 18995 30984
rect 19029 30987 19063 31040
rect 19097 31073 19207 31087
rect 19097 31071 19173 31073
rect 19131 31039 19173 31071
rect 19131 31037 19207 31039
rect 19097 31021 19207 31037
rect 19029 30953 19071 30987
rect 19105 30953 19121 30987
rect 19173 30981 19207 31021
rect 18865 30936 18995 30950
rect 19173 30918 19207 30947
rect 18633 30495 18667 30512
rect 19177 30495 19211 30512
rect 18633 30483 18900 30495
rect 18667 30449 18738 30483
rect 18772 30449 18831 30483
rect 18865 30449 18900 30483
rect 18633 30437 18900 30449
rect 19032 30483 19211 30495
rect 19032 30449 19049 30483
rect 19083 30449 19177 30483
rect 19032 30437 19211 30449
rect 18633 30391 18667 30437
rect 18633 30301 18667 30357
rect 18701 30386 19143 30402
rect 18701 30385 18840 30386
rect 18874 30385 19143 30386
rect 18701 30351 18709 30385
rect 18743 30351 18780 30385
rect 18814 30352 18840 30385
rect 18885 30355 19063 30385
rect 18814 30351 18851 30352
rect 18885 30351 18898 30355
rect 19012 30351 19063 30355
rect 19097 30351 19143 30385
rect 19177 30391 19211 30437
rect 18701 30335 18898 30351
rect 18633 30299 18709 30301
rect 18667 30267 18709 30299
rect 18743 30267 18777 30301
rect 18811 30267 18845 30301
rect 18879 30267 18895 30301
rect 18667 30265 18895 30267
rect 18633 30258 18895 30265
rect 18929 30287 18945 30321
rect 18979 30287 18995 30321
rect 19177 30317 19211 30357
rect 18633 30207 18667 30258
rect 18929 30220 18995 30287
rect 19085 30301 19211 30317
rect 19085 30267 19101 30301
rect 19135 30299 19211 30301
rect 19135 30267 19177 30299
rect 19085 30265 19177 30267
rect 19085 30253 19211 30265
rect 18633 30115 18667 30173
rect 18705 30206 18995 30220
rect 19177 30207 19211 30253
rect 18705 30204 19075 30206
rect 18705 30170 18709 30204
rect 18743 30170 18777 30204
rect 18811 30172 19075 30204
rect 19109 30172 19125 30206
rect 18811 30170 19125 30172
rect 18705 30166 19125 30170
rect 18705 30154 18851 30166
rect 19071 30156 19125 30166
rect 18879 30118 19046 30132
rect 18879 30116 19133 30118
rect 18633 30023 18667 30081
rect 18710 30106 19133 30116
rect 18710 30102 19062 30106
rect 19096 30102 19133 30106
rect 18710 30100 19030 30102
rect 18710 30066 18715 30100
rect 18749 30066 18783 30100
rect 18817 30066 18851 30100
rect 18885 30094 19030 30100
rect 18885 30085 18905 30094
rect 18885 30066 18895 30085
rect 19021 30083 19030 30094
rect 18710 30050 18895 30066
rect 19029 30068 19030 30083
rect 19096 30072 19098 30102
rect 19064 30068 19098 30072
rect 19132 30068 19133 30102
rect 18929 30026 18945 30060
rect 18979 30026 18995 30060
rect 19029 30052 19133 30068
rect 19177 30115 19211 30173
rect 18667 29989 18739 30016
rect 18633 29982 18739 29989
rect 18773 29982 18819 30016
rect 18853 29982 18869 30016
rect 18633 29931 18667 29982
rect 18929 29950 18995 30026
rect 19177 30023 19211 30081
rect 19055 29984 19071 30018
rect 19105 29989 19177 30018
rect 19105 29984 19211 29989
rect 18929 29948 19134 29950
rect 18633 29839 18667 29897
rect 18701 29934 19134 29948
rect 18701 29930 19032 29934
rect 18701 29896 18709 29930
rect 18743 29896 18780 29930
rect 18814 29896 18851 29930
rect 18885 29910 19032 29930
rect 18885 29896 18888 29910
rect 18701 29880 18888 29896
rect 19029 29900 19032 29910
rect 19066 29900 19100 29934
rect 19029 29884 19134 29900
rect 19177 29931 19211 29984
rect 18667 29806 18767 29833
rect 18667 29805 18717 29806
rect 18633 29772 18717 29805
rect 18751 29772 18767 29806
rect 18633 29770 18767 29772
rect 18813 29802 18888 29880
rect 18633 29747 18667 29770
rect 18813 29768 18829 29802
rect 18863 29768 18888 29802
rect 18929 29842 18945 29876
rect 18979 29842 18995 29876
rect 18929 29734 18995 29842
rect 19177 29839 19211 29897
rect 19071 29828 19177 29831
rect 19071 29794 19087 29828
rect 19121 29805 19177 29828
rect 19121 29794 19211 29805
rect 19071 29789 19211 29794
rect 19177 29747 19211 29789
rect 18633 29655 18667 29713
rect 18633 29563 18667 29621
rect 18727 29700 19121 29734
rect 18727 29607 18761 29700
rect 18795 29632 18829 29666
rect 18863 29653 19053 29666
rect 18863 29632 18871 29653
rect 18795 29619 18871 29632
rect 18905 29619 19053 29653
rect 18795 29607 19053 29619
rect 18795 29602 19003 29607
rect 18987 29573 19003 29602
rect 19037 29573 19053 29607
rect 19087 29630 19121 29700
rect 19087 29577 19121 29596
rect 19177 29655 19211 29713
rect 18727 29557 18761 29573
rect 18801 29566 18945 29568
rect 18801 29532 18803 29566
rect 18837 29564 18945 29566
rect 18837 29532 18895 29564
rect 18801 29530 18895 29532
rect 18929 29530 18945 29564
rect 19177 29563 19211 29621
rect 18633 29471 18667 29529
rect 19087 29527 19121 29543
rect 18701 29478 18717 29512
rect 18751 29496 18767 29512
rect 18751 29493 19087 29496
rect 18751 29478 19121 29493
rect 18701 29462 19121 29478
rect 19177 29471 19211 29529
rect 18633 29428 18667 29437
rect 18633 29394 18709 29428
rect 18743 29394 18777 29428
rect 18811 29394 18827 29428
rect 18879 29394 18895 29428
rect 18929 29394 18945 29428
rect 18633 29379 18667 29394
rect 18879 29360 18931 29394
rect 18981 29370 19041 29462
rect 19177 29426 19211 29437
rect 18633 29287 18667 29345
rect 18633 29195 18667 29253
rect 18633 29103 18667 29161
rect 18722 29326 18931 29360
rect 18975 29364 19041 29370
rect 18975 29330 18991 29364
rect 19025 29330 19041 29364
rect 19077 29408 19211 29426
rect 19077 29374 19093 29408
rect 19127 29379 19211 29408
rect 19127 29374 19177 29379
rect 19077 29352 19177 29374
rect 18722 29189 18756 29326
rect 18790 29254 18863 29292
rect 18897 29288 18931 29326
rect 18897 29254 19121 29288
rect 18790 29252 18829 29254
rect 18790 29218 18803 29252
rect 18837 29218 19047 29220
rect 18790 29186 19047 29218
rect 18722 29139 18756 29155
rect 19003 29165 19047 29186
rect 18850 29149 18969 29152
rect 18850 29115 18871 29149
rect 18905 29145 18969 29149
rect 18905 29115 18907 29145
rect 18850 29111 18907 29115
rect 18941 29111 18969 29145
rect 19037 29131 19047 29165
rect 19087 29209 19121 29254
rect 19087 29153 19121 29175
rect 19177 29287 19211 29345
rect 19177 29195 19211 29253
rect 19003 29115 19047 29131
rect 18850 29104 18969 29111
rect 19087 29098 19121 29114
rect 18633 29013 18667 29069
rect 18701 29063 18717 29097
rect 18751 29070 18812 29097
rect 19033 29070 19087 29081
rect 18751 29064 19087 29070
rect 18751 29063 19121 29064
rect 18701 29047 19121 29063
rect 19177 29103 19211 29161
rect 18786 29036 19059 29047
rect 19177 29013 19211 29069
rect 18633 29011 18709 29013
rect 18667 28979 18709 29011
rect 18743 28979 18759 29013
rect 18667 28977 18759 28979
rect 18633 28960 18759 28977
rect 18861 28968 18877 29002
rect 18911 28996 19051 29002
rect 18911 28968 18992 28996
rect 18633 28919 18667 28960
rect 18861 28956 18992 28968
rect 19032 28956 19051 28996
rect 19085 28979 19101 29013
rect 19135 29011 19211 29013
rect 19135 28979 19177 29011
rect 19085 28977 19177 28979
rect 19085 28963 19211 28977
rect 18861 28946 19051 28956
rect 19177 28919 19211 28963
rect 18633 28841 18667 28885
rect 18701 28911 19125 28912
rect 18701 28909 18871 28911
rect 18701 28875 18717 28909
rect 18751 28875 18785 28909
rect 18819 28877 18871 28909
rect 18905 28909 19125 28911
rect 18905 28877 19075 28909
rect 18819 28875 19075 28877
rect 19109 28875 19125 28909
rect 19177 28841 19211 28885
rect 18633 28827 18767 28841
rect 18667 28825 18767 28827
rect 18667 28793 18733 28825
rect 18633 28791 18733 28793
rect 18633 28775 18767 28791
rect 18801 28832 18930 28840
rect 18801 28798 18803 28832
rect 18837 28806 18930 28832
rect 18964 28806 19067 28840
rect 18837 28798 19067 28806
rect 18801 28794 19067 28798
rect 18633 28735 18667 28775
rect 18801 28741 18835 28794
rect 18701 28707 18717 28741
rect 18751 28707 18785 28741
rect 18819 28707 18835 28741
rect 18869 28738 18999 28760
rect 18633 28672 18667 28701
rect 18869 28704 18944 28738
rect 18980 28704 18999 28738
rect 19033 28741 19067 28794
rect 19101 28827 19211 28841
rect 19101 28825 19177 28827
rect 19135 28793 19177 28825
rect 19135 28791 19211 28793
rect 19101 28775 19211 28791
rect 19033 28707 19075 28741
rect 19109 28707 19125 28741
rect 19177 28735 19211 28775
rect 18869 28690 18999 28704
rect 19177 28672 19211 28701
rect 18625 28309 18659 28326
rect 19169 28309 19203 28326
rect 18625 28297 18892 28309
rect 18659 28263 18730 28297
rect 18764 28263 18823 28297
rect 18857 28263 18892 28297
rect 18625 28251 18892 28263
rect 19024 28297 19203 28309
rect 19024 28263 19041 28297
rect 19075 28263 19169 28297
rect 19024 28251 19203 28263
rect 18625 28205 18659 28251
rect 18625 28115 18659 28171
rect 18693 28200 19135 28216
rect 18693 28199 18832 28200
rect 18866 28199 19135 28200
rect 18693 28165 18701 28199
rect 18735 28165 18772 28199
rect 18806 28166 18832 28199
rect 18877 28169 19055 28199
rect 18806 28165 18843 28166
rect 18877 28165 18890 28169
rect 19004 28165 19055 28169
rect 19089 28165 19135 28199
rect 19169 28205 19203 28251
rect 18693 28149 18890 28165
rect 18625 28113 18701 28115
rect 18659 28081 18701 28113
rect 18735 28081 18769 28115
rect 18803 28081 18837 28115
rect 18871 28081 18887 28115
rect 18659 28079 18887 28081
rect 18625 28072 18887 28079
rect 18921 28101 18937 28135
rect 18971 28101 18987 28135
rect 19169 28131 19203 28171
rect 18625 28021 18659 28072
rect 18921 28034 18987 28101
rect 19077 28115 19203 28131
rect 19077 28081 19093 28115
rect 19127 28113 19203 28115
rect 19127 28081 19169 28113
rect 19077 28079 19169 28081
rect 19077 28067 19203 28079
rect 18625 27929 18659 27987
rect 18697 28020 18987 28034
rect 19169 28021 19203 28067
rect 18697 28018 19067 28020
rect 18697 27984 18701 28018
rect 18735 27984 18769 28018
rect 18803 27986 19067 28018
rect 19101 27986 19117 28020
rect 18803 27984 19117 27986
rect 18697 27980 19117 27984
rect 18697 27968 18843 27980
rect 19063 27970 19117 27980
rect 18871 27932 19038 27946
rect 18871 27930 19125 27932
rect 18625 27837 18659 27895
rect 18702 27920 19125 27930
rect 18702 27916 19054 27920
rect 19088 27916 19125 27920
rect 18702 27914 19022 27916
rect 18702 27880 18707 27914
rect 18741 27880 18775 27914
rect 18809 27880 18843 27914
rect 18877 27908 19022 27914
rect 18877 27899 18897 27908
rect 18877 27880 18887 27899
rect 19013 27897 19022 27908
rect 18702 27864 18887 27880
rect 19021 27882 19022 27897
rect 19088 27886 19090 27916
rect 19056 27882 19090 27886
rect 19124 27882 19125 27916
rect 18921 27840 18937 27874
rect 18971 27840 18987 27874
rect 19021 27866 19125 27882
rect 19169 27929 19203 27987
rect 18659 27803 18731 27830
rect 18625 27796 18731 27803
rect 18765 27796 18811 27830
rect 18845 27796 18861 27830
rect 18625 27745 18659 27796
rect 18921 27764 18987 27840
rect 19169 27837 19203 27895
rect 19047 27798 19063 27832
rect 19097 27803 19169 27832
rect 19097 27798 19203 27803
rect 18921 27762 19126 27764
rect 18625 27653 18659 27711
rect 18693 27748 19126 27762
rect 18693 27744 19024 27748
rect 18693 27710 18701 27744
rect 18735 27710 18772 27744
rect 18806 27710 18843 27744
rect 18877 27724 19024 27744
rect 18877 27710 18880 27724
rect 18693 27694 18880 27710
rect 19021 27714 19024 27724
rect 19058 27714 19092 27748
rect 19021 27698 19126 27714
rect 19169 27745 19203 27798
rect 18659 27620 18759 27647
rect 18659 27619 18709 27620
rect 18625 27586 18709 27619
rect 18743 27586 18759 27620
rect 18625 27584 18759 27586
rect 18805 27616 18880 27694
rect 18625 27561 18659 27584
rect 18805 27582 18821 27616
rect 18855 27582 18880 27616
rect 18921 27656 18937 27690
rect 18971 27656 18987 27690
rect 18921 27548 18987 27656
rect 19169 27653 19203 27711
rect 19063 27642 19169 27645
rect 19063 27608 19079 27642
rect 19113 27619 19169 27642
rect 19113 27608 19203 27619
rect 19063 27603 19203 27608
rect 19169 27561 19203 27603
rect 18625 27469 18659 27527
rect 18625 27377 18659 27435
rect 18719 27514 19113 27548
rect 18719 27421 18753 27514
rect 18787 27446 18821 27480
rect 18855 27467 19045 27480
rect 18855 27446 18863 27467
rect 18787 27433 18863 27446
rect 18897 27433 19045 27467
rect 18787 27421 19045 27433
rect 18787 27416 18995 27421
rect 18979 27387 18995 27416
rect 19029 27387 19045 27421
rect 19079 27444 19113 27514
rect 19079 27391 19113 27410
rect 19169 27469 19203 27527
rect 18719 27371 18753 27387
rect 18793 27380 18937 27382
rect 18793 27346 18795 27380
rect 18829 27378 18937 27380
rect 18829 27346 18887 27378
rect 18793 27344 18887 27346
rect 18921 27344 18937 27378
rect 19169 27377 19203 27435
rect 18625 27285 18659 27343
rect 19079 27341 19113 27357
rect 18693 27292 18709 27326
rect 18743 27310 18759 27326
rect 18743 27307 19079 27310
rect 18743 27292 19113 27307
rect 18693 27276 19113 27292
rect 19169 27285 19203 27343
rect 18625 27242 18659 27251
rect 18625 27208 18701 27242
rect 18735 27208 18769 27242
rect 18803 27208 18819 27242
rect 18871 27208 18887 27242
rect 18921 27208 18937 27242
rect 18625 27193 18659 27208
rect 18871 27174 18923 27208
rect 18973 27184 19033 27276
rect 19169 27240 19203 27251
rect 18625 27101 18659 27159
rect 18625 27009 18659 27067
rect 18625 26917 18659 26975
rect 18714 27140 18923 27174
rect 18967 27178 19033 27184
rect 18967 27144 18983 27178
rect 19017 27144 19033 27178
rect 19069 27222 19203 27240
rect 19069 27188 19085 27222
rect 19119 27193 19203 27222
rect 19119 27188 19169 27193
rect 19069 27166 19169 27188
rect 18714 27003 18748 27140
rect 18782 27068 18855 27106
rect 18889 27102 18923 27140
rect 18889 27068 19113 27102
rect 18782 27066 18821 27068
rect 18782 27032 18795 27066
rect 18829 27032 19039 27034
rect 18782 27000 19039 27032
rect 18714 26953 18748 26969
rect 18995 26979 19039 27000
rect 18842 26963 18961 26966
rect 18842 26929 18863 26963
rect 18897 26959 18961 26963
rect 18897 26929 18899 26959
rect 18842 26925 18899 26929
rect 18933 26925 18961 26959
rect 19029 26945 19039 26979
rect 19079 27023 19113 27068
rect 19079 26967 19113 26989
rect 19169 27101 19203 27159
rect 19169 27009 19203 27067
rect 18995 26929 19039 26945
rect 18842 26918 18961 26925
rect 19079 26912 19113 26928
rect 18625 26827 18659 26883
rect 18693 26877 18709 26911
rect 18743 26884 18804 26911
rect 19025 26884 19079 26895
rect 18743 26878 19079 26884
rect 18743 26877 19113 26878
rect 18693 26861 19113 26877
rect 19169 26917 19203 26975
rect 18778 26850 19051 26861
rect 19169 26827 19203 26883
rect 18625 26825 18701 26827
rect 18659 26793 18701 26825
rect 18735 26793 18751 26827
rect 18659 26791 18751 26793
rect 18625 26774 18751 26791
rect 18853 26782 18869 26816
rect 18903 26810 19043 26816
rect 18903 26782 18984 26810
rect 18625 26733 18659 26774
rect 18853 26770 18984 26782
rect 19024 26770 19043 26810
rect 19077 26793 19093 26827
rect 19127 26825 19203 26827
rect 19127 26793 19169 26825
rect 19077 26791 19169 26793
rect 19077 26777 19203 26791
rect 18853 26760 19043 26770
rect 19169 26733 19203 26777
rect 18625 26655 18659 26699
rect 18693 26725 19117 26726
rect 18693 26723 18863 26725
rect 18693 26689 18709 26723
rect 18743 26689 18777 26723
rect 18811 26691 18863 26723
rect 18897 26723 19117 26725
rect 18897 26691 19067 26723
rect 18811 26689 19067 26691
rect 19101 26689 19117 26723
rect 19169 26655 19203 26699
rect 18625 26641 18759 26655
rect 18659 26639 18759 26641
rect 18659 26607 18725 26639
rect 18625 26605 18725 26607
rect 18625 26589 18759 26605
rect 18793 26646 18922 26654
rect 18793 26612 18795 26646
rect 18829 26620 18922 26646
rect 18956 26620 19059 26654
rect 18829 26612 19059 26620
rect 18793 26608 19059 26612
rect 18625 26549 18659 26589
rect 18793 26555 18827 26608
rect 18693 26521 18709 26555
rect 18743 26521 18777 26555
rect 18811 26521 18827 26555
rect 18861 26552 18991 26574
rect 18625 26486 18659 26515
rect 18861 26518 18936 26552
rect 18972 26518 18991 26552
rect 19025 26555 19059 26608
rect 19093 26641 19203 26655
rect 19093 26639 19169 26641
rect 19127 26607 19169 26639
rect 19127 26605 19203 26607
rect 19093 26589 19203 26605
rect 19025 26521 19067 26555
rect 19101 26521 19117 26555
rect 19169 26549 19203 26589
rect 18861 26504 18991 26518
rect 19169 26486 19203 26515
rect 18629 26063 18663 26080
rect 19173 26063 19207 26080
rect 18629 26051 18896 26063
rect 18663 26017 18734 26051
rect 18768 26017 18827 26051
rect 18861 26017 18896 26051
rect 18629 26005 18896 26017
rect 19028 26051 19207 26063
rect 19028 26017 19045 26051
rect 19079 26017 19173 26051
rect 19028 26005 19207 26017
rect 18629 25959 18663 26005
rect 18629 25869 18663 25925
rect 18697 25954 19139 25970
rect 18697 25953 18836 25954
rect 18870 25953 19139 25954
rect 18697 25919 18705 25953
rect 18739 25919 18776 25953
rect 18810 25920 18836 25953
rect 18881 25923 19059 25953
rect 18810 25919 18847 25920
rect 18881 25919 18894 25923
rect 19008 25919 19059 25923
rect 19093 25919 19139 25953
rect 19173 25959 19207 26005
rect 18697 25903 18894 25919
rect 18629 25867 18705 25869
rect 18663 25835 18705 25867
rect 18739 25835 18773 25869
rect 18807 25835 18841 25869
rect 18875 25835 18891 25869
rect 18663 25833 18891 25835
rect 18629 25826 18891 25833
rect 18925 25855 18941 25889
rect 18975 25855 18991 25889
rect 19173 25885 19207 25925
rect 18629 25775 18663 25826
rect 18925 25788 18991 25855
rect 19081 25869 19207 25885
rect 19081 25835 19097 25869
rect 19131 25867 19207 25869
rect 19131 25835 19173 25867
rect 19081 25833 19173 25835
rect 19081 25821 19207 25833
rect 18629 25683 18663 25741
rect 18701 25774 18991 25788
rect 19173 25775 19207 25821
rect 18701 25772 19071 25774
rect 18701 25738 18705 25772
rect 18739 25738 18773 25772
rect 18807 25740 19071 25772
rect 19105 25740 19121 25774
rect 18807 25738 19121 25740
rect 18701 25734 19121 25738
rect 18701 25722 18847 25734
rect 19067 25724 19121 25734
rect 18875 25686 19042 25700
rect 18875 25684 19129 25686
rect 18629 25591 18663 25649
rect 18706 25674 19129 25684
rect 18706 25670 19058 25674
rect 19092 25670 19129 25674
rect 18706 25668 19026 25670
rect 18706 25634 18711 25668
rect 18745 25634 18779 25668
rect 18813 25634 18847 25668
rect 18881 25662 19026 25668
rect 18881 25653 18901 25662
rect 18881 25634 18891 25653
rect 19017 25651 19026 25662
rect 18706 25618 18891 25634
rect 19025 25636 19026 25651
rect 19092 25640 19094 25670
rect 19060 25636 19094 25640
rect 19128 25636 19129 25670
rect 18925 25594 18941 25628
rect 18975 25594 18991 25628
rect 19025 25620 19129 25636
rect 19173 25683 19207 25741
rect 18663 25557 18735 25584
rect 18629 25550 18735 25557
rect 18769 25550 18815 25584
rect 18849 25550 18865 25584
rect 18629 25499 18663 25550
rect 18925 25518 18991 25594
rect 19173 25591 19207 25649
rect 19051 25552 19067 25586
rect 19101 25557 19173 25586
rect 19101 25552 19207 25557
rect 18925 25516 19130 25518
rect 18629 25407 18663 25465
rect 18697 25502 19130 25516
rect 18697 25498 19028 25502
rect 18697 25464 18705 25498
rect 18739 25464 18776 25498
rect 18810 25464 18847 25498
rect 18881 25478 19028 25498
rect 18881 25464 18884 25478
rect 18697 25448 18884 25464
rect 19025 25468 19028 25478
rect 19062 25468 19096 25502
rect 19025 25452 19130 25468
rect 19173 25499 19207 25552
rect 18663 25374 18763 25401
rect 18663 25373 18713 25374
rect 18629 25340 18713 25373
rect 18747 25340 18763 25374
rect 18629 25338 18763 25340
rect 18809 25370 18884 25448
rect 18629 25315 18663 25338
rect 18809 25336 18825 25370
rect 18859 25336 18884 25370
rect 18925 25410 18941 25444
rect 18975 25410 18991 25444
rect 18925 25302 18991 25410
rect 19173 25407 19207 25465
rect 19067 25396 19173 25399
rect 19067 25362 19083 25396
rect 19117 25373 19173 25396
rect 19117 25362 19207 25373
rect 19067 25357 19207 25362
rect 19173 25315 19207 25357
rect 18629 25223 18663 25281
rect 18629 25131 18663 25189
rect 18723 25268 19117 25302
rect 18723 25175 18757 25268
rect 18791 25200 18825 25234
rect 18859 25221 19049 25234
rect 18859 25200 18867 25221
rect 18791 25187 18867 25200
rect 18901 25187 19049 25221
rect 18791 25175 19049 25187
rect 18791 25170 18999 25175
rect 18983 25141 18999 25170
rect 19033 25141 19049 25175
rect 19083 25198 19117 25268
rect 19083 25145 19117 25164
rect 19173 25223 19207 25281
rect 18723 25125 18757 25141
rect 18797 25134 18941 25136
rect 18797 25100 18799 25134
rect 18833 25132 18941 25134
rect 18833 25100 18891 25132
rect 18797 25098 18891 25100
rect 18925 25098 18941 25132
rect 19173 25131 19207 25189
rect 18629 25039 18663 25097
rect 19083 25095 19117 25111
rect 18697 25046 18713 25080
rect 18747 25064 18763 25080
rect 18747 25061 19083 25064
rect 18747 25046 19117 25061
rect 18697 25030 19117 25046
rect 19173 25039 19207 25097
rect 18629 24996 18663 25005
rect 18629 24962 18705 24996
rect 18739 24962 18773 24996
rect 18807 24962 18823 24996
rect 18875 24962 18891 24996
rect 18925 24962 18941 24996
rect 18629 24947 18663 24962
rect 18875 24928 18927 24962
rect 18977 24938 19037 25030
rect 19173 24994 19207 25005
rect 18629 24855 18663 24913
rect 18629 24763 18663 24821
rect 18629 24671 18663 24729
rect 18718 24894 18927 24928
rect 18971 24932 19037 24938
rect 18971 24898 18987 24932
rect 19021 24898 19037 24932
rect 19073 24976 19207 24994
rect 19073 24942 19089 24976
rect 19123 24947 19207 24976
rect 19123 24942 19173 24947
rect 19073 24920 19173 24942
rect 18718 24757 18752 24894
rect 18786 24822 18859 24860
rect 18893 24856 18927 24894
rect 18893 24822 19117 24856
rect 18786 24820 18825 24822
rect 18786 24786 18799 24820
rect 18833 24786 19043 24788
rect 18786 24754 19043 24786
rect 18718 24707 18752 24723
rect 18999 24733 19043 24754
rect 18846 24717 18965 24720
rect 18846 24683 18867 24717
rect 18901 24713 18965 24717
rect 18901 24683 18903 24713
rect 18846 24679 18903 24683
rect 18937 24679 18965 24713
rect 19033 24699 19043 24733
rect 19083 24777 19117 24822
rect 19083 24721 19117 24743
rect 19173 24855 19207 24913
rect 19173 24763 19207 24821
rect 18999 24683 19043 24699
rect 18846 24672 18965 24679
rect 19083 24666 19117 24682
rect 18629 24581 18663 24637
rect 18697 24631 18713 24665
rect 18747 24638 18808 24665
rect 19029 24638 19083 24649
rect 18747 24632 19083 24638
rect 18747 24631 19117 24632
rect 18697 24615 19117 24631
rect 19173 24671 19207 24729
rect 18782 24604 19055 24615
rect 19173 24581 19207 24637
rect 18629 24579 18705 24581
rect 18663 24547 18705 24579
rect 18739 24547 18755 24581
rect 18663 24545 18755 24547
rect 18629 24528 18755 24545
rect 18857 24536 18873 24570
rect 18907 24564 19047 24570
rect 18907 24536 18988 24564
rect 18629 24487 18663 24528
rect 18857 24524 18988 24536
rect 19028 24524 19047 24564
rect 19081 24547 19097 24581
rect 19131 24579 19207 24581
rect 19131 24547 19173 24579
rect 19081 24545 19173 24547
rect 19081 24531 19207 24545
rect 18857 24514 19047 24524
rect 19173 24487 19207 24531
rect 18629 24409 18663 24453
rect 18697 24479 19121 24480
rect 18697 24477 18867 24479
rect 18697 24443 18713 24477
rect 18747 24443 18781 24477
rect 18815 24445 18867 24477
rect 18901 24477 19121 24479
rect 18901 24445 19071 24477
rect 18815 24443 19071 24445
rect 19105 24443 19121 24477
rect 19173 24409 19207 24453
rect 18629 24395 18763 24409
rect 18663 24393 18763 24395
rect 18663 24361 18729 24393
rect 18629 24359 18729 24361
rect 18629 24343 18763 24359
rect 18797 24400 18926 24408
rect 18797 24366 18799 24400
rect 18833 24374 18926 24400
rect 18960 24374 19063 24408
rect 18833 24366 19063 24374
rect 18797 24362 19063 24366
rect 18629 24303 18663 24343
rect 18797 24309 18831 24362
rect 18697 24275 18713 24309
rect 18747 24275 18781 24309
rect 18815 24275 18831 24309
rect 18865 24306 18995 24328
rect 18629 24240 18663 24269
rect 18865 24272 18940 24306
rect 18976 24272 18995 24306
rect 19029 24309 19063 24362
rect 19097 24395 19207 24409
rect 19097 24393 19173 24395
rect 19131 24361 19173 24393
rect 19131 24359 19207 24361
rect 19097 24343 19207 24359
rect 19029 24275 19071 24309
rect 19105 24275 19121 24309
rect 19173 24303 19207 24343
rect 18865 24258 18995 24272
rect 19173 24240 19207 24269
rect 7670 23355 7699 23389
rect 7733 23355 7791 23389
rect 7825 23355 7883 23389
rect 7917 23355 7975 23389
rect 8009 23355 8067 23389
rect 8101 23355 8159 23389
rect 8193 23355 8251 23389
rect 8285 23355 8343 23389
rect 8377 23355 8435 23389
rect 8469 23355 8527 23389
rect 8561 23355 8619 23389
rect 8653 23355 8711 23389
rect 8745 23355 8803 23389
rect 8837 23355 8895 23389
rect 8929 23355 8987 23389
rect 9021 23355 9079 23389
rect 9113 23355 9171 23389
rect 9205 23355 9263 23389
rect 9297 23355 9355 23389
rect 9389 23355 9447 23389
rect 9481 23355 9510 23389
rect 9916 23359 9945 23393
rect 9979 23359 10037 23393
rect 10071 23359 10129 23393
rect 10163 23359 10221 23393
rect 10255 23359 10313 23393
rect 10347 23359 10405 23393
rect 10439 23359 10497 23393
rect 10531 23359 10589 23393
rect 10623 23359 10681 23393
rect 10715 23359 10773 23393
rect 10807 23359 10865 23393
rect 10899 23359 10957 23393
rect 10991 23359 11049 23393
rect 11083 23359 11141 23393
rect 11175 23359 11233 23393
rect 11267 23359 11325 23393
rect 11359 23359 11417 23393
rect 11451 23359 11509 23393
rect 11543 23359 11601 23393
rect 11635 23359 11693 23393
rect 11727 23359 11756 23393
rect 7705 23305 7739 23321
rect 7705 23237 7739 23271
rect 7773 23289 7839 23355
rect 7773 23255 7789 23289
rect 7823 23255 7839 23289
rect 7873 23305 7910 23321
rect 7907 23271 7910 23305
rect 7873 23237 7910 23271
rect 7958 23313 8011 23355
rect 7958 23279 7977 23313
rect 7958 23263 8011 23279
rect 8045 23305 8095 23321
rect 8045 23271 8061 23305
rect 8392 23313 8426 23355
rect 7739 23219 7838 23221
rect 7739 23203 7796 23219
rect 7705 23187 7796 23203
rect 7792 23185 7796 23187
rect 7830 23185 7838 23219
rect 7688 23078 7758 23153
rect 7688 23042 7702 23078
rect 7736 23042 7758 23078
rect 7688 23023 7758 23042
rect 7792 23092 7838 23185
rect 7792 23058 7804 23092
rect 7792 22989 7838 23058
rect 7705 22955 7838 22989
rect 7907 23203 7910 23237
rect 8045 23236 8095 23271
rect 8137 23266 8153 23300
rect 8187 23266 8358 23300
rect 7873 23151 7910 23203
rect 8034 23210 8095 23236
rect 8184 23219 8290 23232
rect 7873 23117 7875 23151
rect 7909 23117 7910 23151
rect 7705 22947 7739 22955
rect 7873 22947 7910 23117
rect 7944 23145 8000 23161
rect 7944 23111 7966 23145
rect 7944 23030 8000 23111
rect 7944 22990 7954 23030
rect 7994 22990 8000 23030
rect 7944 22971 8000 22990
rect 8034 22989 8068 23210
rect 8184 23185 8216 23219
rect 8250 23193 8290 23219
rect 8102 23151 8150 23172
rect 8102 23117 8113 23151
rect 8147 23117 8150 23151
rect 8102 23115 8150 23117
rect 8102 23081 8109 23115
rect 8143 23081 8150 23115
rect 8102 23053 8150 23081
rect 8184 23019 8218 23185
rect 8252 23159 8290 23193
rect 8324 23143 8358 23266
rect 8392 23245 8426 23279
rect 8392 23195 8426 23211
rect 8460 23305 8510 23321
rect 8460 23271 8476 23305
rect 8768 23305 8831 23355
rect 8460 23255 8510 23271
rect 8555 23261 8571 23295
rect 8605 23261 8732 23295
rect 8324 23127 8426 23143
rect 8324 23125 8392 23127
rect 8034 22963 8079 22989
rect 8113 22985 8129 23019
rect 8163 22985 8218 23019
rect 8113 22975 8218 22985
rect 8252 23093 8392 23125
rect 8252 23091 8426 23093
rect 7705 22897 7739 22913
rect 7773 22887 7789 22921
rect 7823 22887 7839 22921
rect 7907 22913 7910 22947
rect 7873 22897 7910 22913
rect 7961 22921 8011 22937
rect 7773 22845 7839 22887
rect 7961 22887 7977 22921
rect 8045 22935 8079 22963
rect 8252 22935 8286 23091
rect 8392 23077 8426 23091
rect 8328 23041 8368 23047
rect 8460 23041 8494 23255
rect 8528 23219 8566 23221
rect 8528 23185 8530 23219
rect 8564 23185 8566 23219
rect 8528 23127 8566 23185
rect 8562 23093 8566 23127
rect 8528 23077 8566 23093
rect 8600 23193 8664 23227
rect 8600 23159 8630 23193
rect 8600 23151 8664 23159
rect 8600 23117 8617 23151
rect 8651 23117 8664 23151
rect 8328 23031 8494 23041
rect 8600 23035 8664 23117
rect 8362 22997 8494 23031
rect 8328 22981 8494 22997
rect 8045 22901 8062 22935
rect 8096 22901 8112 22935
rect 8151 22901 8173 22935
rect 8207 22901 8286 22935
rect 8350 22929 8424 22945
rect 7961 22845 8011 22887
rect 8350 22895 8372 22929
rect 8406 22895 8424 22929
rect 8460 22935 8494 22981
rect 8571 23019 8664 23035
rect 8605 22985 8664 23019
rect 8571 22969 8664 22985
rect 8698 23093 8732 23261
rect 8768 23271 8770 23305
rect 8804 23271 8831 23305
rect 8768 23255 8831 23271
rect 8878 23313 8946 23321
rect 8878 23279 8894 23313
rect 8928 23279 8946 23313
rect 8878 23242 8946 23279
rect 8878 23209 8894 23242
rect 8766 23208 8894 23209
rect 8928 23208 8946 23242
rect 8766 23193 8946 23208
rect 8800 23171 8946 23193
rect 8800 23159 8894 23171
rect 8766 23137 8894 23159
rect 8928 23137 8946 23171
rect 8980 23283 9014 23355
rect 9152 23313 9218 23317
rect 8980 23203 9014 23249
rect 8980 23153 9014 23169
rect 9048 23307 9114 23312
rect 9048 23273 9064 23307
rect 9098 23273 9114 23307
rect 9048 23239 9114 23273
rect 9048 23205 9064 23239
rect 9098 23205 9114 23239
rect 9048 23171 9114 23205
rect 9152 23279 9168 23313
rect 9202 23279 9218 23313
rect 9152 23245 9218 23279
rect 9152 23211 9168 23245
rect 9202 23211 9218 23245
rect 9152 23171 9218 23211
rect 8766 23134 8946 23137
rect 8908 23093 8946 23134
rect 9048 23137 9064 23171
rect 9098 23143 9114 23171
rect 9098 23137 9130 23143
rect 9048 23127 9130 23137
rect 9083 23117 9130 23127
rect 8698 23077 8874 23093
rect 8698 23043 8840 23077
rect 8698 23027 8874 23043
rect 8908 23077 9058 23093
rect 8908 23043 9024 23077
rect 8908 23027 9058 23043
rect 8698 22935 8732 23027
rect 8908 22993 8948 23027
rect 9092 23001 9130 23117
rect 9081 22993 9130 23001
rect 8882 22990 8948 22993
rect 8882 22956 8898 22990
rect 8932 22956 8948 22990
rect 9050 22992 9130 22993
rect 8460 22901 8491 22935
rect 8525 22901 8541 22935
rect 8575 22901 8594 22935
rect 8628 22901 8732 22935
rect 8787 22935 8829 22951
rect 8787 22901 8792 22935
rect 8826 22901 8829 22935
rect 8350 22845 8424 22895
rect 8787 22845 8829 22901
rect 8882 22922 8948 22956
rect 8882 22888 8898 22922
rect 8932 22888 8948 22922
rect 8982 22951 9016 22967
rect 8982 22845 9016 22917
rect 9050 22958 9066 22992
rect 9100 22976 9130 22992
rect 9164 23093 9218 23171
rect 9256 23313 9299 23355
rect 9256 23279 9265 23313
rect 9256 23245 9299 23279
rect 9256 23211 9265 23245
rect 9256 23177 9299 23211
rect 9256 23143 9265 23177
rect 9256 23127 9299 23143
rect 9333 23313 9400 23321
rect 9333 23279 9349 23313
rect 9383 23279 9400 23313
rect 9333 23242 9400 23279
rect 9333 23208 9349 23242
rect 9383 23208 9400 23242
rect 9333 23182 9400 23208
rect 9333 23171 9350 23182
rect 9333 23137 9349 23171
rect 9384 23148 9400 23182
rect 9383 23137 9400 23148
rect 9333 23124 9400 23137
rect 9164 23077 9319 23093
rect 9164 23043 9285 23077
rect 9164 23027 9319 23043
rect 9100 22960 9116 22976
rect 9050 22926 9070 22958
rect 9104 22926 9116 22960
rect 9164 22951 9204 23027
rect 9353 23010 9400 23124
rect 9435 23284 9493 23355
rect 9435 23250 9447 23284
rect 9481 23250 9493 23284
rect 9435 23191 9493 23250
rect 9951 23309 9985 23325
rect 9951 23241 9985 23275
rect 10019 23293 10085 23359
rect 10019 23259 10035 23293
rect 10069 23259 10085 23293
rect 10119 23309 10156 23325
rect 10153 23275 10156 23309
rect 10119 23241 10156 23275
rect 10204 23317 10257 23359
rect 10204 23283 10223 23317
rect 10204 23267 10257 23283
rect 10291 23309 10341 23325
rect 10291 23275 10307 23309
rect 10638 23317 10672 23359
rect 9985 23223 10084 23225
rect 9985 23207 10042 23223
rect 9951 23191 10042 23207
rect 9435 23157 9447 23191
rect 9481 23157 9493 23191
rect 10038 23189 10042 23191
rect 10076 23189 10084 23223
rect 9435 23122 9493 23157
rect 9934 23082 10004 23157
rect 9934 23046 9948 23082
rect 9982 23046 10004 23082
rect 9934 23027 10004 23046
rect 10038 23096 10084 23189
rect 10038 23062 10050 23096
rect 9050 22924 9116 22926
rect 9050 22890 9066 22924
rect 9100 22890 9116 22924
rect 9154 22947 9204 22951
rect 9154 22913 9170 22947
rect 9349 22959 9400 23010
rect 10038 22993 10084 23062
rect 9154 22897 9204 22913
rect 9251 22921 9315 22937
rect 9050 22889 9116 22890
rect 9251 22887 9265 22921
rect 9299 22887 9315 22921
rect 9251 22845 9315 22887
rect 9383 22925 9400 22959
rect 9349 22879 9400 22925
rect 9435 22973 9493 22990
rect 9435 22939 9447 22973
rect 9481 22939 9493 22973
rect 9435 22845 9493 22939
rect 9951 22959 10084 22993
rect 10153 23207 10156 23241
rect 10291 23240 10341 23275
rect 10383 23270 10399 23304
rect 10433 23270 10604 23304
rect 10119 23155 10156 23207
rect 10280 23214 10341 23240
rect 10430 23223 10536 23236
rect 10119 23121 10121 23155
rect 10155 23121 10156 23155
rect 9951 22951 9985 22959
rect 10119 22951 10156 23121
rect 10190 23149 10246 23165
rect 10190 23115 10212 23149
rect 10190 23034 10246 23115
rect 10190 22994 10200 23034
rect 10240 22994 10246 23034
rect 10190 22975 10246 22994
rect 10280 22993 10314 23214
rect 10430 23189 10462 23223
rect 10496 23197 10536 23223
rect 10348 23155 10396 23176
rect 10348 23121 10359 23155
rect 10393 23121 10396 23155
rect 10348 23119 10396 23121
rect 10348 23085 10355 23119
rect 10389 23085 10396 23119
rect 10348 23057 10396 23085
rect 10430 23023 10464 23189
rect 10498 23163 10536 23197
rect 10570 23147 10604 23270
rect 10638 23249 10672 23283
rect 10638 23199 10672 23215
rect 10706 23309 10756 23325
rect 10706 23275 10722 23309
rect 11014 23309 11077 23359
rect 10706 23259 10756 23275
rect 10801 23265 10817 23299
rect 10851 23265 10978 23299
rect 10570 23131 10672 23147
rect 10570 23129 10638 23131
rect 10280 22967 10325 22993
rect 10359 22989 10375 23023
rect 10409 22989 10464 23023
rect 10359 22979 10464 22989
rect 10498 23097 10638 23129
rect 10498 23095 10672 23097
rect 9951 22901 9985 22917
rect 10019 22891 10035 22925
rect 10069 22891 10085 22925
rect 10153 22917 10156 22951
rect 10119 22901 10156 22917
rect 10207 22925 10257 22941
rect 10019 22849 10085 22891
rect 10207 22891 10223 22925
rect 10291 22939 10325 22967
rect 10498 22939 10532 23095
rect 10638 23081 10672 23095
rect 10574 23045 10614 23051
rect 10706 23045 10740 23259
rect 10774 23223 10812 23225
rect 10774 23189 10776 23223
rect 10810 23189 10812 23223
rect 10774 23131 10812 23189
rect 10808 23097 10812 23131
rect 10774 23081 10812 23097
rect 10846 23197 10910 23231
rect 10846 23163 10876 23197
rect 10846 23155 10910 23163
rect 10846 23121 10863 23155
rect 10897 23121 10910 23155
rect 10574 23035 10740 23045
rect 10846 23039 10910 23121
rect 10608 23001 10740 23035
rect 10574 22985 10740 23001
rect 10291 22905 10308 22939
rect 10342 22905 10358 22939
rect 10397 22905 10419 22939
rect 10453 22905 10532 22939
rect 10596 22933 10670 22949
rect 10207 22849 10257 22891
rect 10596 22899 10618 22933
rect 10652 22899 10670 22933
rect 10706 22939 10740 22985
rect 10817 23023 10910 23039
rect 10851 22989 10910 23023
rect 10817 22973 10910 22989
rect 10944 23097 10978 23265
rect 11014 23275 11016 23309
rect 11050 23275 11077 23309
rect 11014 23259 11077 23275
rect 11124 23317 11192 23325
rect 11124 23283 11140 23317
rect 11174 23283 11192 23317
rect 11124 23246 11192 23283
rect 11124 23213 11140 23246
rect 11012 23212 11140 23213
rect 11174 23212 11192 23246
rect 11012 23197 11192 23212
rect 11046 23175 11192 23197
rect 11046 23163 11140 23175
rect 11012 23141 11140 23163
rect 11174 23141 11192 23175
rect 11226 23287 11260 23359
rect 11398 23317 11464 23321
rect 11226 23207 11260 23253
rect 11226 23157 11260 23173
rect 11294 23311 11360 23316
rect 11294 23277 11310 23311
rect 11344 23277 11360 23311
rect 11294 23243 11360 23277
rect 11294 23209 11310 23243
rect 11344 23209 11360 23243
rect 11294 23175 11360 23209
rect 11398 23283 11414 23317
rect 11448 23283 11464 23317
rect 11398 23249 11464 23283
rect 11398 23215 11414 23249
rect 11448 23215 11464 23249
rect 11398 23175 11464 23215
rect 11012 23138 11192 23141
rect 11154 23097 11192 23138
rect 11294 23141 11310 23175
rect 11344 23147 11360 23175
rect 11344 23141 11376 23147
rect 11294 23131 11376 23141
rect 11329 23121 11376 23131
rect 10944 23081 11120 23097
rect 10944 23047 11086 23081
rect 10944 23031 11120 23047
rect 11154 23081 11304 23097
rect 11154 23047 11270 23081
rect 11154 23031 11304 23047
rect 10944 22939 10978 23031
rect 11154 22997 11194 23031
rect 11338 23005 11376 23121
rect 11327 22997 11376 23005
rect 11128 22994 11194 22997
rect 11128 22960 11144 22994
rect 11178 22960 11194 22994
rect 11296 22996 11376 22997
rect 10706 22905 10737 22939
rect 10771 22905 10787 22939
rect 10821 22905 10840 22939
rect 10874 22905 10978 22939
rect 11033 22939 11075 22955
rect 11033 22905 11038 22939
rect 11072 22905 11075 22939
rect 10596 22849 10670 22899
rect 11033 22849 11075 22905
rect 11128 22926 11194 22960
rect 11128 22892 11144 22926
rect 11178 22892 11194 22926
rect 11228 22955 11262 22971
rect 11228 22849 11262 22921
rect 11296 22962 11312 22996
rect 11346 22980 11376 22996
rect 11410 23097 11464 23175
rect 11502 23317 11545 23359
rect 11502 23283 11511 23317
rect 11502 23249 11545 23283
rect 11502 23215 11511 23249
rect 11502 23181 11545 23215
rect 11502 23147 11511 23181
rect 11502 23131 11545 23147
rect 11579 23317 11646 23325
rect 11579 23283 11595 23317
rect 11629 23283 11646 23317
rect 11579 23246 11646 23283
rect 11579 23212 11595 23246
rect 11629 23212 11646 23246
rect 11579 23186 11646 23212
rect 11579 23175 11596 23186
rect 11579 23141 11595 23175
rect 11630 23152 11646 23186
rect 11629 23141 11646 23152
rect 11579 23128 11646 23141
rect 11410 23081 11565 23097
rect 11410 23047 11531 23081
rect 11410 23031 11565 23047
rect 11346 22964 11362 22980
rect 11296 22930 11316 22962
rect 11350 22930 11362 22964
rect 11410 22955 11450 23031
rect 11599 23014 11646 23128
rect 11681 23288 11739 23359
rect 12102 23351 12131 23385
rect 12165 23351 12223 23385
rect 12257 23351 12315 23385
rect 12349 23351 12407 23385
rect 12441 23351 12499 23385
rect 12533 23351 12591 23385
rect 12625 23351 12683 23385
rect 12717 23351 12775 23385
rect 12809 23351 12867 23385
rect 12901 23351 12959 23385
rect 12993 23351 13051 23385
rect 13085 23351 13143 23385
rect 13177 23351 13235 23385
rect 13269 23351 13327 23385
rect 13361 23351 13419 23385
rect 13453 23351 13511 23385
rect 13545 23351 13603 23385
rect 13637 23351 13695 23385
rect 13729 23351 13787 23385
rect 13821 23351 13879 23385
rect 13913 23351 13942 23385
rect 14348 23355 14377 23389
rect 14411 23355 14469 23389
rect 14503 23355 14561 23389
rect 14595 23355 14653 23389
rect 14687 23355 14745 23389
rect 14779 23355 14837 23389
rect 14871 23355 14929 23389
rect 14963 23355 15021 23389
rect 15055 23355 15113 23389
rect 15147 23355 15205 23389
rect 15239 23355 15297 23389
rect 15331 23355 15389 23389
rect 15423 23355 15481 23389
rect 15515 23355 15573 23389
rect 15607 23355 15665 23389
rect 15699 23355 15757 23389
rect 15791 23355 15849 23389
rect 15883 23355 15941 23389
rect 15975 23355 16033 23389
rect 16067 23355 16125 23389
rect 16159 23355 16188 23389
rect 16630 23355 16659 23389
rect 16693 23355 16751 23389
rect 16785 23355 16843 23389
rect 16877 23355 16935 23389
rect 16969 23355 17027 23389
rect 17061 23355 17119 23389
rect 17153 23355 17211 23389
rect 17245 23355 17303 23389
rect 17337 23355 17395 23389
rect 17429 23355 17487 23389
rect 17521 23355 17579 23389
rect 17613 23355 17671 23389
rect 17705 23355 17763 23389
rect 17797 23355 17855 23389
rect 17889 23355 17947 23389
rect 17981 23355 18039 23389
rect 18073 23355 18131 23389
rect 18165 23355 18223 23389
rect 18257 23355 18315 23389
rect 18349 23355 18407 23389
rect 18441 23355 18470 23389
rect 11681 23254 11693 23288
rect 11727 23254 11739 23288
rect 11681 23195 11739 23254
rect 11681 23161 11693 23195
rect 11727 23161 11739 23195
rect 12137 23301 12171 23317
rect 12137 23233 12171 23267
rect 12205 23285 12271 23351
rect 12205 23251 12221 23285
rect 12255 23251 12271 23285
rect 12305 23301 12342 23317
rect 12339 23267 12342 23301
rect 12305 23233 12342 23267
rect 12390 23309 12443 23351
rect 12390 23275 12409 23309
rect 12390 23259 12443 23275
rect 12477 23301 12527 23317
rect 12477 23267 12493 23301
rect 12824 23309 12858 23351
rect 12171 23215 12270 23217
rect 12171 23199 12228 23215
rect 12137 23183 12228 23199
rect 11681 23126 11739 23161
rect 12224 23181 12228 23183
rect 12262 23181 12270 23215
rect 12120 23074 12190 23149
rect 12120 23038 12134 23074
rect 12168 23038 12190 23074
rect 12120 23019 12190 23038
rect 12224 23088 12270 23181
rect 12224 23054 12236 23088
rect 11296 22928 11362 22930
rect 11296 22894 11312 22928
rect 11346 22894 11362 22928
rect 11400 22951 11450 22955
rect 11400 22917 11416 22951
rect 11595 22963 11646 23014
rect 11400 22901 11450 22917
rect 11497 22925 11561 22941
rect 11296 22893 11362 22894
rect 11497 22891 11511 22925
rect 11545 22891 11561 22925
rect 11497 22849 11561 22891
rect 11629 22929 11646 22963
rect 11595 22883 11646 22929
rect 11681 22977 11739 22994
rect 12224 22985 12270 23054
rect 11681 22943 11693 22977
rect 11727 22943 11739 22977
rect 11681 22849 11739 22943
rect 12137 22951 12270 22985
rect 12339 23199 12342 23233
rect 12477 23232 12527 23267
rect 12569 23262 12585 23296
rect 12619 23262 12790 23296
rect 12305 23147 12342 23199
rect 12466 23206 12527 23232
rect 12616 23215 12722 23228
rect 12305 23113 12307 23147
rect 12341 23113 12342 23147
rect 12137 22943 12171 22951
rect 12305 22943 12342 23113
rect 12376 23141 12432 23157
rect 12376 23107 12398 23141
rect 12376 23026 12432 23107
rect 12376 22986 12386 23026
rect 12426 22986 12432 23026
rect 12376 22967 12432 22986
rect 12466 22985 12500 23206
rect 12616 23181 12648 23215
rect 12682 23189 12722 23215
rect 12534 23147 12582 23168
rect 12534 23113 12545 23147
rect 12579 23113 12582 23147
rect 12534 23111 12582 23113
rect 12534 23077 12541 23111
rect 12575 23077 12582 23111
rect 12534 23049 12582 23077
rect 12616 23015 12650 23181
rect 12684 23155 12722 23189
rect 12756 23139 12790 23262
rect 12824 23241 12858 23275
rect 12824 23191 12858 23207
rect 12892 23301 12942 23317
rect 12892 23267 12908 23301
rect 13200 23301 13263 23351
rect 12892 23251 12942 23267
rect 12987 23257 13003 23291
rect 13037 23257 13164 23291
rect 12756 23123 12858 23139
rect 12756 23121 12824 23123
rect 12466 22959 12511 22985
rect 12545 22981 12561 23015
rect 12595 22981 12650 23015
rect 12545 22971 12650 22981
rect 12684 23089 12824 23121
rect 12684 23087 12858 23089
rect 12137 22893 12171 22909
rect 12205 22883 12221 22917
rect 12255 22883 12271 22917
rect 12339 22909 12342 22943
rect 12305 22893 12342 22909
rect 12393 22917 12443 22933
rect 7670 22811 7699 22845
rect 7733 22811 7791 22845
rect 7825 22811 7883 22845
rect 7917 22811 7975 22845
rect 8009 22811 8067 22845
rect 8101 22811 8159 22845
rect 8193 22811 8251 22845
rect 8285 22811 8343 22845
rect 8377 22811 8435 22845
rect 8469 22811 8527 22845
rect 8561 22811 8619 22845
rect 8653 22811 8711 22845
rect 8745 22811 8803 22845
rect 8837 22811 8895 22845
rect 8929 22811 8987 22845
rect 9021 22811 9079 22845
rect 9113 22811 9171 22845
rect 9205 22811 9263 22845
rect 9297 22811 9355 22845
rect 9389 22811 9447 22845
rect 9481 22811 9510 22845
rect 9916 22815 9945 22849
rect 9979 22815 10037 22849
rect 10071 22815 10129 22849
rect 10163 22815 10221 22849
rect 10255 22815 10313 22849
rect 10347 22815 10405 22849
rect 10439 22815 10497 22849
rect 10531 22815 10589 22849
rect 10623 22815 10681 22849
rect 10715 22815 10773 22849
rect 10807 22815 10865 22849
rect 10899 22815 10957 22849
rect 10991 22815 11049 22849
rect 11083 22815 11141 22849
rect 11175 22815 11233 22849
rect 11267 22815 11325 22849
rect 11359 22815 11417 22849
rect 11451 22815 11509 22849
rect 11543 22815 11601 22849
rect 11635 22815 11693 22849
rect 11727 22815 11756 22849
rect 12205 22841 12271 22883
rect 12393 22883 12409 22917
rect 12477 22931 12511 22959
rect 12684 22931 12718 23087
rect 12824 23073 12858 23087
rect 12760 23037 12800 23043
rect 12892 23037 12926 23251
rect 12960 23215 12998 23217
rect 12960 23181 12962 23215
rect 12996 23181 12998 23215
rect 12960 23123 12998 23181
rect 12994 23089 12998 23123
rect 12960 23073 12998 23089
rect 13032 23189 13096 23223
rect 13032 23155 13062 23189
rect 13032 23147 13096 23155
rect 13032 23113 13049 23147
rect 13083 23113 13096 23147
rect 12760 23027 12926 23037
rect 13032 23031 13096 23113
rect 12794 22993 12926 23027
rect 12760 22977 12926 22993
rect 12477 22897 12494 22931
rect 12528 22897 12544 22931
rect 12583 22897 12605 22931
rect 12639 22897 12718 22931
rect 12782 22925 12856 22941
rect 12393 22841 12443 22883
rect 12782 22891 12804 22925
rect 12838 22891 12856 22925
rect 12892 22931 12926 22977
rect 13003 23015 13096 23031
rect 13037 22981 13096 23015
rect 13003 22965 13096 22981
rect 13130 23089 13164 23257
rect 13200 23267 13202 23301
rect 13236 23267 13263 23301
rect 13200 23251 13263 23267
rect 13310 23309 13378 23317
rect 13310 23275 13326 23309
rect 13360 23275 13378 23309
rect 13310 23238 13378 23275
rect 13310 23205 13326 23238
rect 13198 23204 13326 23205
rect 13360 23204 13378 23238
rect 13198 23189 13378 23204
rect 13232 23167 13378 23189
rect 13232 23155 13326 23167
rect 13198 23133 13326 23155
rect 13360 23133 13378 23167
rect 13412 23279 13446 23351
rect 13584 23309 13650 23313
rect 13412 23199 13446 23245
rect 13412 23149 13446 23165
rect 13480 23303 13546 23308
rect 13480 23269 13496 23303
rect 13530 23269 13546 23303
rect 13480 23235 13546 23269
rect 13480 23201 13496 23235
rect 13530 23201 13546 23235
rect 13480 23167 13546 23201
rect 13584 23275 13600 23309
rect 13634 23275 13650 23309
rect 13584 23241 13650 23275
rect 13584 23207 13600 23241
rect 13634 23207 13650 23241
rect 13584 23167 13650 23207
rect 13198 23130 13378 23133
rect 13340 23089 13378 23130
rect 13480 23133 13496 23167
rect 13530 23139 13546 23167
rect 13530 23133 13562 23139
rect 13480 23123 13562 23133
rect 13515 23113 13562 23123
rect 13130 23073 13306 23089
rect 13130 23039 13272 23073
rect 13130 23023 13306 23039
rect 13340 23073 13490 23089
rect 13340 23039 13456 23073
rect 13340 23023 13490 23039
rect 13130 22931 13164 23023
rect 13340 22989 13380 23023
rect 13524 22997 13562 23113
rect 13513 22989 13562 22997
rect 13314 22986 13380 22989
rect 13314 22952 13330 22986
rect 13364 22952 13380 22986
rect 13482 22988 13562 22989
rect 12892 22897 12923 22931
rect 12957 22897 12973 22931
rect 13007 22897 13026 22931
rect 13060 22897 13164 22931
rect 13219 22931 13261 22947
rect 13219 22897 13224 22931
rect 13258 22897 13261 22931
rect 12782 22841 12856 22891
rect 13219 22841 13261 22897
rect 13314 22918 13380 22952
rect 13314 22884 13330 22918
rect 13364 22884 13380 22918
rect 13414 22947 13448 22963
rect 13414 22841 13448 22913
rect 13482 22954 13498 22988
rect 13532 22972 13562 22988
rect 13596 23089 13650 23167
rect 13688 23309 13731 23351
rect 13688 23275 13697 23309
rect 13688 23241 13731 23275
rect 13688 23207 13697 23241
rect 13688 23173 13731 23207
rect 13688 23139 13697 23173
rect 13688 23123 13731 23139
rect 13765 23309 13832 23317
rect 13765 23275 13781 23309
rect 13815 23275 13832 23309
rect 13765 23238 13832 23275
rect 13765 23204 13781 23238
rect 13815 23204 13832 23238
rect 13765 23178 13832 23204
rect 13765 23167 13782 23178
rect 13765 23133 13781 23167
rect 13816 23144 13832 23178
rect 13815 23133 13832 23144
rect 13765 23120 13832 23133
rect 13596 23073 13751 23089
rect 13596 23039 13717 23073
rect 13596 23023 13751 23039
rect 13532 22956 13548 22972
rect 13482 22922 13502 22954
rect 13536 22922 13548 22956
rect 13596 22947 13636 23023
rect 13785 23006 13832 23120
rect 13867 23280 13925 23351
rect 13867 23246 13879 23280
rect 13913 23246 13925 23280
rect 13867 23187 13925 23246
rect 14383 23305 14417 23321
rect 14383 23237 14417 23271
rect 14451 23289 14517 23355
rect 14451 23255 14467 23289
rect 14501 23255 14517 23289
rect 14551 23305 14588 23321
rect 14585 23271 14588 23305
rect 14551 23237 14588 23271
rect 14636 23313 14689 23355
rect 14636 23279 14655 23313
rect 14636 23263 14689 23279
rect 14723 23305 14773 23321
rect 14723 23271 14739 23305
rect 15070 23313 15104 23355
rect 14417 23219 14516 23221
rect 14417 23203 14474 23219
rect 14383 23187 14474 23203
rect 13867 23153 13879 23187
rect 13913 23153 13925 23187
rect 14470 23185 14474 23187
rect 14508 23185 14516 23219
rect 13867 23118 13925 23153
rect 14366 23078 14436 23153
rect 14366 23042 14380 23078
rect 14414 23042 14436 23078
rect 14366 23023 14436 23042
rect 14470 23092 14516 23185
rect 14470 23058 14482 23092
rect 13482 22920 13548 22922
rect 13482 22886 13498 22920
rect 13532 22886 13548 22920
rect 13586 22943 13636 22947
rect 13586 22909 13602 22943
rect 13781 22955 13832 23006
rect 14470 22989 14516 23058
rect 13586 22893 13636 22909
rect 13683 22917 13747 22933
rect 13482 22885 13548 22886
rect 13683 22883 13697 22917
rect 13731 22883 13747 22917
rect 13683 22841 13747 22883
rect 13815 22921 13832 22955
rect 13781 22875 13832 22921
rect 13867 22969 13925 22986
rect 13867 22935 13879 22969
rect 13913 22935 13925 22969
rect 13867 22841 13925 22935
rect 14383 22955 14516 22989
rect 14585 23203 14588 23237
rect 14723 23236 14773 23271
rect 14815 23266 14831 23300
rect 14865 23266 15036 23300
rect 14551 23151 14588 23203
rect 14712 23210 14773 23236
rect 14862 23219 14968 23232
rect 14551 23117 14553 23151
rect 14587 23117 14588 23151
rect 14383 22947 14417 22955
rect 14551 22947 14588 23117
rect 14622 23145 14678 23161
rect 14622 23111 14644 23145
rect 14622 23030 14678 23111
rect 14622 22990 14632 23030
rect 14672 22990 14678 23030
rect 14622 22971 14678 22990
rect 14712 22989 14746 23210
rect 14862 23185 14894 23219
rect 14928 23193 14968 23219
rect 14780 23151 14828 23172
rect 14780 23117 14791 23151
rect 14825 23117 14828 23151
rect 14780 23115 14828 23117
rect 14780 23081 14787 23115
rect 14821 23081 14828 23115
rect 14780 23053 14828 23081
rect 14862 23019 14896 23185
rect 14930 23159 14968 23193
rect 15002 23143 15036 23266
rect 15070 23245 15104 23279
rect 15070 23195 15104 23211
rect 15138 23305 15188 23321
rect 15138 23271 15154 23305
rect 15446 23305 15509 23355
rect 15138 23255 15188 23271
rect 15233 23261 15249 23295
rect 15283 23261 15410 23295
rect 15002 23127 15104 23143
rect 15002 23125 15070 23127
rect 14712 22963 14757 22989
rect 14791 22985 14807 23019
rect 14841 22985 14896 23019
rect 14791 22975 14896 22985
rect 14930 23093 15070 23125
rect 14930 23091 15104 23093
rect 14383 22897 14417 22913
rect 14451 22887 14467 22921
rect 14501 22887 14517 22921
rect 14585 22913 14588 22947
rect 14551 22897 14588 22913
rect 14639 22921 14689 22937
rect 14451 22845 14517 22887
rect 14639 22887 14655 22921
rect 14723 22935 14757 22963
rect 14930 22935 14964 23091
rect 15070 23077 15104 23091
rect 15006 23041 15046 23047
rect 15138 23041 15172 23255
rect 15206 23219 15244 23221
rect 15206 23185 15208 23219
rect 15242 23185 15244 23219
rect 15206 23127 15244 23185
rect 15240 23093 15244 23127
rect 15206 23077 15244 23093
rect 15278 23193 15342 23227
rect 15278 23159 15308 23193
rect 15278 23151 15342 23159
rect 15278 23117 15295 23151
rect 15329 23117 15342 23151
rect 15006 23031 15172 23041
rect 15278 23035 15342 23117
rect 15040 22997 15172 23031
rect 15006 22981 15172 22997
rect 14723 22901 14740 22935
rect 14774 22901 14790 22935
rect 14829 22901 14851 22935
rect 14885 22901 14964 22935
rect 15028 22929 15102 22945
rect 14639 22845 14689 22887
rect 15028 22895 15050 22929
rect 15084 22895 15102 22929
rect 15138 22935 15172 22981
rect 15249 23019 15342 23035
rect 15283 22985 15342 23019
rect 15249 22969 15342 22985
rect 15376 23093 15410 23261
rect 15446 23271 15448 23305
rect 15482 23271 15509 23305
rect 15446 23255 15509 23271
rect 15556 23313 15624 23321
rect 15556 23279 15572 23313
rect 15606 23279 15624 23313
rect 15556 23242 15624 23279
rect 15556 23209 15572 23242
rect 15444 23208 15572 23209
rect 15606 23208 15624 23242
rect 15444 23193 15624 23208
rect 15478 23171 15624 23193
rect 15478 23159 15572 23171
rect 15444 23137 15572 23159
rect 15606 23137 15624 23171
rect 15658 23283 15692 23355
rect 15830 23313 15896 23317
rect 15658 23203 15692 23249
rect 15658 23153 15692 23169
rect 15726 23307 15792 23312
rect 15726 23273 15742 23307
rect 15776 23273 15792 23307
rect 15726 23239 15792 23273
rect 15726 23205 15742 23239
rect 15776 23205 15792 23239
rect 15726 23171 15792 23205
rect 15830 23279 15846 23313
rect 15880 23279 15896 23313
rect 15830 23245 15896 23279
rect 15830 23211 15846 23245
rect 15880 23211 15896 23245
rect 15830 23171 15896 23211
rect 15444 23134 15624 23137
rect 15586 23093 15624 23134
rect 15726 23137 15742 23171
rect 15776 23143 15792 23171
rect 15776 23137 15808 23143
rect 15726 23127 15808 23137
rect 15761 23117 15808 23127
rect 15376 23077 15552 23093
rect 15376 23043 15518 23077
rect 15376 23027 15552 23043
rect 15586 23077 15736 23093
rect 15586 23043 15702 23077
rect 15586 23027 15736 23043
rect 15376 22935 15410 23027
rect 15586 22993 15626 23027
rect 15770 23001 15808 23117
rect 15759 22993 15808 23001
rect 15560 22990 15626 22993
rect 15560 22956 15576 22990
rect 15610 22956 15626 22990
rect 15728 22992 15808 22993
rect 15138 22901 15169 22935
rect 15203 22901 15219 22935
rect 15253 22901 15272 22935
rect 15306 22901 15410 22935
rect 15465 22935 15507 22951
rect 15465 22901 15470 22935
rect 15504 22901 15507 22935
rect 15028 22845 15102 22895
rect 15465 22845 15507 22901
rect 15560 22922 15626 22956
rect 15560 22888 15576 22922
rect 15610 22888 15626 22922
rect 15660 22951 15694 22967
rect 15660 22845 15694 22917
rect 15728 22958 15744 22992
rect 15778 22976 15808 22992
rect 15842 23093 15896 23171
rect 15934 23313 15977 23355
rect 15934 23279 15943 23313
rect 15934 23245 15977 23279
rect 15934 23211 15943 23245
rect 15934 23177 15977 23211
rect 15934 23143 15943 23177
rect 15934 23127 15977 23143
rect 16011 23313 16078 23321
rect 16011 23279 16027 23313
rect 16061 23279 16078 23313
rect 16011 23242 16078 23279
rect 16011 23208 16027 23242
rect 16061 23208 16078 23242
rect 16011 23182 16078 23208
rect 16011 23171 16028 23182
rect 16011 23137 16027 23171
rect 16062 23148 16078 23182
rect 16061 23137 16078 23148
rect 16011 23124 16078 23137
rect 15842 23077 15997 23093
rect 15842 23043 15963 23077
rect 15842 23027 15997 23043
rect 15778 22960 15794 22976
rect 15728 22926 15748 22958
rect 15782 22926 15794 22960
rect 15842 22951 15882 23027
rect 16031 23010 16078 23124
rect 16113 23284 16171 23355
rect 16113 23250 16125 23284
rect 16159 23250 16171 23284
rect 16113 23191 16171 23250
rect 16113 23157 16125 23191
rect 16159 23157 16171 23191
rect 16665 23305 16699 23321
rect 16665 23237 16699 23271
rect 16733 23289 16799 23355
rect 16733 23255 16749 23289
rect 16783 23255 16799 23289
rect 16833 23305 16870 23321
rect 16867 23271 16870 23305
rect 16833 23237 16870 23271
rect 16918 23313 16971 23355
rect 16918 23279 16937 23313
rect 16918 23263 16971 23279
rect 17005 23305 17055 23321
rect 17005 23271 17021 23305
rect 17352 23313 17386 23355
rect 16699 23219 16798 23221
rect 16699 23203 16756 23219
rect 16665 23187 16756 23203
rect 16113 23122 16171 23157
rect 16752 23185 16756 23187
rect 16790 23185 16798 23219
rect 16648 23078 16718 23153
rect 16648 23042 16662 23078
rect 16696 23042 16718 23078
rect 16648 23023 16718 23042
rect 16752 23092 16798 23185
rect 16752 23058 16764 23092
rect 15728 22924 15794 22926
rect 15728 22890 15744 22924
rect 15778 22890 15794 22924
rect 15832 22947 15882 22951
rect 15832 22913 15848 22947
rect 16027 22959 16078 23010
rect 15832 22897 15882 22913
rect 15929 22921 15993 22937
rect 15728 22889 15794 22890
rect 15929 22887 15943 22921
rect 15977 22887 15993 22921
rect 15929 22845 15993 22887
rect 16061 22925 16078 22959
rect 16027 22879 16078 22925
rect 16113 22973 16171 22990
rect 16752 22989 16798 23058
rect 16113 22939 16125 22973
rect 16159 22939 16171 22973
rect 16113 22845 16171 22939
rect 16665 22955 16798 22989
rect 16867 23203 16870 23237
rect 17005 23236 17055 23271
rect 17097 23266 17113 23300
rect 17147 23266 17318 23300
rect 16833 23151 16870 23203
rect 16994 23210 17055 23236
rect 17144 23219 17250 23232
rect 16833 23117 16835 23151
rect 16869 23117 16870 23151
rect 16665 22947 16699 22955
rect 16833 22947 16870 23117
rect 16904 23145 16960 23161
rect 16904 23111 16926 23145
rect 16904 23030 16960 23111
rect 16904 22990 16914 23030
rect 16954 22990 16960 23030
rect 16904 22971 16960 22990
rect 16994 22989 17028 23210
rect 17144 23185 17176 23219
rect 17210 23193 17250 23219
rect 17062 23151 17110 23172
rect 17062 23117 17073 23151
rect 17107 23117 17110 23151
rect 17062 23115 17110 23117
rect 17062 23081 17069 23115
rect 17103 23081 17110 23115
rect 17062 23053 17110 23081
rect 17144 23019 17178 23185
rect 17212 23159 17250 23193
rect 17284 23143 17318 23266
rect 17352 23245 17386 23279
rect 17352 23195 17386 23211
rect 17420 23305 17470 23321
rect 17420 23271 17436 23305
rect 17728 23305 17791 23355
rect 17420 23255 17470 23271
rect 17515 23261 17531 23295
rect 17565 23261 17692 23295
rect 17284 23127 17386 23143
rect 17284 23125 17352 23127
rect 16994 22963 17039 22989
rect 17073 22985 17089 23019
rect 17123 22985 17178 23019
rect 17073 22975 17178 22985
rect 17212 23093 17352 23125
rect 17212 23091 17386 23093
rect 16665 22897 16699 22913
rect 16733 22887 16749 22921
rect 16783 22887 16799 22921
rect 16867 22913 16870 22947
rect 16833 22897 16870 22913
rect 16921 22921 16971 22937
rect 16733 22845 16799 22887
rect 16921 22887 16937 22921
rect 17005 22935 17039 22963
rect 17212 22935 17246 23091
rect 17352 23077 17386 23091
rect 17288 23041 17328 23047
rect 17420 23041 17454 23255
rect 17488 23219 17526 23221
rect 17488 23185 17490 23219
rect 17524 23185 17526 23219
rect 17488 23127 17526 23185
rect 17522 23093 17526 23127
rect 17488 23077 17526 23093
rect 17560 23193 17624 23227
rect 17560 23159 17590 23193
rect 17560 23151 17624 23159
rect 17560 23117 17577 23151
rect 17611 23117 17624 23151
rect 17288 23031 17454 23041
rect 17560 23035 17624 23117
rect 17322 22997 17454 23031
rect 17288 22981 17454 22997
rect 17005 22901 17022 22935
rect 17056 22901 17072 22935
rect 17111 22901 17133 22935
rect 17167 22901 17246 22935
rect 17310 22929 17384 22945
rect 16921 22845 16971 22887
rect 17310 22895 17332 22929
rect 17366 22895 17384 22929
rect 17420 22935 17454 22981
rect 17531 23019 17624 23035
rect 17565 22985 17624 23019
rect 17531 22969 17624 22985
rect 17658 23093 17692 23261
rect 17728 23271 17730 23305
rect 17764 23271 17791 23305
rect 17728 23255 17791 23271
rect 17838 23313 17906 23321
rect 17838 23279 17854 23313
rect 17888 23279 17906 23313
rect 17838 23242 17906 23279
rect 17838 23209 17854 23242
rect 17726 23208 17854 23209
rect 17888 23208 17906 23242
rect 17726 23193 17906 23208
rect 17760 23171 17906 23193
rect 17760 23159 17854 23171
rect 17726 23137 17854 23159
rect 17888 23137 17906 23171
rect 17940 23283 17974 23355
rect 18112 23313 18178 23317
rect 17940 23203 17974 23249
rect 17940 23153 17974 23169
rect 18008 23307 18074 23312
rect 18008 23273 18024 23307
rect 18058 23273 18074 23307
rect 18008 23239 18074 23273
rect 18008 23205 18024 23239
rect 18058 23205 18074 23239
rect 18008 23171 18074 23205
rect 18112 23279 18128 23313
rect 18162 23279 18178 23313
rect 18112 23245 18178 23279
rect 18112 23211 18128 23245
rect 18162 23211 18178 23245
rect 18112 23171 18178 23211
rect 17726 23134 17906 23137
rect 17868 23093 17906 23134
rect 18008 23137 18024 23171
rect 18058 23143 18074 23171
rect 18058 23137 18090 23143
rect 18008 23127 18090 23137
rect 18043 23117 18090 23127
rect 17658 23077 17834 23093
rect 17658 23043 17800 23077
rect 17658 23027 17834 23043
rect 17868 23077 18018 23093
rect 17868 23043 17984 23077
rect 17868 23027 18018 23043
rect 17658 22935 17692 23027
rect 17868 22993 17908 23027
rect 18052 23001 18090 23117
rect 18041 22993 18090 23001
rect 17842 22990 17908 22993
rect 17842 22956 17858 22990
rect 17892 22956 17908 22990
rect 18010 22992 18090 22993
rect 17420 22901 17451 22935
rect 17485 22901 17501 22935
rect 17535 22901 17554 22935
rect 17588 22901 17692 22935
rect 17747 22935 17789 22951
rect 17747 22901 17752 22935
rect 17786 22901 17789 22935
rect 17310 22845 17384 22895
rect 17747 22845 17789 22901
rect 17842 22922 17908 22956
rect 17842 22888 17858 22922
rect 17892 22888 17908 22922
rect 17942 22951 17976 22967
rect 17942 22845 17976 22917
rect 18010 22958 18026 22992
rect 18060 22976 18090 22992
rect 18124 23093 18178 23171
rect 18216 23313 18259 23355
rect 18216 23279 18225 23313
rect 18216 23245 18259 23279
rect 18216 23211 18225 23245
rect 18216 23177 18259 23211
rect 18216 23143 18225 23177
rect 18216 23127 18259 23143
rect 18293 23313 18360 23321
rect 18293 23279 18309 23313
rect 18343 23279 18360 23313
rect 18293 23242 18360 23279
rect 18293 23208 18309 23242
rect 18343 23208 18360 23242
rect 18293 23182 18360 23208
rect 18293 23171 18310 23182
rect 18293 23137 18309 23171
rect 18344 23148 18360 23182
rect 18343 23137 18360 23148
rect 18293 23124 18360 23137
rect 18124 23077 18279 23093
rect 18124 23043 18245 23077
rect 18124 23027 18279 23043
rect 18060 22960 18076 22976
rect 18010 22926 18030 22958
rect 18064 22926 18076 22960
rect 18124 22951 18164 23027
rect 18313 23010 18360 23124
rect 18395 23284 18453 23355
rect 18395 23250 18407 23284
rect 18441 23250 18453 23284
rect 18395 23191 18453 23250
rect 18395 23157 18407 23191
rect 18441 23157 18453 23191
rect 18395 23122 18453 23157
rect 18010 22924 18076 22926
rect 18010 22890 18026 22924
rect 18060 22890 18076 22924
rect 18114 22947 18164 22951
rect 18114 22913 18130 22947
rect 18309 22959 18360 23010
rect 18114 22897 18164 22913
rect 18211 22921 18275 22937
rect 18010 22889 18076 22890
rect 18211 22887 18225 22921
rect 18259 22887 18275 22921
rect 18211 22845 18275 22887
rect 18343 22925 18360 22959
rect 18309 22879 18360 22925
rect 18395 22973 18453 22990
rect 18395 22939 18407 22973
rect 18441 22939 18453 22973
rect 18395 22845 18453 22939
rect 12102 22807 12131 22841
rect 12165 22807 12223 22841
rect 12257 22807 12315 22841
rect 12349 22807 12407 22841
rect 12441 22807 12499 22841
rect 12533 22807 12591 22841
rect 12625 22807 12683 22841
rect 12717 22807 12775 22841
rect 12809 22807 12867 22841
rect 12901 22807 12959 22841
rect 12993 22807 13051 22841
rect 13085 22807 13143 22841
rect 13177 22807 13235 22841
rect 13269 22807 13327 22841
rect 13361 22807 13419 22841
rect 13453 22807 13511 22841
rect 13545 22807 13603 22841
rect 13637 22807 13695 22841
rect 13729 22807 13787 22841
rect 13821 22807 13879 22841
rect 13913 22807 13942 22841
rect 14348 22811 14377 22845
rect 14411 22811 14469 22845
rect 14503 22811 14561 22845
rect 14595 22811 14653 22845
rect 14687 22811 14745 22845
rect 14779 22811 14837 22845
rect 14871 22811 14929 22845
rect 14963 22811 15021 22845
rect 15055 22811 15113 22845
rect 15147 22811 15205 22845
rect 15239 22811 15297 22845
rect 15331 22811 15389 22845
rect 15423 22811 15481 22845
rect 15515 22811 15573 22845
rect 15607 22811 15665 22845
rect 15699 22811 15757 22845
rect 15791 22811 15849 22845
rect 15883 22811 15941 22845
rect 15975 22811 16033 22845
rect 16067 22811 16125 22845
rect 16159 22811 16188 22845
rect 16630 22811 16659 22845
rect 16693 22811 16751 22845
rect 16785 22811 16843 22845
rect 16877 22811 16935 22845
rect 16969 22811 17027 22845
rect 17061 22811 17119 22845
rect 17153 22811 17211 22845
rect 17245 22811 17303 22845
rect 17337 22811 17395 22845
rect 17429 22811 17487 22845
rect 17521 22811 17579 22845
rect 17613 22811 17671 22845
rect 17705 22811 17763 22845
rect 17797 22811 17855 22845
rect 17889 22811 17947 22845
rect 17981 22811 18039 22845
rect 18073 22811 18131 22845
rect 18165 22811 18223 22845
rect 18257 22811 18315 22845
rect 18349 22811 18407 22845
rect 18441 22811 18470 22845
rect 9430 17777 9459 17811
rect 9493 17777 9551 17811
rect 9585 17777 9643 17811
rect 9677 17777 9719 17811
rect 9753 17777 9782 17811
rect 9496 17731 9562 17743
rect 9496 17697 9512 17731
rect 9546 17697 9562 17731
rect 9496 17663 9562 17697
rect 9496 17629 9512 17663
rect 9546 17629 9562 17663
rect 9496 17617 9562 17629
rect 9596 17731 9642 17777
rect 9630 17697 9642 17731
rect 9596 17663 9642 17697
rect 9630 17629 9642 17663
rect 9707 17683 9765 17777
rect 9707 17649 9719 17683
rect 9753 17649 9765 17683
rect 16267 17667 16296 17701
rect 16330 17667 16374 17701
rect 16408 17667 16466 17701
rect 16500 17667 16558 17701
rect 16592 17667 16621 17701
rect 17133 17669 17162 17703
rect 17196 17669 17248 17703
rect 17282 17669 17340 17703
rect 17374 17669 17432 17703
rect 17466 17669 17495 17703
rect 9707 17632 9765 17649
rect 15481 17629 15510 17663
rect 15544 17629 15596 17663
rect 15630 17629 15688 17663
rect 15722 17629 15780 17663
rect 15814 17629 15843 17663
rect 9496 17568 9542 17617
rect 9596 17613 9642 17629
rect 9532 17532 9542 17568
rect 9496 17497 9542 17532
rect 9576 17545 9592 17579
rect 9626 17572 9642 17579
rect 9576 17536 9596 17545
rect 9632 17536 9642 17572
rect 9576 17531 9642 17536
rect 15498 17535 15556 17629
rect 15498 17501 15510 17535
rect 15544 17501 15556 17535
rect 9496 17479 9562 17497
rect 9496 17445 9512 17479
rect 9546 17445 9562 17479
rect 9496 17411 9562 17445
rect 9496 17377 9512 17411
rect 9546 17377 9562 17411
rect 9496 17343 9562 17377
rect 9496 17309 9512 17343
rect 9546 17309 9562 17343
rect 9496 17301 9562 17309
rect 9596 17479 9638 17495
rect 9630 17445 9638 17479
rect 9596 17411 9638 17445
rect 9630 17377 9638 17411
rect 9596 17343 9638 17377
rect 9630 17309 9638 17343
rect 9596 17267 9638 17309
rect 9707 17465 9765 17500
rect 15498 17484 15556 17501
rect 15633 17583 15699 17595
rect 15633 17549 15649 17583
rect 15683 17549 15699 17583
rect 15633 17515 15699 17549
rect 9707 17431 9719 17465
rect 9753 17431 9765 17465
rect 9707 17372 9765 17431
rect 9707 17338 9719 17372
rect 9753 17338 9765 17372
rect 15633 17481 15649 17515
rect 15683 17481 15699 17515
rect 15633 17469 15699 17481
rect 15733 17583 15779 17629
rect 15767 17549 15779 17583
rect 15733 17515 15779 17549
rect 16284 17573 16342 17667
rect 16284 17539 16296 17573
rect 16330 17539 16342 17573
rect 16284 17522 16342 17539
rect 16411 17621 16477 17633
rect 16411 17587 16427 17621
rect 16461 17587 16477 17621
rect 16411 17553 16477 17587
rect 15767 17481 15779 17515
rect 15633 17436 15679 17469
rect 15733 17465 15779 17481
rect 16411 17519 16427 17553
rect 16461 17519 16477 17553
rect 16411 17507 16477 17519
rect 16511 17621 16557 17667
rect 16545 17587 16557 17621
rect 16511 17553 16557 17587
rect 16545 17519 16557 17553
rect 17150 17575 17208 17669
rect 17150 17541 17162 17575
rect 17196 17541 17208 17575
rect 17150 17524 17208 17541
rect 17285 17623 17351 17635
rect 17285 17589 17301 17623
rect 17335 17589 17351 17623
rect 17285 17555 17351 17589
rect 16411 17468 16457 17507
rect 16511 17503 16557 17519
rect 17285 17521 17301 17555
rect 17335 17521 17351 17555
rect 17285 17509 17351 17521
rect 17385 17623 17431 17669
rect 17911 17659 17940 17693
rect 17974 17659 18016 17693
rect 18050 17659 18108 17693
rect 18142 17659 18200 17693
rect 18234 17659 18263 17693
rect 19027 17661 19056 17695
rect 19090 17661 19138 17695
rect 19172 17661 19230 17695
rect 19264 17661 19322 17695
rect 19356 17661 19385 17695
rect 19893 17663 19922 17697
rect 19956 17663 20012 17697
rect 20046 17663 20104 17697
rect 20138 17663 20196 17697
rect 20230 17663 20259 17697
rect 17419 17589 17431 17623
rect 17385 17555 17431 17589
rect 17419 17521 17431 17555
rect 17285 17476 17331 17509
rect 17385 17505 17431 17521
rect 17928 17565 17986 17659
rect 17928 17531 17940 17565
rect 17974 17531 17986 17565
rect 17928 17514 17986 17531
rect 18053 17613 18119 17625
rect 18053 17579 18069 17613
rect 18103 17579 18119 17613
rect 18053 17545 18119 17579
rect 18053 17511 18069 17545
rect 18103 17511 18119 17545
rect 15633 17402 15635 17436
rect 15669 17402 15679 17436
rect 16411 17434 16413 17468
rect 16449 17434 16457 17468
rect 9707 17267 9765 17338
rect 15498 17317 15556 17352
rect 15498 17283 15510 17317
rect 15544 17283 15556 17317
rect 9430 17233 9459 17267
rect 9493 17233 9551 17267
rect 9585 17233 9643 17267
rect 9677 17233 9719 17267
rect 9753 17233 9782 17267
rect 15498 17224 15556 17283
rect 15498 17190 15510 17224
rect 15544 17190 15556 17224
rect 15498 17119 15556 17190
rect 15633 17349 15679 17402
rect 15713 17428 15729 17431
rect 15713 17394 15725 17428
rect 15763 17394 15779 17431
rect 15713 17383 15779 17394
rect 16284 17355 16342 17390
rect 15633 17331 15699 17349
rect 15633 17297 15649 17331
rect 15683 17297 15699 17331
rect 15633 17263 15699 17297
rect 15633 17229 15649 17263
rect 15683 17229 15699 17263
rect 15633 17195 15699 17229
rect 15633 17161 15649 17195
rect 15683 17161 15699 17195
rect 15633 17153 15699 17161
rect 15733 17331 15775 17347
rect 15767 17297 15775 17331
rect 15733 17263 15775 17297
rect 15767 17229 15775 17263
rect 15733 17195 15775 17229
rect 15767 17161 15775 17195
rect 15733 17119 15775 17161
rect 16284 17321 16296 17355
rect 16330 17321 16342 17355
rect 16284 17262 16342 17321
rect 16284 17228 16296 17262
rect 16330 17228 16342 17262
rect 16284 17157 16342 17228
rect 16411 17387 16457 17434
rect 16491 17435 16507 17469
rect 16541 17464 16557 17469
rect 16491 17430 16517 17435
rect 16551 17430 16557 17464
rect 16491 17421 16557 17430
rect 17285 17442 17287 17476
rect 17321 17442 17331 17476
rect 18053 17499 18119 17511
rect 18153 17613 18199 17659
rect 18187 17579 18199 17613
rect 18153 17545 18199 17579
rect 18187 17511 18199 17545
rect 19044 17567 19102 17661
rect 19044 17533 19056 17567
rect 19090 17533 19102 17567
rect 19044 17516 19102 17533
rect 19175 17615 19241 17627
rect 19175 17581 19191 17615
rect 19225 17581 19241 17615
rect 19175 17547 19241 17581
rect 18053 17472 18099 17499
rect 18153 17495 18199 17511
rect 19175 17513 19191 17547
rect 19225 17513 19241 17547
rect 19175 17501 19241 17513
rect 19275 17615 19321 17661
rect 19309 17581 19321 17615
rect 19275 17547 19321 17581
rect 19309 17513 19321 17547
rect 19910 17569 19968 17663
rect 19910 17535 19922 17569
rect 19956 17535 19968 17569
rect 19910 17518 19968 17535
rect 20049 17617 20115 17629
rect 20049 17583 20065 17617
rect 20099 17583 20115 17617
rect 20049 17549 20115 17583
rect 16411 17369 16477 17387
rect 16411 17335 16427 17369
rect 16461 17335 16477 17369
rect 16411 17301 16477 17335
rect 16411 17267 16427 17301
rect 16461 17267 16477 17301
rect 16411 17233 16477 17267
rect 16411 17199 16427 17233
rect 16461 17199 16477 17233
rect 16411 17191 16477 17199
rect 16511 17369 16553 17385
rect 16545 17335 16553 17369
rect 16511 17301 16553 17335
rect 16545 17267 16553 17301
rect 16511 17233 16553 17267
rect 16545 17199 16553 17233
rect 16511 17157 16553 17199
rect 17150 17357 17208 17392
rect 17150 17323 17162 17357
rect 17196 17323 17208 17357
rect 17150 17264 17208 17323
rect 17150 17230 17162 17264
rect 17196 17230 17208 17264
rect 17150 17159 17208 17230
rect 17285 17389 17331 17442
rect 17365 17468 17381 17471
rect 17365 17434 17377 17468
rect 17415 17434 17431 17471
rect 17365 17423 17431 17434
rect 18053 17438 18059 17472
rect 18097 17438 18099 17472
rect 19175 17462 19221 17501
rect 19275 17497 19321 17513
rect 20049 17515 20065 17549
rect 20099 17515 20115 17549
rect 20049 17503 20115 17515
rect 20149 17617 20195 17663
rect 20663 17653 20692 17687
rect 20726 17653 20780 17687
rect 20814 17653 20872 17687
rect 20906 17653 20964 17687
rect 20998 17653 21027 17687
rect 20183 17583 20195 17617
rect 20149 17549 20195 17583
rect 20183 17515 20195 17549
rect 20049 17470 20095 17503
rect 20149 17499 20195 17515
rect 20680 17559 20738 17653
rect 20680 17525 20692 17559
rect 20726 17525 20738 17559
rect 20680 17508 20738 17525
rect 20817 17607 20883 17619
rect 20817 17573 20833 17607
rect 20867 17573 20883 17607
rect 20817 17539 20883 17573
rect 20817 17505 20833 17539
rect 20867 17505 20883 17539
rect 17285 17371 17351 17389
rect 17285 17337 17301 17371
rect 17335 17337 17351 17371
rect 17285 17303 17351 17337
rect 17285 17269 17301 17303
rect 17335 17269 17351 17303
rect 17285 17235 17351 17269
rect 17285 17201 17301 17235
rect 17335 17201 17351 17235
rect 17285 17193 17351 17201
rect 17385 17371 17427 17387
rect 17419 17337 17427 17371
rect 17385 17303 17427 17337
rect 17419 17269 17427 17303
rect 17385 17235 17427 17269
rect 17419 17201 17427 17235
rect 17385 17159 17427 17201
rect 17928 17347 17986 17382
rect 17928 17313 17940 17347
rect 17974 17313 17986 17347
rect 17928 17254 17986 17313
rect 17928 17220 17940 17254
rect 17974 17220 17986 17254
rect 16267 17123 16296 17157
rect 16330 17123 16374 17157
rect 16408 17123 16466 17157
rect 16500 17123 16558 17157
rect 16592 17123 16621 17157
rect 17133 17125 17162 17159
rect 17196 17125 17248 17159
rect 17282 17125 17340 17159
rect 17374 17125 17432 17159
rect 17466 17125 17495 17159
rect 17928 17149 17986 17220
rect 18053 17379 18099 17438
rect 18133 17460 18149 17461
rect 18133 17426 18147 17460
rect 18183 17426 18199 17461
rect 18133 17413 18199 17426
rect 19175 17428 19177 17462
rect 19213 17428 19221 17462
rect 18053 17361 18119 17379
rect 18053 17327 18069 17361
rect 18103 17327 18119 17361
rect 18053 17293 18119 17327
rect 18053 17259 18069 17293
rect 18103 17259 18119 17293
rect 18053 17225 18119 17259
rect 18053 17191 18069 17225
rect 18103 17191 18119 17225
rect 18053 17183 18119 17191
rect 18153 17361 18195 17377
rect 18187 17327 18195 17361
rect 18153 17293 18195 17327
rect 18187 17259 18195 17293
rect 18153 17225 18195 17259
rect 18187 17191 18195 17225
rect 18153 17149 18195 17191
rect 19044 17349 19102 17384
rect 19044 17315 19056 17349
rect 19090 17315 19102 17349
rect 19044 17256 19102 17315
rect 19044 17222 19056 17256
rect 19090 17222 19102 17256
rect 19044 17151 19102 17222
rect 19175 17381 19221 17428
rect 19255 17429 19271 17463
rect 19305 17458 19321 17463
rect 19255 17424 19281 17429
rect 19315 17424 19321 17458
rect 19255 17415 19321 17424
rect 20049 17436 20051 17470
rect 20085 17436 20095 17470
rect 20817 17493 20883 17505
rect 20917 17607 20963 17653
rect 21365 17651 21394 17685
rect 21428 17651 21486 17685
rect 21520 17651 21578 17685
rect 21612 17651 21670 17685
rect 21704 17651 21733 17685
rect 22149 17653 22178 17687
rect 22212 17653 22268 17687
rect 22302 17653 22360 17687
rect 22394 17653 22452 17687
rect 22486 17653 22515 17687
rect 20951 17573 20963 17607
rect 20917 17539 20963 17573
rect 20951 17505 20963 17539
rect 20817 17466 20863 17493
rect 20917 17489 20963 17505
rect 21431 17605 21497 17617
rect 21431 17571 21447 17605
rect 21481 17571 21497 17605
rect 21431 17537 21497 17571
rect 21431 17503 21447 17537
rect 21481 17503 21497 17537
rect 21431 17491 21497 17503
rect 21531 17605 21577 17651
rect 21565 17571 21577 17605
rect 21531 17537 21577 17571
rect 21565 17503 21577 17537
rect 21658 17557 21716 17651
rect 21658 17523 21670 17557
rect 21704 17523 21716 17557
rect 21658 17506 21716 17523
rect 22166 17559 22224 17653
rect 22166 17525 22178 17559
rect 22212 17525 22224 17559
rect 22166 17508 22224 17525
rect 22305 17607 22371 17619
rect 22305 17573 22321 17607
rect 22355 17573 22371 17607
rect 22305 17539 22371 17573
rect 19175 17363 19241 17381
rect 19175 17329 19191 17363
rect 19225 17329 19241 17363
rect 19175 17295 19241 17329
rect 19175 17261 19191 17295
rect 19225 17261 19241 17295
rect 19175 17227 19241 17261
rect 19175 17193 19191 17227
rect 19225 17193 19241 17227
rect 19175 17185 19241 17193
rect 19275 17363 19317 17379
rect 19309 17329 19317 17363
rect 19275 17295 19317 17329
rect 19309 17261 19317 17295
rect 19275 17227 19317 17261
rect 19309 17193 19317 17227
rect 19275 17151 19317 17193
rect 19910 17351 19968 17386
rect 19910 17317 19922 17351
rect 19956 17317 19968 17351
rect 19910 17258 19968 17317
rect 19910 17224 19922 17258
rect 19956 17224 19968 17258
rect 19910 17153 19968 17224
rect 20049 17383 20095 17436
rect 20129 17462 20145 17465
rect 20129 17428 20141 17462
rect 20179 17428 20195 17465
rect 20129 17417 20195 17428
rect 20817 17432 20823 17466
rect 20861 17432 20863 17466
rect 20049 17365 20115 17383
rect 20049 17331 20065 17365
rect 20099 17331 20115 17365
rect 20049 17297 20115 17331
rect 20049 17263 20065 17297
rect 20099 17263 20115 17297
rect 20049 17229 20115 17263
rect 20049 17195 20065 17229
rect 20099 17195 20115 17229
rect 20049 17187 20115 17195
rect 20149 17365 20191 17381
rect 20183 17331 20191 17365
rect 20149 17297 20191 17331
rect 20183 17263 20191 17297
rect 20149 17229 20191 17263
rect 20183 17195 20191 17229
rect 20149 17153 20191 17195
rect 20680 17341 20738 17376
rect 20680 17307 20692 17341
rect 20726 17307 20738 17341
rect 20680 17248 20738 17307
rect 20680 17214 20692 17248
rect 20726 17214 20738 17248
rect 15481 17085 15510 17119
rect 15544 17085 15596 17119
rect 15630 17085 15688 17119
rect 15722 17085 15780 17119
rect 15814 17085 15843 17119
rect 17911 17115 17940 17149
rect 17974 17115 18016 17149
rect 18050 17115 18108 17149
rect 18142 17115 18200 17149
rect 18234 17115 18263 17149
rect 19027 17117 19056 17151
rect 19090 17117 19138 17151
rect 19172 17117 19230 17151
rect 19264 17117 19322 17151
rect 19356 17117 19385 17151
rect 19893 17119 19922 17153
rect 19956 17119 20012 17153
rect 20046 17119 20104 17153
rect 20138 17119 20196 17153
rect 20230 17119 20259 17153
rect 20680 17143 20738 17214
rect 20817 17373 20863 17432
rect 20897 17454 20913 17455
rect 20897 17420 20911 17454
rect 20947 17420 20963 17455
rect 20897 17407 20963 17420
rect 21431 17452 21477 17491
rect 21531 17487 21577 17503
rect 22305 17505 22321 17539
rect 22355 17505 22371 17539
rect 22305 17493 22371 17505
rect 22405 17607 22451 17653
rect 23007 17643 23036 17677
rect 23070 17643 23128 17677
rect 23162 17643 23220 17677
rect 23254 17643 23310 17677
rect 23344 17643 23373 17677
rect 22439 17573 22451 17607
rect 22405 17539 22451 17573
rect 22439 17505 22451 17539
rect 22305 17460 22351 17493
rect 22405 17489 22451 17505
rect 23073 17597 23139 17609
rect 23073 17563 23089 17597
rect 23123 17563 23139 17597
rect 23073 17529 23139 17563
rect 23073 17495 23089 17529
rect 23123 17495 23139 17529
rect 21431 17418 21433 17452
rect 21469 17418 21477 17452
rect 20817 17355 20883 17373
rect 21431 17371 21477 17418
rect 21511 17419 21527 17453
rect 21561 17448 21577 17453
rect 21511 17414 21537 17419
rect 21571 17414 21577 17448
rect 21511 17405 21577 17414
rect 22305 17426 22307 17460
rect 22341 17426 22351 17460
rect 23073 17483 23139 17495
rect 23173 17597 23219 17643
rect 23207 17563 23219 17597
rect 23173 17529 23219 17563
rect 23207 17495 23219 17529
rect 23298 17549 23356 17643
rect 23298 17515 23310 17549
rect 23344 17515 23356 17549
rect 23298 17498 23356 17515
rect 23073 17456 23119 17483
rect 23173 17479 23219 17495
rect 20817 17321 20833 17355
rect 20867 17321 20883 17355
rect 20817 17287 20883 17321
rect 20817 17253 20833 17287
rect 20867 17253 20883 17287
rect 20817 17219 20883 17253
rect 20817 17185 20833 17219
rect 20867 17185 20883 17219
rect 20817 17177 20883 17185
rect 20917 17355 20959 17371
rect 20951 17321 20959 17355
rect 20917 17287 20959 17321
rect 20951 17253 20959 17287
rect 20917 17219 20959 17253
rect 20951 17185 20959 17219
rect 20917 17143 20959 17185
rect 21431 17353 21497 17371
rect 21431 17319 21447 17353
rect 21481 17319 21497 17353
rect 21431 17285 21497 17319
rect 21431 17251 21447 17285
rect 21481 17251 21497 17285
rect 21431 17217 21497 17251
rect 21431 17183 21447 17217
rect 21481 17183 21497 17217
rect 21431 17175 21497 17183
rect 21531 17353 21573 17369
rect 21565 17319 21573 17353
rect 21531 17285 21573 17319
rect 21565 17251 21573 17285
rect 21531 17217 21573 17251
rect 21565 17183 21573 17217
rect 20663 17109 20692 17143
rect 20726 17109 20780 17143
rect 20814 17109 20872 17143
rect 20906 17109 20964 17143
rect 20998 17109 21027 17143
rect 21531 17141 21573 17183
rect 21658 17339 21716 17374
rect 21658 17305 21670 17339
rect 21704 17305 21716 17339
rect 21658 17246 21716 17305
rect 21658 17212 21670 17246
rect 21704 17212 21716 17246
rect 21658 17141 21716 17212
rect 22166 17341 22224 17376
rect 22166 17307 22178 17341
rect 22212 17307 22224 17341
rect 22166 17248 22224 17307
rect 22166 17214 22178 17248
rect 22212 17214 22224 17248
rect 22166 17143 22224 17214
rect 22305 17373 22351 17426
rect 22385 17452 22401 17455
rect 22385 17418 22397 17452
rect 22435 17418 22451 17455
rect 22385 17407 22451 17418
rect 23073 17422 23079 17456
rect 23117 17422 23119 17456
rect 22305 17355 22371 17373
rect 22305 17321 22321 17355
rect 22355 17321 22371 17355
rect 22305 17287 22371 17321
rect 22305 17253 22321 17287
rect 22355 17253 22371 17287
rect 22305 17219 22371 17253
rect 22305 17185 22321 17219
rect 22355 17185 22371 17219
rect 22305 17177 22371 17185
rect 22405 17355 22447 17371
rect 22439 17321 22447 17355
rect 22405 17287 22447 17321
rect 22439 17253 22447 17287
rect 22405 17219 22447 17253
rect 22439 17185 22447 17219
rect 22405 17143 22447 17185
rect 23073 17363 23119 17422
rect 23153 17444 23169 17445
rect 23153 17410 23167 17444
rect 23203 17410 23219 17445
rect 23153 17397 23219 17410
rect 23073 17345 23139 17363
rect 23073 17311 23089 17345
rect 23123 17311 23139 17345
rect 23073 17277 23139 17311
rect 23073 17243 23089 17277
rect 23123 17243 23139 17277
rect 23073 17209 23139 17243
rect 23073 17175 23089 17209
rect 23123 17175 23139 17209
rect 23073 17167 23139 17175
rect 23173 17345 23215 17361
rect 23207 17311 23215 17345
rect 23173 17277 23215 17311
rect 23207 17243 23215 17277
rect 23173 17209 23215 17243
rect 23207 17175 23215 17209
rect 21365 17107 21394 17141
rect 21428 17107 21486 17141
rect 21520 17107 21578 17141
rect 21612 17107 21670 17141
rect 21704 17107 21733 17141
rect 22149 17109 22178 17143
rect 22212 17109 22268 17143
rect 22302 17109 22360 17143
rect 22394 17109 22452 17143
rect 22486 17109 22515 17143
rect 23173 17133 23215 17175
rect 23298 17331 23356 17366
rect 23298 17297 23310 17331
rect 23344 17297 23356 17331
rect 23298 17238 23356 17297
rect 23298 17204 23310 17238
rect 23344 17204 23356 17238
rect 23298 17133 23356 17204
rect 23007 17099 23036 17133
rect 23070 17099 23128 17133
rect 23162 17099 23220 17133
rect 23254 17099 23310 17133
rect 23344 17099 23373 17133
rect 16246 16677 16275 16711
rect 16309 16677 16365 16711
rect 16399 16677 16457 16711
rect 16491 16677 16549 16711
rect 16583 16677 16612 16711
rect 4376 16569 4405 16603
rect 4439 16569 4497 16603
rect 4531 16569 4589 16603
rect 4623 16569 4681 16603
rect 4715 16569 4773 16603
rect 4807 16569 4865 16603
rect 4899 16569 4957 16603
rect 4991 16569 5049 16603
rect 5083 16569 5112 16603
rect 9242 16573 9271 16607
rect 9305 16573 9363 16607
rect 9397 16573 9455 16607
rect 9489 16573 9547 16607
rect 9581 16573 9639 16607
rect 9673 16573 9731 16607
rect 9765 16573 9823 16607
rect 9857 16573 9915 16607
rect 9949 16573 9978 16607
rect 16263 16606 16321 16677
rect 4393 16498 4451 16569
rect 4393 16464 4405 16498
rect 4439 16464 4451 16498
rect 4393 16405 4451 16464
rect 4393 16371 4405 16405
rect 4439 16371 4451 16405
rect 4393 16336 4451 16371
rect 4485 16527 4561 16535
rect 4485 16493 4511 16527
rect 4545 16493 4561 16527
rect 4485 16459 4561 16493
rect 4485 16425 4511 16459
rect 4545 16425 4561 16459
rect 4485 16399 4561 16425
rect 4679 16517 4713 16569
rect 4679 16449 4713 16483
rect 4679 16399 4713 16415
rect 4747 16517 4813 16535
rect 4747 16483 4763 16517
rect 4797 16483 4813 16517
rect 4747 16449 4813 16483
rect 4847 16517 4881 16569
rect 4847 16467 4881 16483
rect 4915 16517 4995 16535
rect 4915 16483 4951 16517
rect 4985 16483 4995 16517
rect 4747 16415 4763 16449
rect 4797 16433 4813 16449
rect 4915 16449 4995 16483
rect 4915 16433 4951 16449
rect 4797 16415 4951 16433
rect 4985 16415 4995 16449
rect 4747 16399 4995 16415
rect 5031 16519 5095 16535
rect 5031 16485 5035 16519
rect 5069 16485 5095 16519
rect 5031 16451 5095 16485
rect 5031 16417 5035 16451
rect 5069 16417 5095 16451
rect 4485 16207 4519 16399
rect 5031 16390 5095 16417
rect 5031 16383 5044 16390
rect 4553 16331 4814 16365
rect 5031 16349 5035 16383
rect 5078 16352 5095 16390
rect 5069 16349 5095 16352
rect 4553 16292 4602 16331
rect 4553 16291 4554 16292
rect 4588 16258 4602 16292
rect 4587 16257 4602 16258
rect 4636 16294 4746 16297
rect 4636 16291 4674 16294
rect 4636 16257 4670 16291
rect 4708 16260 4746 16294
rect 4704 16257 4746 16260
rect 4780 16291 4814 16331
rect 4969 16315 5095 16349
rect 9259 16502 9317 16573
rect 9259 16468 9271 16502
rect 9305 16468 9317 16502
rect 9259 16409 9317 16468
rect 9259 16375 9271 16409
rect 9305 16375 9317 16409
rect 9259 16340 9317 16375
rect 9351 16531 9427 16539
rect 9351 16497 9377 16531
rect 9411 16497 9427 16531
rect 9351 16463 9427 16497
rect 9351 16429 9377 16463
rect 9411 16429 9427 16463
rect 9351 16403 9427 16429
rect 9545 16521 9579 16573
rect 9545 16453 9579 16487
rect 9545 16403 9579 16419
rect 9613 16521 9679 16539
rect 9613 16487 9629 16521
rect 9663 16487 9679 16521
rect 9613 16453 9679 16487
rect 9713 16521 9747 16573
rect 16263 16572 16275 16606
rect 16309 16572 16321 16606
rect 9713 16471 9747 16487
rect 9781 16521 9861 16539
rect 9781 16487 9817 16521
rect 9851 16487 9861 16521
rect 9613 16419 9629 16453
rect 9663 16437 9679 16453
rect 9781 16453 9861 16487
rect 9781 16437 9817 16453
rect 9663 16419 9817 16437
rect 9851 16419 9861 16453
rect 9613 16403 9861 16419
rect 9897 16523 9961 16539
rect 9897 16489 9901 16523
rect 9935 16489 9961 16523
rect 9897 16455 9961 16489
rect 9897 16421 9901 16455
rect 9935 16421 9961 16455
rect 16263 16513 16321 16572
rect 16263 16479 16275 16513
rect 16309 16479 16321 16513
rect 16263 16444 16321 16479
rect 16404 16635 16446 16677
rect 17104 16667 17133 16701
rect 17167 16667 17225 16701
rect 17259 16667 17317 16701
rect 17351 16667 17407 16701
rect 17441 16667 17470 16701
rect 17886 16669 17915 16703
rect 17949 16669 18007 16703
rect 18041 16669 18099 16703
rect 18133 16669 18191 16703
rect 18225 16669 18254 16703
rect 16404 16601 16412 16635
rect 16404 16567 16446 16601
rect 16404 16533 16412 16567
rect 16404 16499 16446 16533
rect 16404 16465 16412 16499
rect 16404 16449 16446 16465
rect 16480 16635 16546 16643
rect 16480 16601 16496 16635
rect 16530 16601 16546 16635
rect 16480 16567 16546 16601
rect 16480 16533 16496 16567
rect 16530 16533 16546 16567
rect 16480 16499 16546 16533
rect 16480 16465 16496 16499
rect 16530 16465 16546 16499
rect 16480 16447 16546 16465
rect 4889 16291 4935 16307
rect 4780 16257 4805 16291
rect 4839 16257 4855 16291
rect 4889 16257 4901 16291
rect 4553 16241 4602 16257
rect 4889 16207 4935 16257
rect 4393 16187 4451 16204
rect 4393 16153 4405 16187
rect 4439 16153 4451 16187
rect 4485 16173 4935 16207
rect 4393 16059 4451 16153
rect 4595 16159 4629 16173
rect 4495 16103 4511 16137
rect 4545 16103 4561 16137
rect 4969 16139 5003 16315
rect 4595 16109 4629 16125
rect 4495 16059 4561 16103
rect 4663 16103 4679 16137
rect 4713 16103 4729 16137
rect 4812 16105 4847 16139
rect 4881 16105 4947 16139
rect 4981 16105 5003 16139
rect 5037 16210 5095 16226
rect 5071 16176 5095 16210
rect 9351 16211 9385 16403
rect 9897 16394 9961 16421
rect 9897 16387 9910 16394
rect 9419 16335 9680 16369
rect 9897 16353 9901 16387
rect 9944 16356 9961 16394
rect 16400 16400 16466 16413
rect 16400 16365 16416 16400
rect 16452 16366 16466 16400
rect 16450 16365 16466 16366
rect 16500 16388 16546 16447
rect 17172 16625 17214 16667
rect 17172 16591 17180 16625
rect 17172 16557 17214 16591
rect 17172 16523 17180 16557
rect 17172 16489 17214 16523
rect 17172 16455 17180 16489
rect 17172 16439 17214 16455
rect 17248 16625 17314 16633
rect 17248 16591 17264 16625
rect 17298 16591 17314 16625
rect 17248 16557 17314 16591
rect 17248 16523 17264 16557
rect 17298 16523 17314 16557
rect 17248 16489 17314 16523
rect 17248 16455 17264 16489
rect 17298 16455 17314 16489
rect 17248 16437 17314 16455
rect 9935 16353 9961 16356
rect 9419 16296 9468 16335
rect 9419 16295 9420 16296
rect 9454 16262 9468 16296
rect 9453 16261 9468 16262
rect 9502 16298 9612 16301
rect 9502 16295 9540 16298
rect 9502 16261 9536 16295
rect 9574 16264 9612 16298
rect 9570 16261 9612 16264
rect 9646 16295 9680 16335
rect 9835 16319 9961 16353
rect 16500 16354 16502 16388
rect 16540 16354 16546 16388
rect 17168 16392 17234 16403
rect 17168 16355 17184 16392
rect 17222 16358 17234 16392
rect 17218 16355 17234 16358
rect 17268 16384 17314 16437
rect 17395 16596 17453 16667
rect 17395 16562 17407 16596
rect 17441 16562 17453 16596
rect 17395 16503 17453 16562
rect 17395 16469 17407 16503
rect 17441 16469 17453 16503
rect 17395 16434 17453 16469
rect 17903 16598 17961 16669
rect 17903 16564 17915 16598
rect 17949 16564 17961 16598
rect 17903 16505 17961 16564
rect 17903 16471 17915 16505
rect 17949 16471 17961 16505
rect 17903 16436 17961 16471
rect 18046 16627 18088 16669
rect 18592 16667 18621 16701
rect 18655 16667 18713 16701
rect 18747 16667 18805 16701
rect 18839 16667 18893 16701
rect 18927 16667 18956 16701
rect 18046 16593 18054 16627
rect 18046 16559 18088 16593
rect 18046 16525 18054 16559
rect 18046 16491 18088 16525
rect 18046 16457 18054 16491
rect 18046 16441 18088 16457
rect 18122 16627 18188 16635
rect 18122 16593 18138 16627
rect 18172 16593 18188 16627
rect 18122 16559 18188 16593
rect 18122 16525 18138 16559
rect 18172 16525 18188 16559
rect 18122 16491 18188 16525
rect 18122 16457 18138 16491
rect 18172 16457 18188 16491
rect 18122 16439 18188 16457
rect 18660 16625 18702 16667
rect 18660 16591 18668 16625
rect 18660 16557 18702 16591
rect 18660 16523 18668 16557
rect 18660 16489 18702 16523
rect 18660 16455 18668 16489
rect 18660 16439 18702 16455
rect 18736 16625 18802 16633
rect 18736 16591 18752 16625
rect 18786 16591 18802 16625
rect 18736 16557 18802 16591
rect 18736 16523 18752 16557
rect 18786 16523 18802 16557
rect 18736 16489 18802 16523
rect 18736 16455 18752 16489
rect 18786 16455 18802 16489
rect 9755 16295 9801 16311
rect 9646 16261 9671 16295
rect 9705 16261 9721 16295
rect 9755 16261 9767 16295
rect 9419 16245 9468 16261
rect 9755 16211 9801 16261
rect 5037 16142 5095 16176
rect 5071 16108 5095 16142
rect 4663 16059 4729 16103
rect 5037 16059 5095 16108
rect 9259 16191 9317 16208
rect 9259 16157 9271 16191
rect 9305 16157 9317 16191
rect 9351 16177 9801 16211
rect 9259 16063 9317 16157
rect 9461 16163 9495 16177
rect 9361 16107 9377 16141
rect 9411 16107 9427 16141
rect 9835 16143 9869 16319
rect 16400 16315 16446 16331
rect 16500 16327 16546 16354
rect 16263 16295 16321 16312
rect 16263 16261 16275 16295
rect 16309 16261 16321 16295
rect 9461 16113 9495 16129
rect 9361 16063 9427 16107
rect 9529 16107 9545 16141
rect 9579 16107 9595 16141
rect 9678 16109 9713 16143
rect 9747 16109 9813 16143
rect 9847 16109 9869 16143
rect 9903 16214 9961 16230
rect 9937 16180 9961 16214
rect 9903 16146 9961 16180
rect 16263 16167 16321 16261
rect 16400 16281 16412 16315
rect 16400 16247 16446 16281
rect 16400 16213 16412 16247
rect 16400 16167 16446 16213
rect 16480 16315 16546 16327
rect 17268 16350 17278 16384
rect 17312 16350 17314 16384
rect 18042 16396 18108 16405
rect 18042 16362 18048 16396
rect 18082 16391 18108 16396
rect 18042 16357 18058 16362
rect 18092 16357 18108 16391
rect 18142 16392 18188 16439
rect 18736 16437 18802 16455
rect 18142 16358 18150 16392
rect 18186 16358 18188 16392
rect 16480 16281 16496 16315
rect 16530 16281 16546 16315
rect 16480 16247 16546 16281
rect 16480 16213 16496 16247
rect 16530 16213 16546 16247
rect 16480 16201 16546 16213
rect 17168 16305 17214 16321
rect 17268 16317 17314 16350
rect 17168 16271 17180 16305
rect 17168 16237 17214 16271
rect 17168 16203 17180 16237
rect 9937 16112 9961 16146
rect 16246 16133 16275 16167
rect 16309 16133 16365 16167
rect 16399 16133 16457 16167
rect 16491 16133 16549 16167
rect 16583 16133 16612 16167
rect 17168 16157 17214 16203
rect 17248 16305 17314 16317
rect 17248 16271 17264 16305
rect 17298 16271 17314 16305
rect 18042 16307 18088 16323
rect 18142 16319 18188 16358
rect 18656 16390 18722 16403
rect 18656 16355 18672 16390
rect 18708 16356 18722 16390
rect 18706 16355 18722 16356
rect 18756 16378 18802 16437
rect 18881 16596 18939 16667
rect 19360 16657 19389 16691
rect 19423 16657 19481 16691
rect 19515 16657 19573 16691
rect 19607 16657 19663 16691
rect 19697 16657 19726 16691
rect 20234 16659 20263 16693
rect 20297 16659 20355 16693
rect 20389 16659 20447 16693
rect 20481 16659 20529 16693
rect 20563 16659 20592 16693
rect 21356 16661 21385 16695
rect 21419 16661 21477 16695
rect 21511 16661 21569 16695
rect 21603 16661 21645 16695
rect 21679 16661 21708 16695
rect 18881 16562 18893 16596
rect 18927 16562 18939 16596
rect 18881 16503 18939 16562
rect 18881 16469 18893 16503
rect 18927 16469 18939 16503
rect 18881 16434 18939 16469
rect 19428 16615 19470 16657
rect 19428 16581 19436 16615
rect 19428 16547 19470 16581
rect 19428 16513 19436 16547
rect 19428 16479 19470 16513
rect 19428 16445 19436 16479
rect 19428 16429 19470 16445
rect 19504 16615 19570 16623
rect 19504 16581 19520 16615
rect 19554 16581 19570 16615
rect 19504 16547 19570 16581
rect 19504 16513 19520 16547
rect 19554 16513 19570 16547
rect 19504 16479 19570 16513
rect 19504 16445 19520 16479
rect 19554 16445 19570 16479
rect 19504 16427 19570 16445
rect 18756 16344 18758 16378
rect 18796 16344 18802 16378
rect 19424 16382 19490 16393
rect 19424 16345 19440 16382
rect 19478 16348 19490 16382
rect 19474 16345 19490 16348
rect 19524 16374 19570 16427
rect 19651 16586 19709 16657
rect 19651 16552 19663 16586
rect 19697 16552 19709 16586
rect 19651 16493 19709 16552
rect 19651 16459 19663 16493
rect 19697 16459 19709 16493
rect 19651 16424 19709 16459
rect 20302 16617 20344 16659
rect 20302 16583 20310 16617
rect 20302 16549 20344 16583
rect 20302 16515 20310 16549
rect 20302 16481 20344 16515
rect 20302 16447 20310 16481
rect 20302 16431 20344 16447
rect 20378 16617 20444 16625
rect 20378 16583 20394 16617
rect 20428 16583 20444 16617
rect 20378 16549 20444 16583
rect 20378 16515 20394 16549
rect 20428 16515 20444 16549
rect 20378 16481 20444 16515
rect 20378 16447 20394 16481
rect 20428 16447 20444 16481
rect 20378 16429 20444 16447
rect 17248 16237 17314 16271
rect 17248 16203 17264 16237
rect 17298 16203 17314 16237
rect 17248 16191 17314 16203
rect 17395 16285 17453 16302
rect 17395 16251 17407 16285
rect 17441 16251 17453 16285
rect 17395 16157 17453 16251
rect 17903 16287 17961 16304
rect 17903 16253 17915 16287
rect 17949 16253 17961 16287
rect 17903 16159 17961 16253
rect 18042 16273 18054 16307
rect 18042 16239 18088 16273
rect 18042 16205 18054 16239
rect 18042 16159 18088 16205
rect 18122 16307 18188 16319
rect 18122 16273 18138 16307
rect 18172 16273 18188 16307
rect 18122 16239 18188 16273
rect 18122 16205 18138 16239
rect 18172 16205 18188 16239
rect 18122 16193 18188 16205
rect 18656 16305 18702 16321
rect 18756 16317 18802 16344
rect 18656 16271 18668 16305
rect 18656 16237 18702 16271
rect 18656 16203 18668 16237
rect 17104 16123 17133 16157
rect 17167 16123 17225 16157
rect 17259 16123 17317 16157
rect 17351 16123 17407 16157
rect 17441 16123 17470 16157
rect 17886 16125 17915 16159
rect 17949 16125 18007 16159
rect 18041 16125 18099 16159
rect 18133 16125 18191 16159
rect 18225 16125 18254 16159
rect 18656 16157 18702 16203
rect 18736 16305 18802 16317
rect 19524 16340 19534 16374
rect 19568 16340 19570 16374
rect 20298 16386 20364 16395
rect 20298 16352 20304 16386
rect 20338 16381 20364 16386
rect 20298 16347 20314 16352
rect 20348 16347 20364 16381
rect 20398 16382 20444 16429
rect 20517 16588 20575 16659
rect 20517 16554 20529 16588
rect 20563 16554 20575 16588
rect 20517 16495 20575 16554
rect 20517 16461 20529 16495
rect 20563 16461 20575 16495
rect 20517 16426 20575 16461
rect 21424 16619 21466 16661
rect 21424 16585 21432 16619
rect 21424 16551 21466 16585
rect 21424 16517 21432 16551
rect 21424 16483 21466 16517
rect 21424 16449 21432 16483
rect 21424 16433 21466 16449
rect 21500 16619 21566 16627
rect 21500 16585 21516 16619
rect 21550 16585 21566 16619
rect 21500 16551 21566 16585
rect 21500 16517 21516 16551
rect 21550 16517 21566 16551
rect 21500 16483 21566 16517
rect 21500 16449 21516 16483
rect 21550 16449 21566 16483
rect 21500 16431 21566 16449
rect 20398 16348 20406 16382
rect 20442 16348 20444 16382
rect 21420 16384 21486 16397
rect 21420 16349 21436 16384
rect 21472 16350 21486 16384
rect 21470 16349 21486 16350
rect 21520 16372 21566 16431
rect 21633 16590 21691 16661
rect 22124 16651 22153 16685
rect 22187 16651 22245 16685
rect 22279 16651 22337 16685
rect 22371 16651 22423 16685
rect 22457 16651 22486 16685
rect 22998 16653 23027 16687
rect 23061 16653 23119 16687
rect 23153 16653 23211 16687
rect 23245 16653 23289 16687
rect 23323 16653 23352 16687
rect 21633 16556 21645 16590
rect 21679 16556 21691 16590
rect 21633 16497 21691 16556
rect 21633 16463 21645 16497
rect 21679 16463 21691 16497
rect 21633 16428 21691 16463
rect 22192 16609 22234 16651
rect 22192 16575 22200 16609
rect 22192 16541 22234 16575
rect 22192 16507 22200 16541
rect 22192 16473 22234 16507
rect 22192 16439 22200 16473
rect 22192 16423 22234 16439
rect 22268 16609 22334 16617
rect 22268 16575 22284 16609
rect 22318 16575 22334 16609
rect 22268 16541 22334 16575
rect 22268 16507 22284 16541
rect 22318 16507 22334 16541
rect 22268 16473 22334 16507
rect 22268 16439 22284 16473
rect 22318 16439 22334 16473
rect 22268 16421 22334 16439
rect 18736 16271 18752 16305
rect 18786 16271 18802 16305
rect 18736 16237 18802 16271
rect 18736 16203 18752 16237
rect 18786 16203 18802 16237
rect 18736 16191 18802 16203
rect 18881 16285 18939 16302
rect 18881 16251 18893 16285
rect 18927 16251 18939 16285
rect 18881 16157 18939 16251
rect 19424 16295 19470 16311
rect 19524 16307 19570 16340
rect 19424 16261 19436 16295
rect 19424 16227 19470 16261
rect 19424 16193 19436 16227
rect 18592 16123 18621 16157
rect 18655 16123 18713 16157
rect 18747 16123 18805 16157
rect 18839 16123 18893 16157
rect 18927 16123 18956 16157
rect 19424 16147 19470 16193
rect 19504 16295 19570 16307
rect 19504 16261 19520 16295
rect 19554 16261 19570 16295
rect 20298 16297 20344 16313
rect 20398 16309 20444 16348
rect 21520 16338 21522 16372
rect 21560 16338 21566 16372
rect 22188 16376 22254 16387
rect 22188 16339 22204 16376
rect 22242 16342 22254 16376
rect 22238 16339 22254 16342
rect 22288 16368 22334 16421
rect 22411 16580 22469 16651
rect 22411 16546 22423 16580
rect 22457 16546 22469 16580
rect 22411 16487 22469 16546
rect 22411 16453 22423 16487
rect 22457 16453 22469 16487
rect 22411 16418 22469 16453
rect 23066 16611 23108 16653
rect 23066 16577 23074 16611
rect 23066 16543 23108 16577
rect 23066 16509 23074 16543
rect 23066 16475 23108 16509
rect 23066 16441 23074 16475
rect 23066 16425 23108 16441
rect 23142 16611 23208 16619
rect 23142 16577 23158 16611
rect 23192 16577 23208 16611
rect 23142 16543 23208 16577
rect 23142 16509 23158 16543
rect 23192 16509 23208 16543
rect 23142 16475 23208 16509
rect 23142 16441 23158 16475
rect 23192 16441 23208 16475
rect 23142 16423 23208 16441
rect 19504 16227 19570 16261
rect 19504 16193 19520 16227
rect 19554 16193 19570 16227
rect 19504 16181 19570 16193
rect 19651 16275 19709 16292
rect 19651 16241 19663 16275
rect 19697 16241 19709 16275
rect 19651 16147 19709 16241
rect 20298 16263 20310 16297
rect 20298 16229 20344 16263
rect 20298 16195 20310 16229
rect 20298 16149 20344 16195
rect 20378 16297 20444 16309
rect 20378 16263 20394 16297
rect 20428 16263 20444 16297
rect 21420 16299 21466 16315
rect 21520 16311 21566 16338
rect 20378 16229 20444 16263
rect 20378 16195 20394 16229
rect 20428 16195 20444 16229
rect 20378 16183 20444 16195
rect 20517 16277 20575 16294
rect 20517 16243 20529 16277
rect 20563 16243 20575 16277
rect 20517 16149 20575 16243
rect 21420 16265 21432 16299
rect 21420 16231 21466 16265
rect 21420 16197 21432 16231
rect 21420 16151 21466 16197
rect 21500 16299 21566 16311
rect 22288 16334 22298 16368
rect 22332 16334 22334 16368
rect 23062 16380 23128 16389
rect 23062 16346 23068 16380
rect 23102 16375 23128 16380
rect 23062 16341 23078 16346
rect 23112 16341 23128 16375
rect 23162 16376 23208 16423
rect 23277 16582 23335 16653
rect 23277 16548 23289 16582
rect 23323 16548 23335 16582
rect 23277 16489 23335 16548
rect 23277 16455 23289 16489
rect 23323 16455 23335 16489
rect 23277 16420 23335 16455
rect 23162 16342 23170 16376
rect 23206 16342 23208 16376
rect 21500 16265 21516 16299
rect 21550 16265 21566 16299
rect 21500 16231 21566 16265
rect 21500 16197 21516 16231
rect 21550 16197 21566 16231
rect 21500 16185 21566 16197
rect 21633 16279 21691 16296
rect 21633 16245 21645 16279
rect 21679 16245 21691 16279
rect 21633 16151 21691 16245
rect 22188 16289 22234 16305
rect 22288 16301 22334 16334
rect 22188 16255 22200 16289
rect 22188 16221 22234 16255
rect 22188 16187 22200 16221
rect 19360 16113 19389 16147
rect 19423 16113 19481 16147
rect 19515 16113 19573 16147
rect 19607 16113 19663 16147
rect 19697 16113 19726 16147
rect 20234 16115 20263 16149
rect 20297 16115 20355 16149
rect 20389 16115 20447 16149
rect 20481 16115 20529 16149
rect 20563 16115 20592 16149
rect 21356 16117 21385 16151
rect 21419 16117 21477 16151
rect 21511 16117 21569 16151
rect 21603 16117 21645 16151
rect 21679 16117 21708 16151
rect 22188 16141 22234 16187
rect 22268 16289 22334 16301
rect 22268 16255 22284 16289
rect 22318 16255 22334 16289
rect 23062 16291 23108 16307
rect 23162 16303 23208 16342
rect 22268 16221 22334 16255
rect 22268 16187 22284 16221
rect 22318 16187 22334 16221
rect 22268 16175 22334 16187
rect 22411 16269 22469 16286
rect 22411 16235 22423 16269
rect 22457 16235 22469 16269
rect 22411 16141 22469 16235
rect 23062 16257 23074 16291
rect 23062 16223 23108 16257
rect 23062 16189 23074 16223
rect 23062 16143 23108 16189
rect 23142 16291 23208 16303
rect 23142 16257 23158 16291
rect 23192 16257 23208 16291
rect 23142 16223 23208 16257
rect 23142 16189 23158 16223
rect 23192 16189 23208 16223
rect 23142 16177 23208 16189
rect 23277 16271 23335 16288
rect 23277 16237 23289 16271
rect 23323 16237 23335 16271
rect 23277 16143 23335 16237
rect 9529 16063 9595 16107
rect 9903 16063 9961 16112
rect 22124 16107 22153 16141
rect 22187 16107 22245 16141
rect 22279 16107 22337 16141
rect 22371 16107 22423 16141
rect 22457 16107 22486 16141
rect 22998 16109 23027 16143
rect 23061 16109 23119 16143
rect 23153 16109 23211 16143
rect 23245 16109 23289 16143
rect 23323 16109 23352 16143
rect 4376 16025 4405 16059
rect 4439 16025 4497 16059
rect 4531 16025 4589 16059
rect 4623 16025 4681 16059
rect 4715 16025 4773 16059
rect 4807 16025 4865 16059
rect 4899 16025 4957 16059
rect 4991 16025 5049 16059
rect 5083 16025 5112 16059
rect 9242 16029 9271 16063
rect 9305 16029 9363 16063
rect 9397 16029 9455 16063
rect 9489 16029 9547 16063
rect 9581 16029 9639 16063
rect 9673 16029 9731 16063
rect 9765 16029 9823 16063
rect 9857 16029 9915 16063
rect 9949 16029 9978 16063
rect 4476 15825 4505 15859
rect 4539 15825 4595 15859
rect 4629 15825 4687 15859
rect 4721 15825 4779 15859
rect 4813 15825 4871 15859
rect 4905 15825 4963 15859
rect 4997 15825 5026 15859
rect 9342 15829 9371 15863
rect 9405 15829 9461 15863
rect 9495 15829 9553 15863
rect 9587 15829 9645 15863
rect 9679 15829 9737 15863
rect 9771 15829 9829 15863
rect 9863 15829 9892 15863
rect 4493 15754 4551 15825
rect 4493 15720 4505 15754
rect 4539 15720 4551 15754
rect 4493 15661 4551 15720
rect 4623 15741 4679 15825
rect 4813 15783 4879 15825
rect 4623 15707 4637 15741
rect 4671 15707 4679 15741
rect 4623 15691 4679 15707
rect 4713 15741 4773 15757
rect 4713 15707 4721 15741
rect 4755 15707 4773 15741
rect 4493 15627 4505 15661
rect 4539 15627 4551 15661
rect 4713 15647 4773 15707
rect 4813 15749 4829 15783
rect 4863 15749 4879 15783
rect 4813 15715 4879 15749
rect 4813 15681 4829 15715
rect 4863 15681 4879 15715
rect 4917 15783 5009 15791
rect 4917 15749 4933 15783
rect 4967 15749 5009 15783
rect 9359 15758 9417 15829
rect 4917 15715 5009 15749
rect 6608 15715 6637 15749
rect 6671 15715 6729 15749
rect 6763 15715 6821 15749
rect 6855 15715 6913 15749
rect 6947 15715 7005 15749
rect 7039 15715 7097 15749
rect 7131 15715 7189 15749
rect 7223 15715 7281 15749
rect 7315 15715 7344 15749
rect 9359 15724 9371 15758
rect 9405 15724 9417 15758
rect 4917 15681 4933 15715
rect 4967 15681 5009 15715
rect 4493 15592 4551 15627
rect 4586 15570 4639 15635
rect 4713 15613 4901 15647
rect 4586 15530 4588 15570
rect 4630 15563 4639 15570
rect 4867 15563 4901 15613
rect 4630 15547 4721 15563
rect 4630 15530 4640 15547
rect 4586 15513 4640 15530
rect 4674 15513 4721 15547
rect 4765 15560 4833 15563
rect 4765 15520 4778 15560
rect 4820 15520 4833 15560
rect 4765 15513 4781 15520
rect 4815 15513 4833 15520
rect 4867 15547 4925 15563
rect 4867 15513 4889 15547
rect 4923 15513 4925 15547
rect 4867 15497 4925 15513
rect 4867 15479 4901 15497
rect 4493 15443 4551 15460
rect 4493 15409 4505 15443
rect 4539 15409 4551 15443
rect 4493 15315 4551 15409
rect 4623 15441 4901 15479
rect 4959 15490 5009 15681
rect 6626 15673 6693 15715
rect 6626 15639 6643 15673
rect 6677 15639 6693 15673
rect 6727 15665 6777 15681
rect 6727 15631 6735 15665
rect 6769 15631 6777 15665
rect 4959 15456 4970 15490
rect 5006 15456 5009 15490
rect 4623 15419 4689 15441
rect 4623 15385 4637 15419
rect 4671 15385 4689 15419
rect 4959 15407 5009 15456
rect 4623 15369 4689 15385
rect 4813 15391 4863 15407
rect 4813 15357 4829 15391
rect 4813 15315 4863 15357
rect 4897 15391 5009 15407
rect 4897 15357 4913 15391
rect 4947 15357 5009 15391
rect 4897 15349 5009 15357
rect 6625 15437 6673 15603
rect 6727 15521 6777 15631
rect 6821 15673 6887 15715
rect 6821 15639 6837 15673
rect 6871 15639 6887 15673
rect 6821 15571 6887 15639
rect 6924 15665 6974 15681
rect 6924 15631 6932 15665
rect 6966 15631 6974 15665
rect 6924 15521 6974 15631
rect 7067 15673 7133 15715
rect 7067 15639 7083 15673
rect 7117 15639 7133 15673
rect 7067 15605 7133 15639
rect 7167 15673 7235 15681
rect 7167 15639 7183 15673
rect 7217 15639 7235 15673
rect 7167 15629 7235 15639
rect 7067 15571 7083 15605
rect 7117 15571 7133 15605
rect 7067 15555 7133 15571
rect 7183 15605 7235 15629
rect 7217 15571 7235 15605
rect 7183 15537 7235 15571
rect 6625 15403 6639 15437
rect 6625 15400 6673 15403
rect 6625 15364 6632 15400
rect 6668 15364 6673 15400
rect 6625 15341 6673 15364
rect 6707 15487 7145 15521
rect 4476 15281 4505 15315
rect 4539 15281 4595 15315
rect 4629 15281 4687 15315
rect 4721 15281 4779 15315
rect 4813 15281 4871 15315
rect 4905 15281 4963 15315
rect 4997 15281 5026 15315
rect 6707 15305 6741 15487
rect 7082 15453 7145 15487
rect 7217 15503 7235 15537
rect 6642 15289 6741 15305
rect 6642 15255 6643 15289
rect 6677 15255 6741 15289
rect 6785 15437 6855 15453
rect 6819 15434 6855 15437
rect 6785 15398 6804 15403
rect 6838 15398 6855 15434
rect 6785 15260 6855 15398
rect 6891 15437 6951 15453
rect 6925 15403 6951 15437
rect 6891 15310 6951 15403
rect 6891 15276 6902 15310
rect 6936 15276 6951 15310
rect 6891 15259 6951 15276
rect 6987 15437 7043 15453
rect 7021 15403 7043 15437
rect 7082 15437 7148 15453
rect 7082 15403 7098 15437
rect 7132 15403 7148 15437
rect 7183 15432 7235 15503
rect 7269 15644 7327 15715
rect 7269 15610 7281 15644
rect 7315 15610 7327 15644
rect 7269 15551 7327 15610
rect 9359 15665 9417 15724
rect 9489 15745 9545 15829
rect 9679 15787 9745 15829
rect 9489 15711 9503 15745
rect 9537 15711 9545 15745
rect 9489 15695 9545 15711
rect 9579 15745 9639 15761
rect 9579 15711 9587 15745
rect 9621 15711 9639 15745
rect 9359 15631 9371 15665
rect 9405 15631 9417 15665
rect 9579 15651 9639 15711
rect 9679 15753 9695 15787
rect 9729 15753 9745 15787
rect 9679 15719 9745 15753
rect 9679 15685 9695 15719
rect 9729 15685 9745 15719
rect 9783 15787 9875 15795
rect 9783 15753 9799 15787
rect 9833 15753 9875 15787
rect 9783 15719 9875 15753
rect 11474 15719 11503 15753
rect 11537 15719 11595 15753
rect 11629 15719 11687 15753
rect 11721 15719 11779 15753
rect 11813 15719 11871 15753
rect 11905 15719 11963 15753
rect 11997 15719 12055 15753
rect 12089 15719 12147 15753
rect 12181 15719 12210 15753
rect 9783 15685 9799 15719
rect 9833 15685 9875 15719
rect 9359 15596 9417 15631
rect 7269 15517 7281 15551
rect 7315 15517 7327 15551
rect 9452 15574 9505 15639
rect 9579 15617 9767 15651
rect 9452 15534 9454 15574
rect 9496 15567 9505 15574
rect 9733 15567 9767 15617
rect 9496 15551 9587 15567
rect 9496 15534 9506 15551
rect 9452 15517 9506 15534
rect 9540 15517 9587 15551
rect 9631 15564 9699 15567
rect 9631 15524 9644 15564
rect 9686 15524 9699 15564
rect 9631 15517 9647 15524
rect 9681 15517 9699 15524
rect 9733 15551 9791 15567
rect 9733 15517 9755 15551
rect 9789 15517 9791 15551
rect 7269 15482 7327 15517
rect 9733 15501 9791 15517
rect 9733 15483 9767 15501
rect 6987 15380 7043 15403
rect 6987 15344 6998 15380
rect 7032 15344 7043 15380
rect 7183 15398 7190 15432
rect 7224 15398 7235 15432
rect 6987 15259 7043 15344
rect 7079 15349 7133 15365
rect 7183 15349 7235 15398
rect 9359 15447 9417 15464
rect 9359 15413 9371 15447
rect 9405 15413 9417 15447
rect 7079 15315 7084 15349
rect 7118 15315 7133 15349
rect 7079 15281 7133 15315
rect 5750 15215 5779 15249
rect 5813 15215 5871 15249
rect 5905 15215 5963 15249
rect 5997 15215 6055 15249
rect 6089 15215 6147 15249
rect 6181 15215 6239 15249
rect 6273 15215 6302 15249
rect 6642 15239 6741 15255
rect 7079 15247 7084 15281
rect 7118 15247 7133 15281
rect 7167 15315 7183 15349
rect 7217 15315 7235 15349
rect 7167 15281 7235 15315
rect 7167 15247 7183 15281
rect 7217 15247 7235 15281
rect 7269 15333 7327 15350
rect 7269 15299 7281 15333
rect 7315 15299 7327 15333
rect 9359 15319 9417 15413
rect 9489 15445 9767 15483
rect 9825 15494 9875 15685
rect 11492 15677 11559 15719
rect 11492 15643 11509 15677
rect 11543 15643 11559 15677
rect 11593 15669 11643 15685
rect 11593 15635 11601 15669
rect 11635 15635 11643 15669
rect 9825 15460 9836 15494
rect 9872 15460 9875 15494
rect 9489 15423 9555 15445
rect 9489 15389 9503 15423
rect 9537 15389 9555 15423
rect 9825 15411 9875 15460
rect 9489 15373 9555 15389
rect 9679 15395 9729 15411
rect 9679 15361 9695 15395
rect 9679 15319 9729 15361
rect 9763 15395 9875 15411
rect 9763 15361 9779 15395
rect 9813 15361 9875 15395
rect 9763 15353 9875 15361
rect 11491 15441 11539 15607
rect 11593 15525 11643 15635
rect 11687 15677 11753 15719
rect 11687 15643 11703 15677
rect 11737 15643 11753 15677
rect 11687 15575 11753 15643
rect 11790 15669 11840 15685
rect 11790 15635 11798 15669
rect 11832 15635 11840 15669
rect 11790 15525 11840 15635
rect 11933 15677 11999 15719
rect 11933 15643 11949 15677
rect 11983 15643 11999 15677
rect 11933 15609 11999 15643
rect 12033 15677 12101 15685
rect 12033 15643 12049 15677
rect 12083 15643 12101 15677
rect 12033 15633 12101 15643
rect 11933 15575 11949 15609
rect 11983 15575 11999 15609
rect 11933 15559 11999 15575
rect 12049 15609 12101 15633
rect 12083 15575 12101 15609
rect 12049 15541 12101 15575
rect 11491 15407 11505 15441
rect 11491 15404 11539 15407
rect 11491 15368 11498 15404
rect 11534 15368 11539 15404
rect 11491 15345 11539 15368
rect 11573 15491 12011 15525
rect 5807 15131 5863 15215
rect 5997 15173 6063 15215
rect 5807 15097 5821 15131
rect 5855 15097 5863 15131
rect 5807 15081 5863 15097
rect 5897 15131 5957 15147
rect 5897 15097 5905 15131
rect 5939 15097 5957 15131
rect 4386 15005 4415 15039
rect 4449 15005 4507 15039
rect 4541 15005 4599 15039
rect 4633 15005 4691 15039
rect 4725 15005 4783 15039
rect 4817 15005 4875 15039
rect 4909 15005 4967 15039
rect 5001 15005 5059 15039
rect 5093 15005 5122 15039
rect 5897 15037 5957 15097
rect 5997 15139 6013 15173
rect 6047 15139 6063 15173
rect 5997 15105 6063 15139
rect 5997 15071 6013 15105
rect 6047 15071 6063 15105
rect 6101 15173 6193 15181
rect 6101 15139 6117 15173
rect 6151 15148 6193 15173
rect 6101 15112 6144 15139
rect 6184 15112 6193 15148
rect 6101 15105 6193 15112
rect 6101 15071 6117 15105
rect 6151 15071 6193 15105
rect 4403 14934 4461 15005
rect 4403 14900 4415 14934
rect 4449 14900 4461 14934
rect 4403 14841 4461 14900
rect 4403 14807 4415 14841
rect 4449 14807 4461 14841
rect 4403 14772 4461 14807
rect 4495 14963 4571 14971
rect 4495 14929 4521 14963
rect 4555 14929 4571 14963
rect 4495 14895 4571 14929
rect 4495 14861 4521 14895
rect 4555 14861 4571 14895
rect 4495 14835 4571 14861
rect 4689 14953 4723 15005
rect 4689 14885 4723 14919
rect 4689 14835 4723 14851
rect 4757 14953 4823 14971
rect 4757 14919 4773 14953
rect 4807 14919 4823 14953
rect 4757 14885 4823 14919
rect 4857 14953 4891 15005
rect 4857 14903 4891 14919
rect 4925 14953 5005 14971
rect 4925 14919 4961 14953
rect 4995 14919 5005 14953
rect 4757 14851 4773 14885
rect 4807 14869 4823 14885
rect 4925 14885 5005 14919
rect 4925 14869 4961 14885
rect 4807 14851 4961 14869
rect 4995 14851 5005 14885
rect 4757 14835 5005 14851
rect 5041 14955 5105 14971
rect 5041 14921 5045 14955
rect 5079 14930 5105 14955
rect 5041 14896 5056 14921
rect 5090 14896 5105 14930
rect 5770 14953 5823 15025
rect 5897 15003 6085 15037
rect 6051 14953 6085 15003
rect 5770 14938 5905 14953
rect 5770 14903 5824 14938
rect 5858 14903 5905 14938
rect 5949 14938 6017 14953
rect 5949 14904 5964 14938
rect 6000 14904 6017 14938
rect 5949 14903 5965 14904
rect 5999 14903 6017 14904
rect 6051 14937 6109 14953
rect 6051 14903 6073 14937
rect 6107 14903 6109 14937
rect 5041 14887 5105 14896
rect 5041 14853 5045 14887
rect 5079 14853 5105 14887
rect 6051 14887 6109 14903
rect 6051 14869 6085 14887
rect 4495 14643 4529 14835
rect 5041 14819 5105 14853
rect 4563 14767 4824 14801
rect 5041 14785 5045 14819
rect 5079 14785 5105 14819
rect 4563 14728 4612 14767
rect 4563 14727 4564 14728
rect 4598 14694 4612 14728
rect 4597 14693 4612 14694
rect 4646 14730 4756 14733
rect 4646 14727 4684 14730
rect 4646 14693 4680 14727
rect 4718 14696 4756 14730
rect 4714 14693 4756 14696
rect 4790 14727 4824 14767
rect 4979 14751 5105 14785
rect 5807 14831 6085 14869
rect 5807 14809 5873 14831
rect 5807 14775 5821 14809
rect 5855 14775 5873 14809
rect 6143 14797 6193 15071
rect 6227 15144 6285 15215
rect 7079 15205 7133 15247
rect 7269 15205 7327 15299
rect 9342 15285 9371 15319
rect 9405 15285 9461 15319
rect 9495 15285 9553 15319
rect 9587 15285 9645 15319
rect 9679 15285 9737 15319
rect 9771 15285 9829 15319
rect 9863 15285 9892 15319
rect 11573 15309 11607 15491
rect 11948 15457 12011 15491
rect 12083 15507 12101 15541
rect 11508 15293 11607 15309
rect 11508 15259 11509 15293
rect 11543 15259 11607 15293
rect 11651 15441 11721 15457
rect 11685 15438 11721 15441
rect 11651 15402 11670 15407
rect 11704 15402 11721 15438
rect 11651 15264 11721 15402
rect 11757 15441 11817 15457
rect 11791 15407 11817 15441
rect 11757 15314 11817 15407
rect 11757 15280 11768 15314
rect 11802 15280 11817 15314
rect 11757 15263 11817 15280
rect 11853 15441 11909 15457
rect 11887 15407 11909 15441
rect 11948 15441 12014 15457
rect 11948 15407 11964 15441
rect 11998 15407 12014 15441
rect 12049 15436 12101 15507
rect 12135 15648 12193 15719
rect 12135 15614 12147 15648
rect 12181 15614 12193 15648
rect 12135 15555 12193 15614
rect 12135 15521 12147 15555
rect 12181 15521 12193 15555
rect 12135 15486 12193 15521
rect 11853 15384 11909 15407
rect 11853 15348 11864 15384
rect 11898 15348 11909 15384
rect 12049 15402 12056 15436
rect 12090 15402 12101 15436
rect 11853 15263 11909 15348
rect 11945 15353 11999 15369
rect 12049 15353 12101 15402
rect 11945 15319 11950 15353
rect 11984 15319 11999 15353
rect 11945 15285 11999 15319
rect 10616 15219 10645 15253
rect 10679 15219 10737 15253
rect 10771 15219 10829 15253
rect 10863 15219 10921 15253
rect 10955 15219 11013 15253
rect 11047 15219 11105 15253
rect 11139 15219 11168 15253
rect 11508 15243 11607 15259
rect 11945 15251 11950 15285
rect 11984 15251 11999 15285
rect 12033 15319 12049 15353
rect 12083 15319 12101 15353
rect 12033 15285 12101 15319
rect 12033 15251 12049 15285
rect 12083 15251 12101 15285
rect 12135 15337 12193 15354
rect 12135 15303 12147 15337
rect 12181 15303 12193 15337
rect 6608 15171 6637 15205
rect 6671 15171 6729 15205
rect 6763 15171 6821 15205
rect 6855 15171 6913 15205
rect 6947 15171 7005 15205
rect 7039 15171 7097 15205
rect 7131 15171 7189 15205
rect 7223 15171 7281 15205
rect 7315 15171 7344 15205
rect 6227 15110 6239 15144
rect 6273 15110 6285 15144
rect 6227 15051 6285 15110
rect 10673 15135 10729 15219
rect 10863 15177 10929 15219
rect 10673 15101 10687 15135
rect 10721 15101 10729 15135
rect 10673 15085 10729 15101
rect 10763 15135 10823 15151
rect 10763 15101 10771 15135
rect 10805 15101 10823 15135
rect 6227 15017 6239 15051
rect 6273 15017 6285 15051
rect 6227 14982 6285 15017
rect 9252 15009 9281 15043
rect 9315 15009 9373 15043
rect 9407 15009 9465 15043
rect 9499 15009 9557 15043
rect 9591 15009 9649 15043
rect 9683 15009 9741 15043
rect 9775 15009 9833 15043
rect 9867 15009 9925 15043
rect 9959 15009 9988 15043
rect 10763 15041 10823 15101
rect 10863 15143 10879 15177
rect 10913 15143 10929 15177
rect 10863 15109 10929 15143
rect 10863 15075 10879 15109
rect 10913 15075 10929 15109
rect 10967 15177 11059 15185
rect 10967 15143 10983 15177
rect 11017 15152 11059 15177
rect 10967 15116 11010 15143
rect 11050 15116 11059 15152
rect 10967 15109 11059 15116
rect 10967 15075 10983 15109
rect 11017 15075 11059 15109
rect 9269 14938 9327 15009
rect 9269 14904 9281 14938
rect 9315 14904 9327 14938
rect 5807 14759 5873 14775
rect 5997 14781 6047 14797
rect 4899 14727 4945 14743
rect 4790 14693 4815 14727
rect 4849 14693 4865 14727
rect 4899 14693 4911 14727
rect 4563 14677 4612 14693
rect 4899 14643 4945 14693
rect 4403 14623 4461 14640
rect 4403 14589 4415 14623
rect 4449 14589 4461 14623
rect 4495 14609 4945 14643
rect 4403 14495 4461 14589
rect 4605 14595 4639 14609
rect 4505 14539 4521 14573
rect 4555 14539 4571 14573
rect 4979 14575 5013 14751
rect 5997 14747 6013 14781
rect 5997 14705 6047 14747
rect 6081 14781 6193 14797
rect 6081 14747 6097 14781
rect 6131 14747 6193 14781
rect 6081 14739 6193 14747
rect 6227 14833 6285 14850
rect 6227 14799 6239 14833
rect 6273 14799 6285 14833
rect 6227 14705 6285 14799
rect 9269 14845 9327 14904
rect 9269 14811 9281 14845
rect 9315 14811 9327 14845
rect 9269 14776 9327 14811
rect 9361 14967 9437 14975
rect 9361 14933 9387 14967
rect 9421 14933 9437 14967
rect 9361 14899 9437 14933
rect 9361 14865 9387 14899
rect 9421 14865 9437 14899
rect 9361 14839 9437 14865
rect 9555 14957 9589 15009
rect 9555 14889 9589 14923
rect 9555 14839 9589 14855
rect 9623 14957 9689 14975
rect 9623 14923 9639 14957
rect 9673 14923 9689 14957
rect 9623 14889 9689 14923
rect 9723 14957 9757 15009
rect 9723 14907 9757 14923
rect 9791 14957 9871 14975
rect 9791 14923 9827 14957
rect 9861 14923 9871 14957
rect 9623 14855 9639 14889
rect 9673 14873 9689 14889
rect 9791 14889 9871 14923
rect 9791 14873 9827 14889
rect 9673 14855 9827 14873
rect 9861 14855 9871 14889
rect 9623 14839 9871 14855
rect 9907 14959 9971 14975
rect 9907 14925 9911 14959
rect 9945 14934 9971 14959
rect 9907 14900 9922 14925
rect 9956 14900 9971 14934
rect 10636 14957 10689 15029
rect 10763 15007 10951 15041
rect 10917 14957 10951 15007
rect 10636 14942 10771 14957
rect 10636 14907 10690 14942
rect 10724 14907 10771 14942
rect 10815 14942 10883 14957
rect 10815 14908 10830 14942
rect 10866 14908 10883 14942
rect 10815 14907 10831 14908
rect 10865 14907 10883 14908
rect 10917 14941 10975 14957
rect 10917 14907 10939 14941
rect 10973 14907 10975 14941
rect 9907 14891 9971 14900
rect 9907 14857 9911 14891
rect 9945 14857 9971 14891
rect 10917 14891 10975 14907
rect 10917 14873 10951 14891
rect 5750 14671 5779 14705
rect 5813 14671 5871 14705
rect 5905 14671 5963 14705
rect 5997 14671 6055 14705
rect 6089 14671 6147 14705
rect 6181 14671 6239 14705
rect 6273 14671 6302 14705
rect 4605 14545 4639 14561
rect 4505 14495 4571 14539
rect 4673 14539 4689 14573
rect 4723 14539 4739 14573
rect 4822 14541 4857 14575
rect 4891 14541 4957 14575
rect 4991 14541 5013 14575
rect 5047 14646 5105 14662
rect 5081 14612 5105 14646
rect 9361 14647 9395 14839
rect 9907 14823 9971 14857
rect 9429 14771 9690 14805
rect 9907 14789 9911 14823
rect 9945 14789 9971 14823
rect 9429 14732 9478 14771
rect 9429 14731 9430 14732
rect 9464 14698 9478 14732
rect 9463 14697 9478 14698
rect 9512 14734 9622 14737
rect 9512 14731 9550 14734
rect 9512 14697 9546 14731
rect 9584 14700 9622 14734
rect 9580 14697 9622 14700
rect 9656 14731 9690 14771
rect 9845 14755 9971 14789
rect 10673 14835 10951 14873
rect 10673 14813 10739 14835
rect 10673 14779 10687 14813
rect 10721 14779 10739 14813
rect 11009 14801 11059 15075
rect 11093 15148 11151 15219
rect 11945 15209 11999 15251
rect 12135 15209 12193 15303
rect 11474 15175 11503 15209
rect 11537 15175 11595 15209
rect 11629 15175 11687 15209
rect 11721 15175 11779 15209
rect 11813 15175 11871 15209
rect 11905 15175 11963 15209
rect 11997 15175 12055 15209
rect 12089 15175 12147 15209
rect 12181 15175 12210 15209
rect 11093 15114 11105 15148
rect 11139 15114 11151 15148
rect 11093 15055 11151 15114
rect 11093 15021 11105 15055
rect 11139 15021 11151 15055
rect 11093 14986 11151 15021
rect 10673 14763 10739 14779
rect 10863 14785 10913 14801
rect 9765 14731 9811 14747
rect 9656 14697 9681 14731
rect 9715 14697 9731 14731
rect 9765 14697 9777 14731
rect 9429 14681 9478 14697
rect 9765 14647 9811 14697
rect 5047 14578 5105 14612
rect 5081 14544 5105 14578
rect 4673 14495 4739 14539
rect 5047 14495 5105 14544
rect 9269 14627 9327 14644
rect 9269 14593 9281 14627
rect 9315 14593 9327 14627
rect 9361 14613 9811 14647
rect 9269 14499 9327 14593
rect 9471 14599 9505 14613
rect 9371 14543 9387 14577
rect 9421 14543 9437 14577
rect 9845 14579 9879 14755
rect 10863 14751 10879 14785
rect 10863 14709 10913 14751
rect 10947 14785 11059 14801
rect 10947 14751 10963 14785
rect 10997 14751 11059 14785
rect 10947 14743 11059 14751
rect 11093 14837 11151 14854
rect 11093 14803 11105 14837
rect 11139 14803 11151 14837
rect 23484 14815 23513 14849
rect 23547 14815 23605 14849
rect 23639 14815 23697 14849
rect 23731 14815 23789 14849
rect 23823 14815 23881 14849
rect 23915 14815 23973 14849
rect 24007 14815 24065 14849
rect 24099 14815 24157 14849
rect 24191 14815 24249 14849
rect 24283 14815 24341 14849
rect 24375 14815 24433 14849
rect 24467 14815 24525 14849
rect 24559 14815 24617 14849
rect 24651 14815 24709 14849
rect 24743 14815 24801 14849
rect 24835 14815 24893 14849
rect 24927 14815 24985 14849
rect 25019 14815 25077 14849
rect 25111 14815 25169 14849
rect 25203 14815 25261 14849
rect 25295 14815 25353 14849
rect 25387 14815 25445 14849
rect 25479 14815 25508 14849
rect 11093 14709 11151 14803
rect 23519 14765 23553 14781
rect 23587 14773 23653 14815
rect 23587 14739 23603 14773
rect 23637 14739 23653 14773
rect 23687 14765 23993 14781
rect 10616 14675 10645 14709
rect 10679 14675 10737 14709
rect 10771 14675 10829 14709
rect 10863 14675 10921 14709
rect 10955 14675 11013 14709
rect 11047 14675 11105 14709
rect 11139 14675 11168 14709
rect 23519 14681 23553 14731
rect 23721 14747 23993 14765
rect 23687 14715 23721 14731
rect 23791 14697 23825 14713
rect 9471 14549 9505 14565
rect 9371 14499 9437 14543
rect 9539 14543 9555 14577
rect 9589 14543 9605 14577
rect 9688 14545 9723 14579
rect 9757 14545 9823 14579
rect 9857 14545 9879 14579
rect 9913 14650 9971 14666
rect 9947 14616 9971 14650
rect 23519 14663 23791 14681
rect 23519 14647 23825 14663
rect 23859 14679 23875 14713
rect 23909 14679 23925 14713
rect 23959 14697 23993 14747
rect 9913 14582 9971 14616
rect 23859 14613 23893 14679
rect 23959 14647 23993 14663
rect 24027 14765 24097 14781
rect 24027 14731 24063 14765
rect 24131 14773 24197 14815
rect 24131 14739 24147 14773
rect 24181 14739 24197 14773
rect 24249 14747 24451 14781
rect 24027 14613 24097 14731
rect 24249 14697 24283 14747
rect 9947 14548 9971 14582
rect 9539 14499 9605 14543
rect 9913 14499 9971 14548
rect 23514 14580 23583 14611
rect 23514 14546 23530 14580
rect 23568 14546 23583 14580
rect 23514 14537 23583 14546
rect 23514 14503 23549 14537
rect 4386 14461 4415 14495
rect 4449 14461 4507 14495
rect 4541 14461 4599 14495
rect 4633 14461 4691 14495
rect 4725 14461 4783 14495
rect 4817 14461 4875 14495
rect 4909 14461 4967 14495
rect 5001 14461 5059 14495
rect 5093 14461 5122 14495
rect 9252 14465 9281 14499
rect 9315 14465 9373 14499
rect 9407 14465 9465 14499
rect 9499 14465 9557 14499
rect 9591 14465 9649 14499
rect 9683 14465 9741 14499
rect 9775 14465 9833 14499
rect 9867 14465 9925 14499
rect 9959 14465 9988 14499
rect 23514 14487 23583 14503
rect 23645 14562 23732 14611
rect 23645 14537 23672 14562
rect 23708 14528 23732 14562
rect 23679 14503 23732 14528
rect 23645 14487 23732 14503
rect 23766 14579 23893 14613
rect 23766 14475 23800 14579
rect 23936 14567 24097 14613
rect 24137 14650 24197 14687
rect 24137 14616 24150 14650
rect 24186 14616 24197 14650
rect 24249 14645 24283 14663
rect 24317 14679 24333 14713
rect 24367 14679 24383 14713
rect 24317 14645 24349 14679
rect 24417 14705 24451 14747
rect 24496 14773 24562 14815
rect 24496 14739 24512 14773
rect 24546 14739 24562 14773
rect 24596 14765 24630 14781
rect 24680 14773 24750 14815
rect 24680 14739 24700 14773
rect 24734 14739 24750 14773
rect 24784 14765 24821 14781
rect 24596 14705 24630 14731
rect 24818 14731 24821 14765
rect 24784 14715 24821 14731
rect 24417 14671 24630 14705
rect 23936 14545 24008 14567
rect 23900 14511 23916 14545
rect 23950 14543 24008 14545
rect 23950 14511 23974 14543
rect 23900 14509 23974 14511
rect 23519 14415 23721 14449
rect 23519 14390 23553 14415
rect 23519 14340 23553 14356
rect 23587 14347 23603 14381
rect 23637 14347 23653 14381
rect 23587 14305 23653 14347
rect 23687 14373 23721 14415
rect 23766 14441 23790 14475
rect 23766 14407 23784 14441
rect 23818 14407 23834 14441
rect 23868 14415 23902 14440
rect 23868 14373 23902 14381
rect 23936 14424 24008 14509
rect 24137 14541 24197 14616
rect 24317 14611 24383 14645
rect 24137 14507 24150 14541
rect 24184 14507 24197 14541
rect 24137 14487 24197 14507
rect 24231 14577 24383 14611
rect 24231 14472 24265 14577
rect 24444 14552 24493 14623
rect 24299 14507 24315 14541
rect 24444 14518 24456 14552
rect 24492 14549 24493 14552
rect 24444 14515 24459 14518
rect 24349 14507 24365 14509
rect 24444 14499 24493 14515
rect 24534 14588 24600 14623
rect 24534 14554 24556 14588
rect 24592 14554 24600 14588
rect 24534 14549 24600 14554
rect 24534 14515 24566 14549
rect 24534 14499 24600 14515
rect 24695 14562 24753 14623
rect 24695 14537 24712 14562
rect 24746 14528 24753 14562
rect 24729 14503 24753 14528
rect 24695 14487 24753 14503
rect 24787 14543 24821 14715
rect 24880 14765 24922 14781
rect 24880 14731 24888 14765
rect 24956 14773 25213 14781
rect 24956 14739 24972 14773
rect 25006 14747 25213 14773
rect 25006 14739 25022 14747
rect 24880 14715 24922 14731
rect 24787 14509 24811 14543
rect 24231 14457 24294 14472
rect 23936 14390 23972 14424
rect 24006 14390 24008 14424
rect 23936 14374 24008 14390
rect 24044 14433 24102 14449
rect 24044 14399 24056 14433
rect 24090 14399 24102 14433
rect 23687 14339 23902 14373
rect 24044 14305 24102 14399
rect 24160 14431 24194 14447
rect 24228 14423 24244 14457
rect 24278 14423 24294 14457
rect 24228 14407 24294 14423
rect 24328 14465 24362 14473
rect 24328 14457 24632 14465
rect 24362 14431 24632 14457
rect 24328 14407 24362 14423
rect 24583 14397 24632 14431
rect 24787 14419 24821 14509
rect 24880 14475 24914 14715
rect 25053 14685 25069 14713
rect 24962 14679 25069 14685
rect 25103 14679 25119 14713
rect 24962 14645 24995 14679
rect 25029 14645 25119 14679
rect 24962 14639 25119 14645
rect 25179 14655 25213 14747
rect 25247 14773 25313 14815
rect 25247 14739 25263 14773
rect 25297 14739 25313 14773
rect 25347 14765 25399 14781
rect 25381 14731 25399 14765
rect 24880 14441 24894 14475
rect 24160 14373 24194 14397
rect 24514 14381 24548 14397
rect 24409 14373 24430 14381
rect 24160 14347 24430 14373
rect 24464 14347 24480 14381
rect 24160 14339 24480 14347
rect 24583 14363 24598 14397
rect 24786 14403 24821 14419
rect 24962 14405 24996 14639
rect 25179 14621 25309 14655
rect 25122 14509 25138 14543
rect 25172 14509 25179 14543
rect 25275 14537 25309 14621
rect 25112 14473 25160 14475
rect 25112 14457 25161 14473
rect 25275 14465 25309 14503
rect 25112 14441 25127 14457
rect 25126 14423 25127 14441
rect 25126 14407 25161 14423
rect 25195 14431 25309 14465
rect 25347 14594 25399 14731
rect 25347 14560 25356 14594
rect 25390 14560 25399 14594
rect 25433 14744 25491 14815
rect 25433 14710 25445 14744
rect 25479 14710 25491 14744
rect 25433 14651 25491 14710
rect 25433 14617 25445 14651
rect 25479 14617 25491 14651
rect 25433 14582 25491 14617
rect 24583 14347 24632 14363
rect 24686 14347 24702 14381
rect 24736 14347 24752 14381
rect 24820 14369 24821 14403
rect 24786 14353 24821 14369
rect 24890 14389 24996 14405
rect 24924 14371 24996 14389
rect 25030 14389 25064 14405
rect 24514 14305 24548 14347
rect 24686 14305 24752 14347
rect 24890 14339 24924 14355
rect 25195 14373 25229 14431
rect 25064 14355 25229 14373
rect 25030 14339 25229 14355
rect 25263 14381 25297 14397
rect 25263 14305 25297 14347
rect 25347 14389 25399 14560
rect 25381 14355 25399 14389
rect 25347 14339 25399 14355
rect 25433 14433 25491 14450
rect 25433 14399 25445 14433
rect 25479 14399 25491 14433
rect 25433 14305 25491 14399
rect 4486 14261 4515 14295
rect 4549 14261 4605 14295
rect 4639 14261 4697 14295
rect 4731 14261 4789 14295
rect 4823 14261 4881 14295
rect 4915 14261 4973 14295
rect 5007 14261 5036 14295
rect 4503 14190 4561 14261
rect 4503 14156 4515 14190
rect 4549 14156 4561 14190
rect 4503 14097 4561 14156
rect 4633 14177 4689 14261
rect 4823 14219 4889 14261
rect 5732 14249 5761 14283
rect 5795 14249 5853 14283
rect 5887 14249 5945 14283
rect 5979 14249 6037 14283
rect 6071 14249 6129 14283
rect 6163 14249 6221 14283
rect 6255 14249 6313 14283
rect 6347 14249 6405 14283
rect 6439 14249 6468 14283
rect 4633 14143 4647 14177
rect 4681 14143 4689 14177
rect 4633 14127 4689 14143
rect 4723 14177 4783 14193
rect 4723 14143 4731 14177
rect 4765 14143 4783 14177
rect 4503 14063 4515 14097
rect 4549 14063 4561 14097
rect 4723 14083 4783 14143
rect 4823 14185 4839 14219
rect 4873 14185 4889 14219
rect 4823 14151 4889 14185
rect 4823 14117 4839 14151
rect 4873 14117 4889 14151
rect 4927 14219 5019 14227
rect 4927 14185 4943 14219
rect 4977 14185 5019 14219
rect 4927 14151 5019 14185
rect 4927 14117 4943 14151
rect 4977 14117 5019 14151
rect 4503 14028 4561 14063
rect 4596 14006 4649 14071
rect 4723 14049 4911 14083
rect 4596 13966 4598 14006
rect 4640 13999 4649 14006
rect 4877 13999 4911 14049
rect 4640 13983 4731 13999
rect 4640 13966 4650 13983
rect 4596 13949 4650 13966
rect 4684 13949 4731 13983
rect 4775 13996 4843 13999
rect 4775 13956 4788 13996
rect 4830 13956 4843 13996
rect 4775 13949 4791 13956
rect 4825 13949 4843 13956
rect 4877 13983 4935 13999
rect 4877 13949 4899 13983
rect 4933 13949 4935 13983
rect 4877 13933 4935 13949
rect 4877 13915 4911 13933
rect 4503 13879 4561 13896
rect 4503 13845 4515 13879
rect 4549 13845 4561 13879
rect 4503 13751 4561 13845
rect 4633 13877 4911 13915
rect 4969 13884 5019 14117
rect 5749 14178 5807 14249
rect 5749 14144 5761 14178
rect 5795 14144 5807 14178
rect 5842 14207 5909 14249
rect 5842 14173 5859 14207
rect 5893 14173 5909 14207
rect 5943 14199 5993 14215
rect 5749 14085 5807 14144
rect 5943 14165 5951 14199
rect 5985 14165 5993 14199
rect 5749 14051 5761 14085
rect 5795 14051 5807 14085
rect 5749 14016 5807 14051
rect 5841 13976 5889 14137
rect 5943 14055 5993 14165
rect 6037 14207 6103 14249
rect 6037 14173 6053 14207
rect 6087 14173 6103 14207
rect 6037 14105 6103 14173
rect 6140 14199 6190 14215
rect 6140 14165 6148 14199
rect 6182 14165 6190 14199
rect 6140 14055 6190 14165
rect 6283 14207 6349 14249
rect 7722 14233 7751 14267
rect 7785 14233 7843 14267
rect 7877 14233 7935 14267
rect 7969 14233 8027 14267
rect 8061 14233 8119 14267
rect 8153 14233 8211 14267
rect 8245 14233 8303 14267
rect 8337 14233 8366 14267
rect 9350 14265 9379 14299
rect 9413 14265 9471 14299
rect 9505 14265 9563 14299
rect 9597 14265 9655 14299
rect 9689 14265 9747 14299
rect 9781 14265 9839 14299
rect 9873 14265 9902 14299
rect 6283 14173 6299 14207
rect 6333 14173 6349 14207
rect 6283 14139 6349 14173
rect 6383 14207 6451 14215
rect 6383 14173 6399 14207
rect 6433 14173 6451 14207
rect 8105 14191 8161 14233
rect 6383 14163 6451 14173
rect 6283 14105 6299 14139
rect 6333 14105 6349 14139
rect 6283 14089 6349 14105
rect 6399 14139 6451 14163
rect 6433 14105 6451 14139
rect 7740 14179 8071 14189
rect 7740 14166 7979 14179
rect 7740 14132 7896 14166
rect 7932 14145 7979 14166
rect 8013 14145 8071 14179
rect 7932 14132 8071 14145
rect 7740 14131 8071 14132
rect 8105 14157 8118 14191
rect 8152 14157 8161 14191
rect 6399 14071 6451 14105
rect 8105 14123 8161 14157
rect 5841 13942 5850 13976
rect 5884 13971 5889 13976
rect 5841 13937 5855 13942
rect 4633 13855 4699 13877
rect 4633 13821 4647 13855
rect 4681 13821 4699 13855
rect 4969 13850 4978 13884
rect 5014 13850 5019 13884
rect 4969 13843 5019 13850
rect 4633 13805 4699 13821
rect 4823 13827 4873 13843
rect 4823 13793 4839 13827
rect 4823 13751 4873 13793
rect 4907 13827 5019 13843
rect 4907 13793 4923 13827
rect 4957 13793 5019 13827
rect 4907 13785 5019 13793
rect 5749 13867 5807 13884
rect 5841 13875 5889 13937
rect 5923 14021 6361 14055
rect 5749 13833 5761 13867
rect 5795 13833 5807 13867
rect 5923 13839 5957 14021
rect 6298 13987 6361 14021
rect 6433 14037 6451 14071
rect 4486 13717 4515 13751
rect 4549 13717 4605 13751
rect 4639 13717 4697 13751
rect 4731 13717 4789 13751
rect 4823 13717 4881 13751
rect 4915 13717 4973 13751
rect 5007 13717 5036 13751
rect 5749 13739 5807 13833
rect 5858 13823 5957 13839
rect 5858 13789 5859 13823
rect 5893 13789 5957 13823
rect 6001 13971 6071 13987
rect 6035 13937 6071 13971
rect 6001 13880 6071 13937
rect 6001 13846 6020 13880
rect 6054 13846 6071 13880
rect 6001 13794 6071 13846
rect 6107 13971 6167 13987
rect 6141 13937 6167 13971
rect 6107 13920 6167 13937
rect 6107 13886 6118 13920
rect 6152 13886 6167 13920
rect 6107 13793 6167 13886
rect 6203 13971 6259 13987
rect 6237 13970 6259 13971
rect 6203 13932 6212 13937
rect 6248 13932 6259 13970
rect 6298 13971 6364 13987
rect 6298 13937 6314 13971
rect 6348 13937 6364 13971
rect 6203 13793 6259 13932
rect 6295 13883 6349 13899
rect 6399 13883 6451 14037
rect 7740 14063 8058 14097
rect 8105 14089 8118 14123
rect 8152 14089 8161 14123
rect 8105 14073 8161 14089
rect 8203 14160 8257 14199
rect 8237 14126 8257 14160
rect 8203 14092 8257 14126
rect 8237 14076 8257 14092
rect 7740 14060 7804 14063
rect 7740 14026 7757 14060
rect 7791 14026 7804 14060
rect 8024 14039 8058 14063
rect 7740 14005 7804 14026
rect 7740 13955 7810 13971
rect 7740 13938 7757 13955
rect 7791 13938 7810 13955
rect 6295 13849 6300 13883
rect 6334 13849 6349 13883
rect 6295 13815 6349 13849
rect 5858 13773 5957 13789
rect 6295 13781 6300 13815
rect 6334 13781 6349 13815
rect 6383 13852 6399 13883
rect 6383 13814 6394 13852
rect 6433 13849 6451 13883
rect 6794 13875 6823 13909
rect 6857 13875 6915 13909
rect 6949 13875 7007 13909
rect 7041 13875 7099 13909
rect 7133 13875 7191 13909
rect 7225 13875 7279 13909
rect 7313 13875 7342 13909
rect 7740 13904 7752 13938
rect 7792 13904 7810 13938
rect 7844 13960 7986 14029
rect 8024 14005 8169 14039
rect 8203 14036 8212 14058
rect 8254 14036 8257 14076
rect 8203 14005 8257 14036
rect 8135 13971 8169 14005
rect 7844 13918 7880 13960
rect 7930 13918 7986 13960
rect 7844 13905 7986 13918
rect 8020 13956 8101 13971
rect 8020 13920 8052 13956
rect 8090 13955 8101 13956
rect 8093 13921 8101 13955
rect 8090 13920 8101 13921
rect 8020 13905 8101 13920
rect 8135 13955 8189 13971
rect 8135 13921 8155 13955
rect 8135 13905 8189 13921
rect 6432 13815 6451 13849
rect 6383 13781 6399 13814
rect 6433 13781 6451 13815
rect 7023 13817 7089 13875
rect 7023 13783 7039 13817
rect 7073 13783 7089 13817
rect 6295 13739 6349 13781
rect 7023 13749 7089 13783
rect 5732 13705 5761 13739
rect 5795 13705 5853 13739
rect 5887 13705 5945 13739
rect 5979 13705 6037 13739
rect 6071 13705 6129 13739
rect 6163 13705 6221 13739
rect 6255 13705 6313 13739
rect 6347 13705 6405 13739
rect 6439 13705 6468 13739
rect 6848 13697 6926 13716
rect 7023 13715 7039 13749
rect 7073 13715 7089 13749
rect 7123 13833 7230 13841
rect 7123 13799 7139 13833
rect 7173 13799 7230 13833
rect 7123 13765 7230 13799
rect 7123 13731 7139 13765
rect 7173 13764 7230 13765
rect 7123 13730 7162 13731
rect 7196 13730 7230 13764
rect 7123 13717 7230 13730
rect 6848 13663 6870 13697
rect 6904 13681 6926 13697
rect 6904 13663 7133 13681
rect 6848 13647 7133 13663
rect 6823 13597 6894 13613
rect 6823 13563 6860 13597
rect 6823 13554 6894 13563
rect 6823 13520 6834 13554
rect 6868 13520 6894 13554
rect 6823 13501 6894 13520
rect 6928 13467 6962 13647
rect 6996 13604 7049 13613
rect 6996 13597 7012 13604
rect 7046 13570 7049 13604
rect 7030 13563 7049 13570
rect 6996 13501 7049 13563
rect 7099 13597 7133 13647
rect 7099 13547 7133 13563
rect 7167 13513 7230 13717
rect 7267 13804 7325 13875
rect 7740 13857 7810 13904
rect 8135 13871 8169 13905
rect 7847 13837 8169 13871
rect 8223 13858 8257 14005
rect 8291 14162 8349 14233
rect 8291 14128 8303 14162
rect 8337 14128 8349 14162
rect 8291 14069 8349 14128
rect 8291 14035 8303 14069
rect 8337 14035 8349 14069
rect 8291 14000 8349 14035
rect 9367 14194 9425 14265
rect 9367 14160 9379 14194
rect 9413 14160 9425 14194
rect 9367 14101 9425 14160
rect 9499 14181 9555 14265
rect 9689 14223 9755 14265
rect 10598 14253 10627 14287
rect 10661 14253 10719 14287
rect 10753 14253 10811 14287
rect 10845 14253 10903 14287
rect 10937 14253 10995 14287
rect 11029 14253 11087 14287
rect 11121 14253 11179 14287
rect 11213 14253 11271 14287
rect 11305 14253 11334 14287
rect 23484 14271 23513 14305
rect 23547 14271 23605 14305
rect 23639 14271 23697 14305
rect 23731 14271 23789 14305
rect 23823 14271 23881 14305
rect 23915 14271 23973 14305
rect 24007 14271 24065 14305
rect 24099 14271 24157 14305
rect 24191 14271 24249 14305
rect 24283 14271 24341 14305
rect 24375 14271 24433 14305
rect 24467 14271 24525 14305
rect 24559 14271 24617 14305
rect 24651 14271 24709 14305
rect 24743 14271 24801 14305
rect 24835 14271 24893 14305
rect 24927 14271 24985 14305
rect 25019 14271 25077 14305
rect 25111 14271 25169 14305
rect 25203 14271 25261 14305
rect 25295 14271 25353 14305
rect 25387 14271 25445 14305
rect 25479 14271 25508 14305
rect 9499 14147 9513 14181
rect 9547 14147 9555 14181
rect 9499 14131 9555 14147
rect 9589 14181 9649 14197
rect 9589 14147 9597 14181
rect 9631 14147 9649 14181
rect 9367 14067 9379 14101
rect 9413 14067 9425 14101
rect 9589 14087 9649 14147
rect 9689 14189 9705 14223
rect 9739 14189 9755 14223
rect 9689 14155 9755 14189
rect 9689 14121 9705 14155
rect 9739 14121 9755 14155
rect 9793 14223 9885 14231
rect 9793 14189 9809 14223
rect 9843 14189 9885 14223
rect 9793 14155 9885 14189
rect 9793 14121 9809 14155
rect 9843 14121 9885 14155
rect 9367 14032 9425 14067
rect 9462 14010 9515 14075
rect 9589 14053 9777 14087
rect 9462 13970 9464 14010
rect 9506 14003 9515 14010
rect 9743 14003 9777 14053
rect 9506 13987 9597 14003
rect 9506 13970 9516 13987
rect 9462 13953 9516 13970
rect 9550 13953 9597 13987
rect 9641 14000 9709 14003
rect 9641 13960 9654 14000
rect 9696 13960 9709 14000
rect 9641 13953 9657 13960
rect 9691 13953 9709 13960
rect 9743 13987 9801 14003
rect 9743 13953 9765 13987
rect 9799 13953 9801 13987
rect 9743 13937 9801 13953
rect 9743 13919 9777 13937
rect 9367 13883 9425 13900
rect 8203 13841 8257 13858
rect 7267 13770 7279 13804
rect 7313 13770 7325 13804
rect 7267 13711 7325 13770
rect 7741 13789 7757 13823
rect 7791 13789 7807 13823
rect 7741 13723 7807 13789
rect 7847 13817 7881 13837
rect 8021 13817 8055 13837
rect 7847 13767 7881 13783
rect 7921 13769 7937 13803
rect 7971 13769 7987 13803
rect 7921 13723 7987 13769
rect 8237 13807 8257 13841
rect 8021 13767 8055 13783
rect 8089 13769 8115 13803
rect 8149 13769 8165 13803
rect 8203 13789 8257 13807
rect 8291 13851 8349 13868
rect 8291 13817 8303 13851
rect 8337 13817 8349 13851
rect 8089 13723 8165 13769
rect 8291 13723 8349 13817
rect 9367 13849 9379 13883
rect 9413 13849 9425 13883
rect 9367 13755 9425 13849
rect 9499 13881 9777 13919
rect 9835 13888 9885 14121
rect 10615 14182 10673 14253
rect 10615 14148 10627 14182
rect 10661 14148 10673 14182
rect 10708 14211 10775 14253
rect 10708 14177 10725 14211
rect 10759 14177 10775 14211
rect 10809 14203 10859 14219
rect 10615 14089 10673 14148
rect 10809 14169 10817 14203
rect 10851 14169 10859 14203
rect 10615 14055 10627 14089
rect 10661 14055 10673 14089
rect 10615 14020 10673 14055
rect 10707 13980 10755 14141
rect 10809 14059 10859 14169
rect 10903 14211 10969 14253
rect 10903 14177 10919 14211
rect 10953 14177 10969 14211
rect 10903 14109 10969 14177
rect 11006 14203 11056 14219
rect 11006 14169 11014 14203
rect 11048 14169 11056 14203
rect 11006 14059 11056 14169
rect 11149 14211 11215 14253
rect 12588 14237 12617 14271
rect 12651 14237 12709 14271
rect 12743 14237 12801 14271
rect 12835 14237 12893 14271
rect 12927 14237 12985 14271
rect 13019 14237 13077 14271
rect 13111 14237 13169 14271
rect 13203 14237 13232 14271
rect 11149 14177 11165 14211
rect 11199 14177 11215 14211
rect 11149 14143 11215 14177
rect 11249 14211 11317 14219
rect 11249 14177 11265 14211
rect 11299 14177 11317 14211
rect 12971 14195 13027 14237
rect 11249 14167 11317 14177
rect 11149 14109 11165 14143
rect 11199 14109 11215 14143
rect 11149 14093 11215 14109
rect 11265 14143 11317 14167
rect 11299 14109 11317 14143
rect 12606 14183 12937 14193
rect 12606 14170 12845 14183
rect 12606 14136 12762 14170
rect 12798 14149 12845 14170
rect 12879 14149 12937 14183
rect 12798 14136 12937 14149
rect 12606 14135 12937 14136
rect 12971 14161 12984 14195
rect 13018 14161 13027 14195
rect 11265 14075 11317 14109
rect 12971 14127 13027 14161
rect 10707 13946 10716 13980
rect 10750 13975 10755 13980
rect 10707 13941 10721 13946
rect 9499 13859 9565 13881
rect 9499 13825 9513 13859
rect 9547 13825 9565 13859
rect 9835 13854 9844 13888
rect 9880 13854 9885 13888
rect 9835 13847 9885 13854
rect 9499 13809 9565 13825
rect 9689 13831 9739 13847
rect 9689 13797 9705 13831
rect 9689 13755 9739 13797
rect 9773 13831 9885 13847
rect 9773 13797 9789 13831
rect 9823 13797 9885 13831
rect 9773 13789 9885 13797
rect 10615 13871 10673 13888
rect 10707 13879 10755 13941
rect 10789 14025 11227 14059
rect 10615 13837 10627 13871
rect 10661 13837 10673 13871
rect 10789 13843 10823 14025
rect 11164 13991 11227 14025
rect 11299 14041 11317 14075
rect 7267 13677 7279 13711
rect 7313 13677 7325 13711
rect 7722 13689 7751 13723
rect 7785 13689 7843 13723
rect 7877 13689 7935 13723
rect 7969 13689 8027 13723
rect 8061 13689 8119 13723
rect 8153 13689 8211 13723
rect 8245 13689 8303 13723
rect 8337 13689 8366 13723
rect 9350 13721 9379 13755
rect 9413 13721 9471 13755
rect 9505 13721 9563 13755
rect 9597 13721 9655 13755
rect 9689 13721 9747 13755
rect 9781 13721 9839 13755
rect 9873 13721 9902 13755
rect 10615 13743 10673 13837
rect 10724 13827 10823 13843
rect 10724 13793 10725 13827
rect 10759 13793 10823 13827
rect 10867 13975 10937 13991
rect 10901 13941 10937 13975
rect 10867 13884 10937 13941
rect 10867 13850 10886 13884
rect 10920 13850 10937 13884
rect 10867 13798 10937 13850
rect 10973 13975 11033 13991
rect 11007 13941 11033 13975
rect 10973 13924 11033 13941
rect 10973 13890 10984 13924
rect 11018 13890 11033 13924
rect 10973 13797 11033 13890
rect 11069 13975 11125 13991
rect 11103 13974 11125 13975
rect 11069 13936 11078 13941
rect 11114 13936 11125 13974
rect 11164 13975 11230 13991
rect 11164 13941 11180 13975
rect 11214 13941 11230 13975
rect 11069 13797 11125 13936
rect 11161 13887 11215 13903
rect 11265 13887 11317 14041
rect 12606 14067 12924 14101
rect 12971 14093 12984 14127
rect 13018 14093 13027 14127
rect 12971 14077 13027 14093
rect 13069 14164 13123 14203
rect 13103 14130 13123 14164
rect 13069 14096 13123 14130
rect 13103 14080 13123 14096
rect 12606 14064 12670 14067
rect 12606 14030 12623 14064
rect 12657 14030 12670 14064
rect 12890 14043 12924 14067
rect 12606 14009 12670 14030
rect 12606 13959 12676 13975
rect 12606 13942 12623 13959
rect 12657 13942 12676 13959
rect 11161 13853 11166 13887
rect 11200 13853 11215 13887
rect 11161 13819 11215 13853
rect 10724 13777 10823 13793
rect 11161 13785 11166 13819
rect 11200 13785 11215 13819
rect 11249 13856 11265 13887
rect 11249 13818 11260 13856
rect 11299 13853 11317 13887
rect 11660 13879 11689 13913
rect 11723 13879 11781 13913
rect 11815 13879 11873 13913
rect 11907 13879 11965 13913
rect 11999 13879 12057 13913
rect 12091 13879 12147 13913
rect 12181 13879 12210 13913
rect 12606 13908 12618 13942
rect 12658 13908 12676 13942
rect 12710 13964 12852 14033
rect 12890 14009 13035 14043
rect 13069 14040 13078 14062
rect 13120 14040 13123 14080
rect 13069 14009 13123 14040
rect 13001 13975 13035 14009
rect 12710 13922 12746 13964
rect 12796 13922 12852 13964
rect 12710 13909 12852 13922
rect 12886 13960 12967 13975
rect 12886 13924 12918 13960
rect 12956 13959 12967 13960
rect 12959 13925 12967 13959
rect 12956 13924 12967 13925
rect 12886 13909 12967 13924
rect 13001 13959 13055 13975
rect 13001 13925 13021 13959
rect 13001 13909 13055 13925
rect 11298 13819 11317 13853
rect 11249 13785 11265 13818
rect 11299 13785 11317 13819
rect 11889 13821 11955 13879
rect 11889 13787 11905 13821
rect 11939 13787 11955 13821
rect 11161 13743 11215 13785
rect 11889 13753 11955 13787
rect 10598 13709 10627 13743
rect 10661 13709 10719 13743
rect 10753 13709 10811 13743
rect 10845 13709 10903 13743
rect 10937 13709 10995 13743
rect 11029 13709 11087 13743
rect 11121 13709 11179 13743
rect 11213 13709 11271 13743
rect 11305 13709 11334 13743
rect 11714 13701 11792 13720
rect 11889 13719 11905 13753
rect 11939 13719 11955 13753
rect 11989 13837 12096 13845
rect 11989 13803 12005 13837
rect 12039 13803 12096 13837
rect 11989 13769 12096 13803
rect 11989 13735 12005 13769
rect 12039 13768 12096 13769
rect 11989 13734 12028 13735
rect 12062 13734 12096 13768
rect 11989 13721 12096 13734
rect 7267 13642 7325 13677
rect 11714 13667 11736 13701
rect 11770 13685 11792 13701
rect 11770 13667 11999 13685
rect 11714 13651 11999 13667
rect 7107 13511 7230 13513
rect 7107 13477 7123 13511
rect 7157 13477 7230 13511
rect 11689 13601 11760 13617
rect 11689 13567 11726 13601
rect 11689 13558 11760 13567
rect 11689 13524 11700 13558
rect 11734 13524 11760 13558
rect 6844 13451 6892 13467
rect 5856 13407 5885 13441
rect 5919 13407 5977 13441
rect 6011 13407 6069 13441
rect 6103 13407 6161 13441
rect 6195 13407 6253 13441
rect 6287 13407 6345 13441
rect 6379 13407 6408 13441
rect 6844 13417 6858 13451
rect 4378 13337 4407 13371
rect 4441 13337 4499 13371
rect 4533 13337 4591 13371
rect 4625 13337 4683 13371
rect 4717 13337 4775 13371
rect 4809 13337 4867 13371
rect 4901 13337 4959 13371
rect 4993 13337 5051 13371
rect 5085 13337 5114 13371
rect 4395 13266 4453 13337
rect 4395 13232 4407 13266
rect 4441 13232 4453 13266
rect 4395 13173 4453 13232
rect 4395 13139 4407 13173
rect 4441 13139 4453 13173
rect 4395 13104 4453 13139
rect 4487 13295 4563 13303
rect 4487 13261 4513 13295
rect 4547 13261 4563 13295
rect 4487 13227 4563 13261
rect 4487 13193 4513 13227
rect 4547 13193 4563 13227
rect 4487 13167 4563 13193
rect 4681 13285 4715 13337
rect 4681 13217 4715 13251
rect 4681 13167 4715 13183
rect 4749 13285 4815 13303
rect 4749 13251 4765 13285
rect 4799 13251 4815 13285
rect 4749 13217 4815 13251
rect 4849 13285 4883 13337
rect 5873 13336 5931 13407
rect 4849 13235 4883 13251
rect 4917 13285 4997 13303
rect 4917 13251 4953 13285
rect 4987 13251 4997 13285
rect 4749 13183 4765 13217
rect 4799 13201 4815 13217
rect 4917 13217 4997 13251
rect 4917 13201 4953 13217
rect 4799 13183 4953 13201
rect 4987 13183 4997 13217
rect 4749 13167 4997 13183
rect 5033 13287 5097 13303
rect 5033 13253 5037 13287
rect 5071 13253 5097 13287
rect 5033 13220 5097 13253
rect 5033 13219 5048 13220
rect 5033 13185 5037 13219
rect 5082 13186 5097 13220
rect 5071 13185 5097 13186
rect 4487 12975 4521 13167
rect 5033 13151 5097 13185
rect 5873 13302 5885 13336
rect 5919 13302 5931 13336
rect 5873 13243 5931 13302
rect 5965 13296 6086 13407
rect 6121 13356 6217 13373
rect 6155 13334 6217 13356
rect 6121 13305 6146 13322
rect 6182 13305 6217 13334
rect 6251 13365 6302 13407
rect 6251 13331 6255 13365
rect 6289 13331 6302 13365
rect 6251 13298 6302 13331
rect 6336 13351 6391 13373
rect 6844 13365 6892 13417
rect 6928 13451 6984 13467
rect 6928 13417 6942 13451
rect 6976 13417 6984 13451
rect 6928 13401 6984 13417
rect 7030 13451 7073 13467
rect 7030 13417 7038 13451
rect 7072 13417 7073 13451
rect 7030 13365 7073 13417
rect 7107 13443 7230 13477
rect 7107 13409 7123 13443
rect 7157 13409 7230 13443
rect 7107 13399 7230 13409
rect 7267 13493 7325 13510
rect 11689 13505 11760 13524
rect 7267 13459 7279 13493
rect 7313 13459 7325 13493
rect 11794 13471 11828 13651
rect 11862 13608 11915 13617
rect 11862 13601 11878 13608
rect 11912 13574 11915 13608
rect 11896 13567 11915 13574
rect 11862 13505 11915 13567
rect 11965 13601 11999 13651
rect 11965 13551 11999 13567
rect 12033 13517 12096 13721
rect 12135 13808 12193 13879
rect 12606 13861 12676 13908
rect 13001 13875 13035 13909
rect 12713 13841 13035 13875
rect 13089 13862 13123 14009
rect 13157 14166 13215 14237
rect 13157 14132 13169 14166
rect 13203 14132 13215 14166
rect 13157 14073 13215 14132
rect 13157 14039 13169 14073
rect 13203 14039 13215 14073
rect 13157 14004 13215 14039
rect 13069 13845 13123 13862
rect 12135 13774 12147 13808
rect 12181 13774 12193 13808
rect 12135 13715 12193 13774
rect 12607 13793 12623 13827
rect 12657 13793 12673 13827
rect 12607 13727 12673 13793
rect 12713 13821 12747 13841
rect 12887 13821 12921 13841
rect 12713 13771 12747 13787
rect 12787 13773 12803 13807
rect 12837 13773 12853 13807
rect 12787 13727 12853 13773
rect 13103 13811 13123 13845
rect 12887 13771 12921 13787
rect 12955 13773 12981 13807
rect 13015 13773 13031 13807
rect 13069 13793 13123 13811
rect 13157 13855 13215 13872
rect 13157 13821 13169 13855
rect 13203 13821 13215 13855
rect 12955 13727 13031 13773
rect 13157 13727 13215 13821
rect 12135 13681 12147 13715
rect 12181 13681 12193 13715
rect 12588 13693 12617 13727
rect 12651 13693 12709 13727
rect 12743 13693 12801 13727
rect 12835 13693 12893 13727
rect 12927 13693 12985 13727
rect 13019 13693 13077 13727
rect 13111 13693 13169 13727
rect 13203 13693 13232 13727
rect 12135 13646 12193 13681
rect 11973 13515 12096 13517
rect 11973 13481 11989 13515
rect 12023 13481 12096 13515
rect 7267 13365 7325 13459
rect 11710 13455 11758 13471
rect 10722 13411 10751 13445
rect 10785 13411 10843 13445
rect 10877 13411 10935 13445
rect 10969 13411 11027 13445
rect 11061 13411 11119 13445
rect 11153 13411 11211 13445
rect 11245 13411 11274 13445
rect 11710 13421 11724 13455
rect 6336 13317 6339 13351
rect 6373 13317 6391 13351
rect 6794 13331 6823 13365
rect 6857 13331 6915 13365
rect 6949 13331 7007 13365
rect 7041 13331 7099 13365
rect 7133 13331 7191 13365
rect 7225 13331 7279 13365
rect 7313 13331 7342 13365
rect 9244 13341 9273 13375
rect 9307 13341 9365 13375
rect 9399 13341 9457 13375
rect 9491 13341 9549 13375
rect 9583 13341 9641 13375
rect 9675 13341 9733 13375
rect 9767 13341 9825 13375
rect 9859 13341 9917 13375
rect 9951 13341 9980 13375
rect 5965 13276 6088 13296
rect 5873 13209 5885 13243
rect 5919 13209 5931 13243
rect 6051 13271 6088 13276
rect 6336 13283 6391 13317
rect 6051 13256 6117 13271
rect 5873 13174 5931 13209
rect 5965 13226 6017 13242
rect 5965 13192 5983 13226
rect 6051 13222 6067 13256
rect 6101 13222 6117 13256
rect 6151 13237 6302 13257
rect 6151 13207 6160 13237
rect 6148 13203 6160 13207
rect 6194 13203 6302 13237
rect 6336 13249 6339 13283
rect 6373 13278 6391 13283
rect 6336 13240 6342 13249
rect 6380 13240 6391 13278
rect 6336 13233 6391 13240
rect 6148 13200 6302 13203
rect 6145 13198 6302 13200
rect 6144 13195 6323 13198
rect 6140 13192 6323 13195
rect 4555 13099 4816 13133
rect 5033 13117 5037 13151
rect 5071 13117 5097 13151
rect 5965 13152 6017 13192
rect 6136 13190 6323 13192
rect 6131 13188 6323 13190
rect 6117 13182 6323 13188
rect 6113 13176 6323 13182
rect 6109 13170 6323 13176
rect 6103 13165 6323 13170
rect 6096 13158 6323 13165
rect 6090 13157 6323 13158
rect 6090 13156 6168 13157
rect 6090 13154 6163 13156
rect 6090 13153 6160 13154
rect 6090 13152 6157 13153
rect 5965 13151 6157 13152
rect 5965 13149 6155 13151
rect 5965 13148 6153 13149
rect 5965 13146 6151 13148
rect 5965 13144 6150 13146
rect 5965 13143 6149 13144
rect 5965 13140 6147 13143
rect 5965 13137 6146 13140
rect 5965 13132 6144 13137
rect 5965 13118 6143 13132
rect 6277 13129 6323 13157
rect 4555 13060 4604 13099
rect 4555 13059 4556 13060
rect 4590 13026 4604 13060
rect 4589 13025 4604 13026
rect 4638 13062 4748 13065
rect 4638 13059 4676 13062
rect 4638 13025 4672 13059
rect 4710 13028 4748 13062
rect 4706 13025 4748 13028
rect 4782 13059 4816 13099
rect 4971 13083 5097 13117
rect 5965 13083 6075 13084
rect 4891 13059 4937 13075
rect 4782 13025 4807 13059
rect 4841 13025 4857 13059
rect 4891 13025 4903 13059
rect 4555 13009 4604 13025
rect 4891 12975 4937 13025
rect 4395 12955 4453 12972
rect 4395 12921 4407 12955
rect 4441 12921 4453 12955
rect 4487 12941 4937 12975
rect 4395 12827 4453 12921
rect 4597 12927 4631 12941
rect 4497 12871 4513 12905
rect 4547 12871 4563 12905
rect 4971 12907 5005 13083
rect 5965 13049 5983 13083
rect 6017 13060 6075 13083
rect 5873 13025 5931 13042
rect 4597 12877 4631 12893
rect 4497 12827 4563 12871
rect 4665 12871 4681 12905
rect 4715 12871 4731 12905
rect 4814 12873 4849 12907
rect 4883 12873 4949 12907
rect 4983 12873 5005 12907
rect 5039 12978 5097 12994
rect 5073 12944 5097 12978
rect 5039 12910 5097 12944
rect 5073 12876 5097 12910
rect 5873 12991 5885 13025
rect 5919 12991 5931 13025
rect 5965 13026 5994 13049
rect 6028 13026 6075 13060
rect 5965 13007 6075 13026
rect 5873 12897 5931 12991
rect 6109 12973 6143 13118
rect 5965 12939 5983 12973
rect 6017 12939 6143 12973
rect 6177 13089 6193 13123
rect 6227 13089 6243 13123
rect 6177 13066 6243 13089
rect 6277 13095 6289 13129
rect 6277 13078 6323 13095
rect 6177 13032 6196 13066
rect 6232 13038 6243 13066
rect 6177 12941 6221 13032
rect 6357 13027 6391 13233
rect 9261 13270 9319 13341
rect 9261 13236 9273 13270
rect 9307 13236 9319 13270
rect 9261 13177 9319 13236
rect 9261 13143 9273 13177
rect 9307 13143 9319 13177
rect 9261 13108 9319 13143
rect 9353 13299 9429 13307
rect 9353 13265 9379 13299
rect 9413 13265 9429 13299
rect 9353 13231 9429 13265
rect 9353 13197 9379 13231
rect 9413 13197 9429 13231
rect 9353 13171 9429 13197
rect 9547 13289 9581 13341
rect 9547 13221 9581 13255
rect 9547 13171 9581 13187
rect 9615 13289 9681 13307
rect 9615 13255 9631 13289
rect 9665 13255 9681 13289
rect 9615 13221 9681 13255
rect 9715 13289 9749 13341
rect 10739 13340 10797 13411
rect 9715 13239 9749 13255
rect 9783 13289 9863 13307
rect 9783 13255 9819 13289
rect 9853 13255 9863 13289
rect 9615 13187 9631 13221
rect 9665 13205 9681 13221
rect 9783 13221 9863 13255
rect 9783 13205 9819 13221
rect 9665 13187 9819 13205
rect 9853 13187 9863 13221
rect 9615 13171 9863 13187
rect 9899 13291 9963 13307
rect 9899 13257 9903 13291
rect 9937 13257 9963 13291
rect 9899 13224 9963 13257
rect 9899 13223 9914 13224
rect 9899 13189 9903 13223
rect 9948 13190 9963 13224
rect 9937 13189 9963 13190
rect 6255 12989 6305 13005
rect 6289 12955 6305 12989
rect 6255 12897 6305 12955
rect 6339 12999 6391 13027
rect 6373 12965 6391 12999
rect 9353 12979 9387 13171
rect 9899 13155 9963 13189
rect 10739 13306 10751 13340
rect 10785 13306 10797 13340
rect 10739 13247 10797 13306
rect 10831 13300 10952 13411
rect 10987 13360 11083 13377
rect 11021 13338 11083 13360
rect 10987 13309 11012 13326
rect 11048 13309 11083 13338
rect 11117 13369 11168 13411
rect 11117 13335 11121 13369
rect 11155 13335 11168 13369
rect 11117 13302 11168 13335
rect 11202 13355 11257 13377
rect 11710 13369 11758 13421
rect 11794 13455 11850 13471
rect 11794 13421 11808 13455
rect 11842 13421 11850 13455
rect 11794 13405 11850 13421
rect 11896 13455 11939 13471
rect 11896 13421 11904 13455
rect 11938 13421 11939 13455
rect 11896 13369 11939 13421
rect 11973 13447 12096 13481
rect 11973 13413 11989 13447
rect 12023 13413 12096 13447
rect 11973 13403 12096 13413
rect 12135 13497 12193 13514
rect 12135 13463 12147 13497
rect 12181 13463 12193 13497
rect 12135 13369 12193 13463
rect 11202 13321 11205 13355
rect 11239 13321 11257 13355
rect 11660 13335 11689 13369
rect 11723 13335 11781 13369
rect 11815 13335 11873 13369
rect 11907 13335 11965 13369
rect 11999 13335 12057 13369
rect 12091 13335 12147 13369
rect 12181 13335 12210 13369
rect 10831 13280 10954 13300
rect 10739 13213 10751 13247
rect 10785 13213 10797 13247
rect 10917 13275 10954 13280
rect 11202 13287 11257 13321
rect 10917 13260 10983 13275
rect 10739 13178 10797 13213
rect 10831 13230 10883 13246
rect 10831 13196 10849 13230
rect 10917 13226 10933 13260
rect 10967 13226 10983 13260
rect 11017 13241 11168 13261
rect 11017 13211 11026 13241
rect 11014 13207 11026 13211
rect 11060 13207 11168 13241
rect 11202 13253 11205 13287
rect 11239 13282 11257 13287
rect 11202 13244 11208 13253
rect 11246 13244 11257 13282
rect 11202 13237 11257 13244
rect 11014 13204 11168 13207
rect 11011 13202 11168 13204
rect 11010 13199 11189 13202
rect 11006 13196 11189 13199
rect 9421 13103 9682 13137
rect 9899 13121 9903 13155
rect 9937 13121 9963 13155
rect 10831 13156 10883 13196
rect 11002 13194 11189 13196
rect 10997 13192 11189 13194
rect 10983 13186 11189 13192
rect 10979 13180 11189 13186
rect 10975 13174 11189 13180
rect 10969 13169 11189 13174
rect 10962 13162 11189 13169
rect 10956 13161 11189 13162
rect 10956 13160 11034 13161
rect 10956 13158 11029 13160
rect 10956 13157 11026 13158
rect 10956 13156 11023 13157
rect 10831 13155 11023 13156
rect 10831 13153 11021 13155
rect 10831 13152 11019 13153
rect 10831 13150 11017 13152
rect 10831 13148 11016 13150
rect 10831 13147 11015 13148
rect 10831 13144 11013 13147
rect 10831 13141 11012 13144
rect 10831 13136 11010 13141
rect 10831 13122 11009 13136
rect 11143 13133 11189 13161
rect 9421 13064 9470 13103
rect 9421 13063 9422 13064
rect 9456 13030 9470 13064
rect 9455 13029 9470 13030
rect 9504 13066 9614 13069
rect 9504 13063 9542 13066
rect 9504 13029 9538 13063
rect 9576 13032 9614 13066
rect 9572 13029 9614 13032
rect 9648 13063 9682 13103
rect 9837 13087 9963 13121
rect 10831 13087 10941 13088
rect 9757 13063 9803 13079
rect 9648 13029 9673 13063
rect 9707 13029 9723 13063
rect 9757 13029 9769 13063
rect 9421 13013 9470 13029
rect 9757 12979 9803 13029
rect 6339 12931 6391 12965
rect 9261 12959 9319 12976
rect 9261 12925 9273 12959
rect 9307 12925 9319 12959
rect 9353 12945 9803 12979
rect 4665 12827 4731 12871
rect 5039 12827 5097 12876
rect 5856 12863 5885 12897
rect 5919 12863 5977 12897
rect 6011 12863 6069 12897
rect 6103 12863 6161 12897
rect 6195 12863 6253 12897
rect 6287 12863 6345 12897
rect 6379 12863 6408 12897
rect 9261 12831 9319 12925
rect 9463 12931 9497 12945
rect 9363 12875 9379 12909
rect 9413 12875 9429 12909
rect 9837 12911 9871 13087
rect 10831 13053 10849 13087
rect 10883 13064 10941 13087
rect 10739 13029 10797 13046
rect 9463 12881 9497 12897
rect 9363 12831 9429 12875
rect 9531 12875 9547 12909
rect 9581 12875 9597 12909
rect 9680 12877 9715 12911
rect 9749 12877 9815 12911
rect 9849 12877 9871 12911
rect 9905 12982 9963 12998
rect 9939 12948 9963 12982
rect 9905 12914 9963 12948
rect 9939 12880 9963 12914
rect 10739 12995 10751 13029
rect 10785 12995 10797 13029
rect 10831 13030 10860 13053
rect 10894 13030 10941 13064
rect 10831 13011 10941 13030
rect 10739 12901 10797 12995
rect 10975 12977 11009 13122
rect 10831 12943 10849 12977
rect 10883 12943 11009 12977
rect 11043 13093 11059 13127
rect 11093 13093 11109 13127
rect 11043 13070 11109 13093
rect 11143 13099 11155 13133
rect 11143 13082 11189 13099
rect 11043 13036 11062 13070
rect 11098 13042 11109 13070
rect 11043 12945 11087 13036
rect 11223 13031 11257 13237
rect 11121 12993 11171 13009
rect 11155 12959 11171 12993
rect 11121 12901 11171 12959
rect 11205 13003 11257 13031
rect 11239 12969 11257 13003
rect 11205 12935 11257 12969
rect 9531 12831 9597 12875
rect 9905 12831 9963 12880
rect 10722 12867 10751 12901
rect 10785 12867 10843 12901
rect 10877 12867 10935 12901
rect 10969 12867 11027 12901
rect 11061 12867 11119 12901
rect 11153 12867 11211 12901
rect 11245 12867 11274 12901
rect 4378 12793 4407 12827
rect 4441 12793 4499 12827
rect 4533 12793 4591 12827
rect 4625 12793 4683 12827
rect 4717 12793 4775 12827
rect 4809 12793 4867 12827
rect 4901 12793 4959 12827
rect 4993 12793 5051 12827
rect 5085 12793 5114 12827
rect 9244 12797 9273 12831
rect 9307 12797 9365 12831
rect 9399 12797 9457 12831
rect 9491 12797 9549 12831
rect 9583 12797 9641 12831
rect 9675 12797 9733 12831
rect 9767 12797 9825 12831
rect 9859 12797 9917 12831
rect 9951 12797 9980 12831
rect 4478 12593 4507 12627
rect 4541 12593 4597 12627
rect 4631 12593 4689 12627
rect 4723 12593 4781 12627
rect 4815 12593 4873 12627
rect 4907 12593 4965 12627
rect 4999 12593 5028 12627
rect 9342 12597 9371 12631
rect 9405 12597 9463 12631
rect 9497 12597 9555 12631
rect 9589 12597 9647 12631
rect 9681 12597 9739 12631
rect 9773 12597 9831 12631
rect 9865 12597 9894 12631
rect 4495 12522 4553 12593
rect 4495 12488 4507 12522
rect 4541 12488 4553 12522
rect 4495 12429 4553 12488
rect 4625 12509 4681 12593
rect 4815 12551 4881 12593
rect 4625 12475 4639 12509
rect 4673 12475 4681 12509
rect 4625 12459 4681 12475
rect 4715 12509 4775 12525
rect 4715 12475 4723 12509
rect 4757 12475 4775 12509
rect 4495 12395 4507 12429
rect 4541 12395 4553 12429
rect 4715 12415 4775 12475
rect 4815 12517 4831 12551
rect 4865 12517 4881 12551
rect 4815 12483 4881 12517
rect 4815 12449 4831 12483
rect 4865 12449 4881 12483
rect 4919 12551 5011 12559
rect 4919 12517 4935 12551
rect 4969 12517 5011 12551
rect 4919 12483 5011 12517
rect 4919 12449 4935 12483
rect 4969 12449 5011 12483
rect 4495 12360 4553 12395
rect 4588 12338 4641 12403
rect 4715 12381 4903 12415
rect 4588 12298 4590 12338
rect 4632 12331 4641 12338
rect 4869 12331 4903 12381
rect 4961 12370 5011 12449
rect 9359 12526 9417 12597
rect 9359 12492 9371 12526
rect 9405 12492 9417 12526
rect 9359 12433 9417 12492
rect 9491 12513 9547 12597
rect 9681 12555 9747 12597
rect 9491 12479 9505 12513
rect 9539 12479 9547 12513
rect 9491 12463 9547 12479
rect 9581 12513 9641 12529
rect 9581 12479 9589 12513
rect 9623 12479 9641 12513
rect 5852 12387 5881 12421
rect 5915 12387 5973 12421
rect 6007 12387 6065 12421
rect 6099 12387 6157 12421
rect 6191 12387 6249 12421
rect 6283 12387 6341 12421
rect 6375 12387 6404 12421
rect 9359 12399 9371 12433
rect 9405 12399 9417 12433
rect 9581 12419 9641 12479
rect 9681 12521 9697 12555
rect 9731 12521 9747 12555
rect 9681 12487 9747 12521
rect 9681 12453 9697 12487
rect 9731 12453 9747 12487
rect 9785 12555 9877 12563
rect 9785 12521 9801 12555
rect 9835 12521 9877 12555
rect 9785 12487 9877 12521
rect 9785 12453 9801 12487
rect 9835 12453 9877 12487
rect 4961 12336 4970 12370
rect 5006 12336 5011 12370
rect 4632 12315 4723 12331
rect 4632 12298 4642 12315
rect 4588 12281 4642 12298
rect 4676 12281 4723 12315
rect 4767 12328 4835 12331
rect 4767 12288 4780 12328
rect 4822 12288 4835 12328
rect 4767 12281 4783 12288
rect 4817 12281 4835 12288
rect 4869 12315 4927 12331
rect 4869 12281 4891 12315
rect 4925 12281 4927 12315
rect 4869 12265 4927 12281
rect 4869 12247 4903 12265
rect 4495 12211 4553 12228
rect 4495 12177 4507 12211
rect 4541 12177 4553 12211
rect 4495 12083 4553 12177
rect 4625 12209 4903 12247
rect 4625 12187 4691 12209
rect 4625 12153 4639 12187
rect 4673 12153 4691 12187
rect 4961 12175 5011 12336
rect 4625 12137 4691 12153
rect 4815 12159 4865 12175
rect 4815 12125 4831 12159
rect 4815 12083 4865 12125
rect 4899 12159 5011 12175
rect 4899 12125 4915 12159
rect 4949 12125 5011 12159
rect 5869 12316 5927 12387
rect 5869 12282 5881 12316
rect 5915 12282 5927 12316
rect 5869 12223 5927 12282
rect 6001 12303 6057 12387
rect 6191 12345 6257 12387
rect 9359 12364 9417 12399
rect 6001 12269 6015 12303
rect 6049 12269 6057 12303
rect 6001 12253 6057 12269
rect 6091 12303 6151 12319
rect 6091 12269 6099 12303
rect 6133 12269 6151 12303
rect 5869 12189 5881 12223
rect 5915 12189 5927 12223
rect 6091 12209 6151 12269
rect 6191 12311 6207 12345
rect 6241 12311 6257 12345
rect 6191 12277 6257 12311
rect 6191 12243 6207 12277
rect 6241 12243 6257 12277
rect 6295 12345 6387 12353
rect 6295 12311 6311 12345
rect 6345 12311 6387 12345
rect 6295 12277 6387 12311
rect 9454 12342 9507 12407
rect 9581 12385 9769 12419
rect 9454 12302 9456 12342
rect 9498 12335 9507 12342
rect 9735 12335 9769 12385
rect 9827 12374 9877 12453
rect 10718 12391 10747 12425
rect 10781 12391 10839 12425
rect 10873 12391 10931 12425
rect 10965 12391 11023 12425
rect 11057 12391 11115 12425
rect 11149 12391 11207 12425
rect 11241 12391 11270 12425
rect 9827 12340 9836 12374
rect 9872 12340 9877 12374
rect 9498 12319 9589 12335
rect 9498 12302 9508 12319
rect 9454 12285 9508 12302
rect 9542 12285 9589 12319
rect 9633 12332 9701 12335
rect 9633 12292 9646 12332
rect 9688 12292 9701 12332
rect 9633 12285 9649 12292
rect 9683 12285 9701 12292
rect 9735 12319 9793 12335
rect 9735 12285 9757 12319
rect 9791 12285 9793 12319
rect 6295 12243 6311 12277
rect 6345 12243 6387 12277
rect 9735 12269 9793 12285
rect 9735 12251 9769 12269
rect 5869 12154 5927 12189
rect 4899 12117 5011 12125
rect 5964 12125 6017 12197
rect 6091 12175 6279 12209
rect 6245 12125 6279 12175
rect 6337 12196 6387 12243
rect 6337 12162 6346 12196
rect 6380 12162 6387 12196
rect 5964 12112 6099 12125
rect 4478 12049 4507 12083
rect 4541 12049 4597 12083
rect 4631 12049 4689 12083
rect 4723 12049 4781 12083
rect 4815 12049 4873 12083
rect 4907 12049 4965 12083
rect 4999 12049 5028 12083
rect 5964 12075 6018 12112
rect 6054 12078 6099 12112
rect 6052 12075 6099 12078
rect 6143 12110 6211 12125
rect 6143 12076 6158 12110
rect 6194 12076 6211 12110
rect 6143 12075 6159 12076
rect 6193 12075 6211 12076
rect 6245 12109 6303 12125
rect 6245 12075 6267 12109
rect 6301 12075 6303 12109
rect 6245 12059 6303 12075
rect 6245 12041 6279 12059
rect 5869 12005 5927 12022
rect 5869 11971 5881 12005
rect 5915 11971 5927 12005
rect 5869 11877 5927 11971
rect 6001 12003 6279 12041
rect 6001 11981 6067 12003
rect 6001 11947 6015 11981
rect 6049 11947 6067 11981
rect 6337 11969 6387 12162
rect 9359 12215 9417 12232
rect 9359 12181 9371 12215
rect 9405 12181 9417 12215
rect 9359 12087 9417 12181
rect 9491 12213 9769 12251
rect 9491 12191 9557 12213
rect 9491 12157 9505 12191
rect 9539 12157 9557 12191
rect 9827 12179 9877 12340
rect 9491 12141 9557 12157
rect 9681 12163 9731 12179
rect 9681 12129 9697 12163
rect 9681 12087 9731 12129
rect 9765 12163 9877 12179
rect 9765 12129 9781 12163
rect 9815 12129 9877 12163
rect 10735 12320 10793 12391
rect 10735 12286 10747 12320
rect 10781 12286 10793 12320
rect 10735 12227 10793 12286
rect 10867 12307 10923 12391
rect 11057 12349 11123 12391
rect 10867 12273 10881 12307
rect 10915 12273 10923 12307
rect 10867 12257 10923 12273
rect 10957 12307 11017 12323
rect 10957 12273 10965 12307
rect 10999 12273 11017 12307
rect 10735 12193 10747 12227
rect 10781 12193 10793 12227
rect 10957 12213 11017 12273
rect 11057 12315 11073 12349
rect 11107 12315 11123 12349
rect 11057 12281 11123 12315
rect 11057 12247 11073 12281
rect 11107 12247 11123 12281
rect 11161 12349 11253 12357
rect 11161 12315 11177 12349
rect 11211 12315 11253 12349
rect 11161 12281 11253 12315
rect 11161 12247 11177 12281
rect 11211 12247 11253 12281
rect 10735 12158 10793 12193
rect 9765 12121 9877 12129
rect 10830 12129 10883 12201
rect 10957 12179 11145 12213
rect 11111 12129 11145 12179
rect 11203 12200 11253 12247
rect 11203 12166 11212 12200
rect 11246 12166 11253 12200
rect 10830 12116 10965 12129
rect 9342 12053 9371 12087
rect 9405 12053 9463 12087
rect 9497 12053 9555 12087
rect 9589 12053 9647 12087
rect 9681 12053 9739 12087
rect 9773 12053 9831 12087
rect 9865 12053 9894 12087
rect 10830 12079 10884 12116
rect 10920 12082 10965 12116
rect 10918 12079 10965 12082
rect 11009 12114 11077 12129
rect 11009 12080 11024 12114
rect 11060 12080 11077 12114
rect 11009 12079 11025 12080
rect 11059 12079 11077 12080
rect 11111 12113 11169 12129
rect 11111 12079 11133 12113
rect 11167 12079 11169 12113
rect 11111 12063 11169 12079
rect 11111 12045 11145 12063
rect 6001 11931 6067 11947
rect 6191 11953 6241 11969
rect 6191 11919 6207 11953
rect 6191 11877 6241 11919
rect 6275 11953 6387 11969
rect 6275 11919 6291 11953
rect 6325 11919 6387 11953
rect 6275 11911 6387 11919
rect 10735 12009 10793 12026
rect 10735 11975 10747 12009
rect 10781 11975 10793 12009
rect 10735 11881 10793 11975
rect 10867 12007 11145 12045
rect 10867 11985 10933 12007
rect 10867 11951 10881 11985
rect 10915 11951 10933 11985
rect 11203 11973 11253 12166
rect 10867 11935 10933 11951
rect 11057 11957 11107 11973
rect 11057 11923 11073 11957
rect 11057 11881 11107 11923
rect 11141 11957 11253 11973
rect 11141 11923 11157 11957
rect 11191 11923 11253 11957
rect 11141 11915 11253 11923
rect 5852 11843 5881 11877
rect 5915 11843 5973 11877
rect 6007 11843 6065 11877
rect 6099 11843 6157 11877
rect 6191 11843 6249 11877
rect 6283 11843 6341 11877
rect 6375 11843 6404 11877
rect 10718 11847 10747 11881
rect 10781 11847 10839 11881
rect 10873 11847 10931 11881
rect 10965 11847 11023 11881
rect 11057 11847 11115 11881
rect 11149 11847 11207 11881
rect 11241 11847 11270 11881
rect 4388 11773 4417 11807
rect 4451 11773 4509 11807
rect 4543 11773 4601 11807
rect 4635 11773 4693 11807
rect 4727 11773 4785 11807
rect 4819 11773 4877 11807
rect 4911 11773 4969 11807
rect 5003 11773 5061 11807
rect 5095 11773 5124 11807
rect 9254 11777 9283 11811
rect 9317 11777 9375 11811
rect 9409 11777 9467 11811
rect 9501 11777 9559 11811
rect 9593 11777 9651 11811
rect 9685 11777 9743 11811
rect 9777 11777 9835 11811
rect 9869 11777 9927 11811
rect 9961 11777 9990 11811
rect 4405 11702 4463 11773
rect 4405 11668 4417 11702
rect 4451 11668 4463 11702
rect 4405 11609 4463 11668
rect 4405 11575 4417 11609
rect 4451 11575 4463 11609
rect 4405 11540 4463 11575
rect 4497 11731 4573 11739
rect 4497 11697 4523 11731
rect 4557 11697 4573 11731
rect 4497 11663 4573 11697
rect 4497 11629 4523 11663
rect 4557 11629 4573 11663
rect 4497 11603 4573 11629
rect 4691 11721 4725 11773
rect 4691 11653 4725 11687
rect 4691 11603 4725 11619
rect 4759 11721 4825 11739
rect 4759 11687 4775 11721
rect 4809 11687 4825 11721
rect 4759 11653 4825 11687
rect 4859 11721 4893 11773
rect 4859 11671 4893 11687
rect 4927 11721 5007 11739
rect 4927 11687 4963 11721
rect 4997 11687 5007 11721
rect 4759 11619 4775 11653
rect 4809 11637 4825 11653
rect 4927 11653 5007 11687
rect 4927 11637 4963 11653
rect 4809 11619 4963 11637
rect 4997 11619 5007 11653
rect 4759 11603 5007 11619
rect 5043 11723 5107 11739
rect 5043 11689 5047 11723
rect 5081 11689 5107 11723
rect 5043 11656 5107 11689
rect 5043 11655 5048 11656
rect 5043 11621 5047 11655
rect 5084 11622 5107 11656
rect 5081 11621 5107 11622
rect 4497 11411 4531 11603
rect 5043 11587 5107 11621
rect 4565 11535 4826 11569
rect 5043 11553 5047 11587
rect 5081 11553 5107 11587
rect 4565 11496 4614 11535
rect 4565 11495 4566 11496
rect 4600 11462 4614 11496
rect 4599 11461 4614 11462
rect 4648 11498 4758 11501
rect 4648 11495 4686 11498
rect 4648 11461 4682 11495
rect 4720 11464 4758 11498
rect 4716 11461 4758 11464
rect 4792 11495 4826 11535
rect 4981 11519 5107 11553
rect 9271 11706 9329 11777
rect 9271 11672 9283 11706
rect 9317 11672 9329 11706
rect 9271 11613 9329 11672
rect 9271 11579 9283 11613
rect 9317 11579 9329 11613
rect 9271 11544 9329 11579
rect 9363 11735 9439 11743
rect 9363 11701 9389 11735
rect 9423 11701 9439 11735
rect 9363 11667 9439 11701
rect 9363 11633 9389 11667
rect 9423 11633 9439 11667
rect 9363 11607 9439 11633
rect 9557 11725 9591 11777
rect 9557 11657 9591 11691
rect 9557 11607 9591 11623
rect 9625 11725 9691 11743
rect 9625 11691 9641 11725
rect 9675 11691 9691 11725
rect 9625 11657 9691 11691
rect 9725 11725 9759 11777
rect 9725 11675 9759 11691
rect 9793 11725 9873 11743
rect 9793 11691 9829 11725
rect 9863 11691 9873 11725
rect 9625 11623 9641 11657
rect 9675 11641 9691 11657
rect 9793 11657 9873 11691
rect 9793 11641 9829 11657
rect 9675 11623 9829 11641
rect 9863 11623 9873 11657
rect 9625 11607 9873 11623
rect 9909 11727 9973 11743
rect 9909 11693 9913 11727
rect 9947 11693 9973 11727
rect 9909 11660 9973 11693
rect 9909 11659 9914 11660
rect 9909 11625 9913 11659
rect 9950 11626 9973 11660
rect 9947 11625 9973 11626
rect 4901 11495 4947 11511
rect 4792 11461 4817 11495
rect 4851 11461 4867 11495
rect 4901 11461 4913 11495
rect 4565 11445 4614 11461
rect 4901 11411 4947 11461
rect 4405 11391 4463 11408
rect 4405 11357 4417 11391
rect 4451 11357 4463 11391
rect 4497 11377 4947 11411
rect 4405 11263 4463 11357
rect 4607 11363 4641 11377
rect 4507 11307 4523 11341
rect 4557 11307 4573 11341
rect 4981 11343 5015 11519
rect 4607 11313 4641 11329
rect 4507 11263 4573 11307
rect 4675 11307 4691 11341
rect 4725 11307 4741 11341
rect 4824 11309 4859 11343
rect 4893 11309 4959 11343
rect 4993 11309 5015 11343
rect 5049 11414 5107 11430
rect 5083 11380 5107 11414
rect 9363 11415 9397 11607
rect 9909 11591 9973 11625
rect 9431 11539 9692 11573
rect 9909 11557 9913 11591
rect 9947 11557 9973 11591
rect 9431 11500 9480 11539
rect 9431 11499 9432 11500
rect 9466 11466 9480 11500
rect 9465 11465 9480 11466
rect 9514 11502 9624 11505
rect 9514 11499 9552 11502
rect 9514 11465 9548 11499
rect 9586 11468 9624 11502
rect 9582 11465 9624 11468
rect 9658 11499 9692 11539
rect 9847 11523 9973 11557
rect 9767 11499 9813 11515
rect 9658 11465 9683 11499
rect 9717 11465 9733 11499
rect 9767 11465 9779 11499
rect 9431 11449 9480 11465
rect 9767 11415 9813 11465
rect 5049 11346 5107 11380
rect 5083 11312 5107 11346
rect 4675 11263 4741 11307
rect 5049 11263 5107 11312
rect 9271 11395 9329 11412
rect 9271 11361 9283 11395
rect 9317 11361 9329 11395
rect 9363 11381 9813 11415
rect 9271 11267 9329 11361
rect 9473 11367 9507 11381
rect 9373 11311 9389 11345
rect 9423 11311 9439 11345
rect 9847 11347 9881 11523
rect 9473 11317 9507 11333
rect 9373 11267 9439 11311
rect 9541 11311 9557 11345
rect 9591 11311 9607 11345
rect 9690 11313 9725 11347
rect 9759 11313 9825 11347
rect 9859 11313 9881 11347
rect 9915 11418 9973 11434
rect 9949 11384 9973 11418
rect 9915 11350 9973 11384
rect 9949 11316 9973 11350
rect 9541 11267 9607 11311
rect 9915 11267 9973 11316
rect 4388 11229 4417 11263
rect 4451 11229 4509 11263
rect 4543 11229 4601 11263
rect 4635 11229 4693 11263
rect 4727 11229 4785 11263
rect 4819 11229 4877 11263
rect 4911 11229 4969 11263
rect 5003 11229 5061 11263
rect 5095 11229 5124 11263
rect 9254 11233 9283 11267
rect 9317 11233 9375 11267
rect 9409 11233 9467 11267
rect 9501 11233 9559 11267
rect 9593 11233 9651 11267
rect 9685 11233 9743 11267
rect 9777 11233 9835 11267
rect 9869 11233 9927 11267
rect 9961 11233 9990 11267
rect 4486 11029 4515 11063
rect 4549 11029 4607 11063
rect 4641 11029 4699 11063
rect 4733 11029 4791 11063
rect 4825 11029 4883 11063
rect 4917 11029 4975 11063
rect 5009 11029 5038 11063
rect 9352 11033 9381 11067
rect 9415 11033 9473 11067
rect 9507 11033 9565 11067
rect 9599 11033 9657 11067
rect 9691 11033 9749 11067
rect 9783 11033 9841 11067
rect 9875 11033 9904 11067
rect 4503 10958 4561 11029
rect 4503 10924 4515 10958
rect 4549 10924 4561 10958
rect 4503 10865 4561 10924
rect 4635 10945 4691 11029
rect 4825 10987 4891 11029
rect 4635 10911 4649 10945
rect 4683 10911 4691 10945
rect 4635 10895 4691 10911
rect 4725 10945 4785 10961
rect 4725 10911 4733 10945
rect 4767 10911 4785 10945
rect 4503 10831 4515 10865
rect 4549 10831 4561 10865
rect 4725 10851 4785 10911
rect 4825 10953 4841 10987
rect 4875 10953 4891 10987
rect 4825 10919 4891 10953
rect 4825 10885 4841 10919
rect 4875 10885 4891 10919
rect 4929 10987 5021 10995
rect 4929 10953 4945 10987
rect 4979 10953 5021 10987
rect 4929 10919 5021 10953
rect 4929 10885 4945 10919
rect 4979 10885 5021 10919
rect 4503 10796 4561 10831
rect 4598 10774 4651 10839
rect 4725 10817 4913 10851
rect 4598 10734 4600 10774
rect 4642 10767 4651 10774
rect 4879 10767 4913 10817
rect 4642 10751 4733 10767
rect 4642 10734 4652 10751
rect 4598 10717 4652 10734
rect 4686 10717 4733 10751
rect 4777 10764 4845 10767
rect 4777 10724 4790 10764
rect 4832 10724 4845 10764
rect 4777 10717 4793 10724
rect 4827 10717 4845 10724
rect 4879 10751 4937 10767
rect 4879 10717 4901 10751
rect 4935 10717 4937 10751
rect 4879 10701 4937 10717
rect 4971 10730 5021 10885
rect 9369 10962 9427 11033
rect 9369 10928 9381 10962
rect 9415 10928 9427 10962
rect 9369 10869 9427 10928
rect 9501 10949 9557 11033
rect 9691 10991 9757 11033
rect 9501 10915 9515 10949
rect 9549 10915 9557 10949
rect 9501 10899 9557 10915
rect 9591 10949 9651 10965
rect 9591 10915 9599 10949
rect 9633 10915 9651 10949
rect 9369 10835 9381 10869
rect 9415 10835 9427 10869
rect 9591 10855 9651 10915
rect 9691 10957 9707 10991
rect 9741 10957 9757 10991
rect 9691 10923 9757 10957
rect 9691 10889 9707 10923
rect 9741 10889 9757 10923
rect 9795 10991 9887 10999
rect 9795 10957 9811 10991
rect 9845 10957 9887 10991
rect 9795 10923 9887 10957
rect 9795 10889 9811 10923
rect 9845 10889 9887 10923
rect 9369 10800 9427 10835
rect 4879 10683 4913 10701
rect 4503 10647 4561 10664
rect 4503 10613 4515 10647
rect 4549 10613 4561 10647
rect 4503 10519 4561 10613
rect 4635 10645 4913 10683
rect 4971 10694 4982 10730
rect 5016 10694 5021 10730
rect 9464 10778 9517 10843
rect 9591 10821 9779 10855
rect 9464 10738 9466 10778
rect 9508 10771 9517 10778
rect 9745 10771 9779 10821
rect 9508 10755 9599 10771
rect 9508 10738 9518 10755
rect 9464 10721 9518 10738
rect 9552 10721 9599 10755
rect 9643 10768 9711 10771
rect 9643 10728 9656 10768
rect 9698 10728 9711 10768
rect 9643 10721 9659 10728
rect 9693 10721 9711 10728
rect 9745 10755 9803 10771
rect 9745 10721 9767 10755
rect 9801 10721 9803 10755
rect 4635 10623 4701 10645
rect 4635 10589 4649 10623
rect 4683 10589 4701 10623
rect 4971 10611 5021 10694
rect 9745 10705 9803 10721
rect 9837 10734 9887 10889
rect 9745 10687 9779 10705
rect 4635 10573 4701 10589
rect 4825 10595 4875 10611
rect 4825 10561 4841 10595
rect 4825 10519 4875 10561
rect 4909 10595 5021 10611
rect 4909 10561 4925 10595
rect 4959 10561 5021 10595
rect 4909 10553 5021 10561
rect 9369 10651 9427 10668
rect 9369 10617 9381 10651
rect 9415 10617 9427 10651
rect 9369 10523 9427 10617
rect 9501 10649 9779 10687
rect 9837 10698 9848 10734
rect 9882 10698 9887 10734
rect 9501 10627 9567 10649
rect 9501 10593 9515 10627
rect 9549 10593 9567 10627
rect 9837 10615 9887 10698
rect 9501 10577 9567 10593
rect 9691 10599 9741 10615
rect 9691 10565 9707 10599
rect 9691 10523 9741 10565
rect 9775 10599 9887 10615
rect 9775 10565 9791 10599
rect 9825 10565 9887 10599
rect 9775 10557 9887 10565
rect 4486 10485 4515 10519
rect 4549 10485 4607 10519
rect 4641 10485 4699 10519
rect 4733 10485 4791 10519
rect 4825 10485 4883 10519
rect 4917 10485 4975 10519
rect 5009 10485 5038 10519
rect 9352 10489 9381 10523
rect 9415 10489 9473 10523
rect 9507 10489 9565 10523
rect 9599 10489 9657 10523
rect 9691 10489 9749 10523
rect 9783 10489 9841 10523
rect 9875 10489 9904 10523
rect 6112 6583 6141 6617
rect 6175 6583 6233 6617
rect 6267 6583 6325 6617
rect 6359 6583 6407 6617
rect 6441 6583 6470 6617
rect 6178 6537 6244 6549
rect 6178 6503 6194 6537
rect 6228 6503 6244 6537
rect 6178 6469 6244 6503
rect 6178 6435 6194 6469
rect 6228 6435 6244 6469
rect 6178 6423 6244 6435
rect 6278 6537 6324 6583
rect 6312 6503 6324 6537
rect 6278 6469 6324 6503
rect 6312 6435 6324 6469
rect 6395 6489 6453 6583
rect 6395 6455 6407 6489
rect 6441 6455 6453 6489
rect 6395 6438 6453 6455
rect 6178 6382 6224 6423
rect 6278 6419 6324 6435
rect 6212 6348 6224 6382
rect 6178 6303 6224 6348
rect 6258 6350 6274 6385
rect 6308 6350 6324 6385
rect 6258 6337 6324 6350
rect 6178 6285 6244 6303
rect 6178 6251 6194 6285
rect 6228 6251 6244 6285
rect 6178 6217 6244 6251
rect 6178 6183 6194 6217
rect 6228 6183 6244 6217
rect 6178 6149 6244 6183
rect 6178 6115 6194 6149
rect 6228 6115 6244 6149
rect 6178 6107 6244 6115
rect 6278 6285 6320 6301
rect 6312 6251 6320 6285
rect 6278 6217 6320 6251
rect 6312 6183 6320 6217
rect 6278 6149 6320 6183
rect 6312 6115 6320 6149
rect 6278 6073 6320 6115
rect 6395 6271 6453 6306
rect 6395 6237 6407 6271
rect 6441 6237 6453 6271
rect 6395 6178 6453 6237
rect 6395 6144 6407 6178
rect 6441 6144 6453 6178
rect 6395 6073 6453 6144
rect 6112 6039 6141 6073
rect 6175 6039 6233 6073
rect 6267 6039 6325 6073
rect 6359 6039 6407 6073
rect 6441 6039 6470 6073
rect 9928 5951 9957 5985
rect 9991 5951 10047 5985
rect 10081 5951 10139 5985
rect 10173 5951 10231 5985
rect 10265 5951 10323 5985
rect 10357 5951 10415 5985
rect 10449 5951 10507 5985
rect 10541 5951 10599 5985
rect 10633 5951 10691 5985
rect 10725 5951 10783 5985
rect 10817 5951 10875 5985
rect 10909 5951 10967 5985
rect 11001 5951 11059 5985
rect 11093 5951 11151 5985
rect 11185 5951 11243 5985
rect 11277 5951 11335 5985
rect 11369 5951 11427 5985
rect 11461 5951 11490 5985
rect 9945 5857 10003 5951
rect 9945 5823 9957 5857
rect 9991 5823 10003 5857
rect 9945 5806 10003 5823
rect 10042 5873 10122 5917
rect 10171 5913 10237 5951
rect 10171 5879 10187 5913
rect 10221 5879 10237 5913
rect 10271 5901 10473 5917
rect 10042 5839 10088 5873
rect 10271 5867 10439 5901
rect 10271 5845 10305 5867
rect 10439 5849 10473 5867
rect 10540 5896 10574 5917
rect 10608 5913 10674 5951
rect 10608 5879 10624 5913
rect 10658 5879 10674 5913
rect 10708 5896 10742 5917
rect 10042 5806 10122 5839
rect 10157 5811 10305 5845
rect 10540 5845 10574 5862
rect 10776 5904 10842 5951
rect 10776 5870 10792 5904
rect 10826 5870 10842 5904
rect 10896 5896 10930 5917
rect 10708 5845 10742 5862
rect 9945 5639 10003 5674
rect 9945 5605 9957 5639
rect 9991 5605 10003 5639
rect 1746 5531 1775 5565
rect 1809 5531 1865 5565
rect 1899 5531 1957 5565
rect 1991 5531 2049 5565
rect 2083 5531 2141 5565
rect 2175 5531 2233 5565
rect 2267 5531 2325 5565
rect 2359 5531 2417 5565
rect 2451 5531 2509 5565
rect 2543 5531 2601 5565
rect 2635 5531 2693 5565
rect 2727 5531 2785 5565
rect 2819 5531 2877 5565
rect 2911 5531 2969 5565
rect 3003 5531 3061 5565
rect 3095 5531 3153 5565
rect 3187 5531 3245 5565
rect 3279 5531 3308 5565
rect 1763 5437 1821 5531
rect 1763 5403 1775 5437
rect 1809 5403 1821 5437
rect 1763 5386 1821 5403
rect 1860 5453 1940 5497
rect 1989 5493 2055 5531
rect 1989 5459 2005 5493
rect 2039 5459 2055 5493
rect 2089 5481 2291 5497
rect 1860 5419 1906 5453
rect 2089 5447 2257 5481
rect 2089 5425 2123 5447
rect 2257 5429 2291 5447
rect 2358 5476 2392 5497
rect 2426 5493 2492 5531
rect 2426 5459 2442 5493
rect 2476 5459 2492 5493
rect 2526 5476 2560 5497
rect 1860 5386 1940 5419
rect 1975 5391 2123 5425
rect 2358 5425 2392 5442
rect 2594 5484 2660 5531
rect 2594 5450 2610 5484
rect 2644 5450 2660 5484
rect 2714 5476 2748 5497
rect 2526 5425 2560 5442
rect 1763 5219 1821 5254
rect 1763 5185 1775 5219
rect 1809 5185 1821 5219
rect 1763 5126 1821 5185
rect 1763 5092 1775 5126
rect 1809 5092 1821 5126
rect 1763 5021 1821 5092
rect 1860 5251 1926 5386
rect 1975 5349 2009 5391
rect 1960 5333 2009 5349
rect 2216 5361 2228 5395
rect 2262 5361 2315 5395
rect 2358 5391 2560 5425
rect 2782 5493 2848 5531
rect 2782 5459 2798 5493
rect 2832 5459 2848 5493
rect 2882 5476 2916 5497
rect 2714 5425 2748 5442
rect 2882 5425 2916 5442
rect 2714 5391 2916 5425
rect 2966 5476 3086 5497
rect 3000 5442 3086 5476
rect 3139 5489 3205 5531
rect 3880 5523 3909 5557
rect 3943 5523 3999 5557
rect 4033 5523 4091 5557
rect 4125 5523 4183 5557
rect 4217 5523 4275 5557
rect 4309 5523 4367 5557
rect 4401 5523 4459 5557
rect 4493 5523 4551 5557
rect 4585 5523 4643 5557
rect 4677 5523 4735 5557
rect 4769 5523 4827 5557
rect 4861 5523 4919 5557
rect 4953 5523 5011 5557
rect 5045 5523 5103 5557
rect 5137 5523 5195 5557
rect 5229 5523 5287 5557
rect 5321 5523 5379 5557
rect 5413 5523 5442 5557
rect 5830 5523 5859 5557
rect 5893 5523 5951 5557
rect 5985 5523 6043 5557
rect 6077 5523 6135 5557
rect 6169 5523 6227 5557
rect 6261 5523 6319 5557
rect 6353 5523 6411 5557
rect 6445 5523 6503 5557
rect 6537 5523 6595 5557
rect 6629 5523 6687 5557
rect 6721 5523 6779 5557
rect 6813 5523 6871 5557
rect 6905 5523 6963 5557
rect 6997 5523 7055 5557
rect 7089 5523 7147 5557
rect 7181 5523 7239 5557
rect 7273 5523 7331 5557
rect 7365 5523 7394 5557
rect 7832 5529 7861 5563
rect 7895 5529 7953 5563
rect 7987 5529 8045 5563
rect 8079 5529 8137 5563
rect 8171 5529 8229 5563
rect 8263 5529 8321 5563
rect 8355 5529 8413 5563
rect 8447 5529 8505 5563
rect 8539 5529 8597 5563
rect 8631 5529 8689 5563
rect 8723 5529 8781 5563
rect 8815 5529 8873 5563
rect 8907 5529 8965 5563
rect 8999 5529 9057 5563
rect 9091 5529 9149 5563
rect 9183 5529 9241 5563
rect 9275 5529 9333 5563
rect 9367 5529 9396 5563
rect 9945 5546 10003 5605
rect 3139 5455 3155 5489
rect 3189 5455 3205 5489
rect 2966 5421 3086 5442
rect 3239 5453 3291 5497
rect 2966 5395 3205 5421
rect 2966 5361 2968 5395
rect 3002 5387 3205 5395
rect 3002 5361 3014 5387
rect 2216 5357 2315 5361
rect 1994 5299 2009 5333
rect 1960 5283 2009 5299
rect 2043 5327 2059 5341
rect 2043 5293 2044 5327
rect 2093 5307 2131 5341
rect 2216 5323 2299 5357
rect 2333 5323 2349 5357
rect 2383 5323 2399 5357
rect 2433 5327 2458 5357
rect 2078 5293 2131 5307
rect 2383 5293 2412 5323
rect 2446 5293 2458 5327
rect 2517 5298 2750 5355
rect 3171 5349 3205 5387
rect 3273 5419 3291 5453
rect 3239 5382 3291 5419
rect 1860 5213 1940 5251
rect 1860 5179 1906 5213
rect 1860 5123 1940 5179
rect 1975 5161 2009 5283
rect 2097 5229 2136 5259
rect 2097 5195 2131 5229
rect 2170 5225 2181 5259
rect 2517 5245 2551 5298
rect 2165 5195 2181 5225
rect 2227 5229 2484 5245
rect 2261 5211 2484 5229
rect 2518 5211 2551 5245
rect 2596 5259 2668 5261
rect 2630 5245 2668 5259
rect 2596 5211 2601 5225
rect 2635 5211 2668 5245
rect 2261 5195 2277 5211
rect 2596 5195 2668 5211
rect 2716 5229 2750 5298
rect 2784 5327 2862 5342
rect 3060 5333 3126 5349
rect 3060 5327 3092 5333
rect 2818 5326 2862 5327
rect 2818 5293 2828 5326
rect 2784 5292 2828 5293
rect 2784 5276 2862 5292
rect 2900 5293 2924 5327
rect 2958 5293 2974 5327
rect 3094 5293 3126 5299
rect 2900 5229 2934 5293
rect 3092 5283 3126 5293
rect 3171 5333 3222 5349
rect 3171 5299 3188 5333
rect 3171 5283 3222 5299
rect 2716 5195 2934 5229
rect 3002 5225 3048 5259
rect 2968 5222 3048 5225
rect 3171 5223 3205 5283
rect 3256 5251 3291 5382
rect 3897 5429 3955 5523
rect 3897 5395 3909 5429
rect 3943 5395 3955 5429
rect 3897 5378 3955 5395
rect 3994 5445 4074 5489
rect 4123 5485 4189 5523
rect 4123 5451 4139 5485
rect 4173 5451 4189 5485
rect 4223 5473 4425 5489
rect 3994 5411 4040 5445
rect 4223 5439 4391 5473
rect 4223 5417 4257 5439
rect 4391 5421 4425 5439
rect 4492 5468 4526 5489
rect 4560 5485 4626 5523
rect 4560 5451 4576 5485
rect 4610 5451 4626 5485
rect 4660 5468 4694 5489
rect 3994 5378 4074 5411
rect 4109 5383 4257 5417
rect 4492 5417 4526 5434
rect 4728 5476 4794 5523
rect 4728 5442 4744 5476
rect 4778 5442 4794 5476
rect 4848 5468 4882 5489
rect 4660 5417 4694 5434
rect 2227 5194 2277 5195
rect 1975 5127 2108 5161
rect 2227 5160 2236 5194
rect 2270 5160 2277 5194
rect 2968 5188 3014 5222
rect 2968 5172 3048 5188
rect 2227 5157 2277 5160
rect 1860 5089 1906 5123
rect 2074 5123 2108 5127
rect 2358 5127 2560 5161
rect 2074 5105 2291 5123
rect 1860 5055 1940 5089
rect 1974 5059 1990 5093
rect 2024 5059 2040 5093
rect 1974 5021 2040 5059
rect 2074 5071 2257 5105
rect 2074 5055 2291 5071
rect 2358 5110 2392 5127
rect 2526 5110 2560 5127
rect 2358 5055 2392 5076
rect 2426 5059 2442 5093
rect 2476 5059 2492 5093
rect 2426 5021 2492 5059
rect 2701 5127 2916 5161
rect 3087 5159 3205 5223
rect 3239 5210 3291 5251
rect 3273 5186 3291 5210
rect 3087 5135 3121 5159
rect 2701 5110 2748 5127
rect 2526 5055 2560 5076
rect 2594 5063 2610 5097
rect 2644 5063 2660 5097
rect 2594 5021 2660 5063
rect 2701 5076 2714 5110
rect 2882 5110 2916 5127
rect 2701 5055 2748 5076
rect 2782 5059 2798 5093
rect 2832 5059 2848 5093
rect 2782 5021 2848 5059
rect 2882 5055 2916 5076
rect 2966 5110 3121 5135
rect 3239 5150 3244 5176
rect 3284 5150 3291 5186
rect 3000 5076 3121 5110
rect 2966 5055 3121 5076
rect 3155 5101 3205 5118
rect 3189 5067 3205 5101
rect 3155 5021 3205 5067
rect 3239 5116 3291 5150
rect 3273 5082 3291 5116
rect 3239 5055 3291 5082
rect 3897 5211 3955 5246
rect 3897 5177 3909 5211
rect 3943 5177 3955 5211
rect 3897 5118 3955 5177
rect 3897 5084 3909 5118
rect 3943 5084 3955 5118
rect 1746 4987 1775 5021
rect 1809 4987 1865 5021
rect 1899 4987 1957 5021
rect 1991 4987 2049 5021
rect 2083 4987 2141 5021
rect 2175 4987 2233 5021
rect 2267 4987 2325 5021
rect 2359 4987 2417 5021
rect 2451 4987 2509 5021
rect 2543 4987 2601 5021
rect 2635 4987 2693 5021
rect 2727 4987 2785 5021
rect 2819 4987 2877 5021
rect 2911 4987 2969 5021
rect 3003 4987 3061 5021
rect 3095 4987 3153 5021
rect 3187 4987 3245 5021
rect 3279 4987 3308 5021
rect 3897 5013 3955 5084
rect 3994 5243 4060 5378
rect 4109 5341 4143 5383
rect 4094 5325 4143 5341
rect 4350 5353 4362 5387
rect 4396 5353 4449 5387
rect 4492 5383 4694 5417
rect 4916 5485 4982 5523
rect 4916 5451 4932 5485
rect 4966 5451 4982 5485
rect 5016 5468 5050 5489
rect 4848 5417 4882 5434
rect 5016 5417 5050 5434
rect 4848 5383 5050 5417
rect 5100 5468 5220 5489
rect 5134 5434 5220 5468
rect 5273 5481 5339 5523
rect 5273 5447 5289 5481
rect 5323 5447 5339 5481
rect 5100 5413 5220 5434
rect 5373 5445 5425 5489
rect 5100 5387 5339 5413
rect 5100 5353 5102 5387
rect 5136 5379 5339 5387
rect 5136 5353 5148 5379
rect 4350 5349 4449 5353
rect 4128 5291 4143 5325
rect 4094 5275 4143 5291
rect 4177 5319 4193 5333
rect 4177 5285 4178 5319
rect 4227 5299 4265 5333
rect 4350 5315 4433 5349
rect 4467 5315 4483 5349
rect 4517 5315 4533 5349
rect 4567 5319 4592 5349
rect 4212 5285 4265 5299
rect 4517 5285 4546 5315
rect 4580 5285 4592 5319
rect 4651 5290 4884 5347
rect 5305 5341 5339 5379
rect 5407 5411 5425 5445
rect 5373 5374 5425 5411
rect 5847 5429 5905 5523
rect 5847 5395 5859 5429
rect 5893 5395 5905 5429
rect 5847 5378 5905 5395
rect 5946 5445 6026 5489
rect 6075 5485 6141 5523
rect 6075 5451 6091 5485
rect 6125 5451 6141 5485
rect 6175 5473 6377 5489
rect 5946 5411 5992 5445
rect 6175 5439 6343 5473
rect 6175 5417 6209 5439
rect 6343 5421 6377 5439
rect 6444 5468 6478 5489
rect 6512 5485 6578 5523
rect 6512 5451 6528 5485
rect 6562 5451 6578 5485
rect 6612 5468 6646 5489
rect 5946 5378 6026 5411
rect 6061 5383 6209 5417
rect 6444 5417 6478 5434
rect 6680 5476 6746 5523
rect 6680 5442 6696 5476
rect 6730 5442 6746 5476
rect 6800 5468 6834 5489
rect 6612 5417 6646 5434
rect 3994 5205 4074 5243
rect 3994 5171 4040 5205
rect 3994 5115 4074 5171
rect 4109 5153 4143 5275
rect 4231 5221 4270 5251
rect 4231 5187 4265 5221
rect 4304 5217 4315 5251
rect 4651 5237 4685 5290
rect 4299 5187 4315 5217
rect 4361 5221 4618 5237
rect 4395 5203 4618 5221
rect 4652 5203 4685 5237
rect 4730 5251 4802 5253
rect 4764 5237 4802 5251
rect 4730 5203 4735 5217
rect 4769 5203 4802 5237
rect 4395 5187 4411 5203
rect 4730 5187 4802 5203
rect 4850 5221 4884 5290
rect 4918 5319 4996 5334
rect 5194 5325 5260 5341
rect 5194 5319 5226 5325
rect 4952 5318 4996 5319
rect 4952 5285 4962 5318
rect 4918 5284 4962 5285
rect 4918 5268 4996 5284
rect 5034 5285 5058 5319
rect 5092 5285 5108 5319
rect 5228 5285 5260 5291
rect 5034 5221 5068 5285
rect 5226 5275 5260 5285
rect 5305 5325 5356 5341
rect 5305 5291 5322 5325
rect 5305 5275 5356 5291
rect 4850 5187 5068 5221
rect 5136 5217 5182 5251
rect 5102 5214 5182 5217
rect 5305 5215 5339 5275
rect 5390 5243 5425 5374
rect 4361 5184 4411 5187
rect 4109 5119 4242 5153
rect 4361 5150 4368 5184
rect 4402 5150 4411 5184
rect 5102 5180 5148 5214
rect 5102 5164 5182 5180
rect 4361 5149 4411 5150
rect 3994 5081 4040 5115
rect 4208 5115 4242 5119
rect 4492 5119 4694 5153
rect 4208 5097 4425 5115
rect 3994 5047 4074 5081
rect 4108 5051 4124 5085
rect 4158 5051 4174 5085
rect 4108 5013 4174 5051
rect 4208 5063 4391 5097
rect 4208 5047 4425 5063
rect 4492 5102 4526 5119
rect 4660 5102 4694 5119
rect 4492 5047 4526 5068
rect 4560 5051 4576 5085
rect 4610 5051 4626 5085
rect 4560 5013 4626 5051
rect 4835 5119 5050 5153
rect 5221 5151 5339 5215
rect 5373 5202 5425 5243
rect 5407 5178 5425 5202
rect 5221 5127 5255 5151
rect 4835 5102 4882 5119
rect 4660 5047 4694 5068
rect 4728 5055 4744 5089
rect 4778 5055 4794 5089
rect 4728 5013 4794 5055
rect 4835 5068 4848 5102
rect 5016 5102 5050 5119
rect 4835 5047 4882 5068
rect 4916 5051 4932 5085
rect 4966 5051 4982 5085
rect 4916 5013 4982 5051
rect 5016 5047 5050 5068
rect 5100 5102 5255 5127
rect 5373 5142 5384 5168
rect 5418 5142 5425 5178
rect 5134 5068 5255 5102
rect 5100 5047 5255 5068
rect 5289 5093 5339 5110
rect 5323 5059 5339 5093
rect 5289 5013 5339 5059
rect 5373 5108 5425 5142
rect 5407 5074 5425 5108
rect 5373 5047 5425 5074
rect 5847 5211 5905 5246
rect 5847 5177 5859 5211
rect 5893 5177 5905 5211
rect 5847 5118 5905 5177
rect 5847 5084 5859 5118
rect 5893 5084 5905 5118
rect 5847 5013 5905 5084
rect 5946 5243 6012 5378
rect 6061 5341 6095 5383
rect 6046 5325 6095 5341
rect 6302 5353 6314 5387
rect 6348 5353 6401 5387
rect 6444 5383 6646 5417
rect 6868 5485 6934 5523
rect 6868 5451 6884 5485
rect 6918 5451 6934 5485
rect 6968 5468 7002 5489
rect 6800 5417 6834 5434
rect 6968 5417 7002 5434
rect 6800 5383 7002 5417
rect 7052 5468 7172 5489
rect 7086 5434 7172 5468
rect 7225 5481 7291 5523
rect 7225 5447 7241 5481
rect 7275 5447 7291 5481
rect 7052 5413 7172 5434
rect 7325 5445 7377 5489
rect 7052 5387 7291 5413
rect 7052 5353 7054 5387
rect 7088 5379 7291 5387
rect 7088 5353 7100 5379
rect 6302 5349 6401 5353
rect 6080 5291 6095 5325
rect 6046 5275 6095 5291
rect 6129 5319 6145 5333
rect 6129 5285 6130 5319
rect 6179 5299 6217 5333
rect 6302 5315 6385 5349
rect 6419 5315 6435 5349
rect 6469 5315 6485 5349
rect 6519 5319 6544 5349
rect 6164 5285 6217 5299
rect 6469 5285 6498 5315
rect 6532 5285 6544 5319
rect 6603 5290 6836 5347
rect 7257 5341 7291 5379
rect 7359 5411 7377 5445
rect 7325 5374 7377 5411
rect 7849 5435 7907 5529
rect 7849 5401 7861 5435
rect 7895 5401 7907 5435
rect 7849 5384 7907 5401
rect 7948 5451 8028 5495
rect 8077 5491 8143 5529
rect 8077 5457 8093 5491
rect 8127 5457 8143 5491
rect 8177 5479 8379 5495
rect 7948 5417 7994 5451
rect 8177 5445 8345 5479
rect 8177 5423 8211 5445
rect 8345 5427 8379 5445
rect 8446 5474 8480 5495
rect 8514 5491 8580 5529
rect 8514 5457 8530 5491
rect 8564 5457 8580 5491
rect 8614 5474 8648 5495
rect 7948 5384 8028 5417
rect 8063 5389 8211 5423
rect 8446 5423 8480 5440
rect 8682 5482 8748 5529
rect 8682 5448 8698 5482
rect 8732 5448 8748 5482
rect 8802 5474 8836 5495
rect 8614 5423 8648 5440
rect 5946 5205 6026 5243
rect 5946 5171 5992 5205
rect 5946 5115 6026 5171
rect 6061 5153 6095 5275
rect 6183 5221 6222 5251
rect 6183 5187 6217 5221
rect 6256 5217 6267 5251
rect 6603 5237 6637 5290
rect 6251 5187 6267 5217
rect 6313 5221 6570 5237
rect 6347 5203 6570 5221
rect 6604 5203 6637 5237
rect 6682 5251 6754 5253
rect 6716 5237 6754 5251
rect 6682 5203 6687 5217
rect 6721 5203 6754 5237
rect 6347 5187 6363 5203
rect 6682 5187 6754 5203
rect 6802 5221 6836 5290
rect 6870 5319 6948 5334
rect 7146 5325 7212 5341
rect 7146 5319 7178 5325
rect 6904 5318 6948 5319
rect 6904 5285 6914 5318
rect 6870 5284 6914 5285
rect 6870 5268 6948 5284
rect 6986 5285 7010 5319
rect 7044 5285 7060 5319
rect 7180 5285 7212 5291
rect 6986 5221 7020 5285
rect 7178 5275 7212 5285
rect 7257 5325 7308 5341
rect 7257 5291 7274 5325
rect 7257 5275 7308 5291
rect 6802 5187 7020 5221
rect 7088 5217 7134 5251
rect 7054 5214 7134 5217
rect 7257 5215 7291 5275
rect 7342 5243 7377 5374
rect 6313 5184 6363 5187
rect 6061 5119 6194 5153
rect 6313 5150 6320 5184
rect 6354 5150 6363 5184
rect 7054 5180 7100 5214
rect 7054 5164 7134 5180
rect 6313 5149 6363 5150
rect 5946 5081 5992 5115
rect 6160 5115 6194 5119
rect 6444 5119 6646 5153
rect 6160 5097 6377 5115
rect 5946 5047 6026 5081
rect 6060 5051 6076 5085
rect 6110 5051 6126 5085
rect 6060 5013 6126 5051
rect 6160 5063 6343 5097
rect 6160 5047 6377 5063
rect 6444 5102 6478 5119
rect 6612 5102 6646 5119
rect 6444 5047 6478 5068
rect 6512 5051 6528 5085
rect 6562 5051 6578 5085
rect 6512 5013 6578 5051
rect 6787 5119 7002 5153
rect 7173 5151 7291 5215
rect 7325 5202 7377 5243
rect 7359 5178 7377 5202
rect 7173 5127 7207 5151
rect 6787 5102 6834 5119
rect 6612 5047 6646 5068
rect 6680 5055 6696 5089
rect 6730 5055 6746 5089
rect 6680 5013 6746 5055
rect 6787 5068 6800 5102
rect 6968 5102 7002 5119
rect 6787 5047 6834 5068
rect 6868 5051 6884 5085
rect 6918 5051 6934 5085
rect 6868 5013 6934 5051
rect 6968 5047 7002 5068
rect 7052 5102 7207 5127
rect 7325 5142 7336 5168
rect 7370 5142 7377 5178
rect 7086 5068 7207 5102
rect 7052 5047 7207 5068
rect 7241 5093 7291 5110
rect 7275 5059 7291 5093
rect 7241 5013 7291 5059
rect 7325 5108 7377 5142
rect 7359 5074 7377 5108
rect 7325 5047 7377 5074
rect 7849 5217 7907 5252
rect 7849 5183 7861 5217
rect 7895 5183 7907 5217
rect 7849 5124 7907 5183
rect 7849 5090 7861 5124
rect 7895 5090 7907 5124
rect 7849 5019 7907 5090
rect 7948 5249 8014 5384
rect 8063 5347 8097 5389
rect 8048 5331 8097 5347
rect 8304 5359 8316 5393
rect 8350 5359 8403 5393
rect 8446 5389 8648 5423
rect 8870 5491 8936 5529
rect 8870 5457 8886 5491
rect 8920 5457 8936 5491
rect 8970 5474 9004 5495
rect 8802 5423 8836 5440
rect 8970 5423 9004 5440
rect 8802 5389 9004 5423
rect 9054 5474 9174 5495
rect 9088 5440 9174 5474
rect 9227 5487 9293 5529
rect 9945 5512 9957 5546
rect 9991 5512 10003 5546
rect 9227 5453 9243 5487
rect 9277 5453 9293 5487
rect 9054 5419 9174 5440
rect 9327 5451 9379 5495
rect 9054 5393 9293 5419
rect 9054 5359 9056 5393
rect 9090 5385 9293 5393
rect 9090 5359 9102 5385
rect 8304 5355 8403 5359
rect 8082 5297 8097 5331
rect 8048 5281 8097 5297
rect 8131 5325 8147 5339
rect 8131 5291 8132 5325
rect 8181 5305 8219 5339
rect 8304 5321 8387 5355
rect 8421 5321 8437 5355
rect 8471 5321 8487 5355
rect 8521 5325 8546 5355
rect 8166 5291 8219 5305
rect 8471 5291 8500 5321
rect 8534 5291 8546 5325
rect 8605 5296 8838 5353
rect 9259 5347 9293 5385
rect 9361 5417 9379 5451
rect 9945 5441 10003 5512
rect 10042 5671 10108 5806
rect 10157 5769 10191 5811
rect 10142 5753 10191 5769
rect 10398 5781 10410 5815
rect 10444 5781 10497 5815
rect 10540 5811 10742 5845
rect 10964 5913 11030 5951
rect 10964 5879 10980 5913
rect 11014 5879 11030 5913
rect 11064 5896 11098 5917
rect 10896 5845 10930 5862
rect 11064 5845 11098 5862
rect 10896 5811 11098 5845
rect 11148 5896 11268 5917
rect 11182 5862 11268 5896
rect 11321 5909 11387 5951
rect 11988 5939 12017 5973
rect 12051 5939 12109 5973
rect 12143 5939 12201 5973
rect 12235 5939 12293 5973
rect 12327 5939 12385 5973
rect 12419 5939 12477 5973
rect 12511 5939 12569 5973
rect 12603 5939 12661 5973
rect 12695 5939 12753 5973
rect 12787 5939 12845 5973
rect 12879 5939 12937 5973
rect 12971 5939 13029 5973
rect 13063 5939 13121 5973
rect 13155 5939 13213 5973
rect 13247 5939 13305 5973
rect 13339 5939 13397 5973
rect 13431 5939 13489 5973
rect 13523 5939 13552 5973
rect 13946 5947 13975 5981
rect 14009 5947 14067 5981
rect 14101 5947 14159 5981
rect 14193 5947 14251 5981
rect 14285 5947 14343 5981
rect 14377 5947 14435 5981
rect 14469 5947 14527 5981
rect 14561 5947 14619 5981
rect 14653 5947 14711 5981
rect 14745 5947 14803 5981
rect 14837 5947 14895 5981
rect 14929 5947 14987 5981
rect 15021 5947 15079 5981
rect 15113 5947 15171 5981
rect 15205 5947 15263 5981
rect 15297 5947 15355 5981
rect 15389 5947 15447 5981
rect 15481 5947 15510 5981
rect 15942 5953 15971 5987
rect 16005 5953 16061 5987
rect 16095 5953 16153 5987
rect 16187 5953 16245 5987
rect 16279 5953 16337 5987
rect 16371 5953 16429 5987
rect 16463 5953 16521 5987
rect 16555 5953 16613 5987
rect 16647 5953 16705 5987
rect 16739 5953 16797 5987
rect 16831 5953 16889 5987
rect 16923 5953 16981 5987
rect 17015 5953 17073 5987
rect 17107 5953 17165 5987
rect 17199 5953 17257 5987
rect 17291 5953 17349 5987
rect 17383 5953 17441 5987
rect 17475 5953 17504 5987
rect 11321 5875 11337 5909
rect 11371 5875 11387 5909
rect 11148 5841 11268 5862
rect 11421 5873 11473 5917
rect 11148 5815 11387 5841
rect 11148 5781 11150 5815
rect 11184 5807 11387 5815
rect 11184 5781 11196 5807
rect 10398 5777 10497 5781
rect 10176 5719 10191 5753
rect 10142 5703 10191 5719
rect 10225 5747 10241 5761
rect 10225 5713 10226 5747
rect 10275 5727 10313 5761
rect 10398 5743 10481 5777
rect 10515 5743 10531 5777
rect 10565 5743 10581 5777
rect 10615 5747 10640 5777
rect 10260 5713 10313 5727
rect 10565 5713 10594 5743
rect 10628 5713 10640 5747
rect 10699 5718 10932 5775
rect 11353 5769 11387 5807
rect 11455 5839 11473 5873
rect 11421 5802 11473 5839
rect 10042 5633 10122 5671
rect 10042 5599 10088 5633
rect 10042 5543 10122 5599
rect 10157 5581 10191 5703
rect 10279 5649 10318 5679
rect 10279 5615 10313 5649
rect 10352 5645 10363 5679
rect 10699 5665 10733 5718
rect 10347 5615 10363 5645
rect 10409 5649 10666 5665
rect 10443 5631 10666 5649
rect 10700 5631 10733 5665
rect 10778 5679 10850 5681
rect 10812 5665 10850 5679
rect 10778 5631 10783 5645
rect 10817 5631 10850 5665
rect 10443 5615 10459 5631
rect 10778 5615 10850 5631
rect 10898 5649 10932 5718
rect 10966 5747 11044 5762
rect 11242 5753 11308 5769
rect 11242 5747 11274 5753
rect 11000 5746 11044 5747
rect 11000 5713 11010 5746
rect 10966 5712 11010 5713
rect 10966 5696 11044 5712
rect 11082 5713 11106 5747
rect 11140 5713 11156 5747
rect 11276 5713 11308 5719
rect 11082 5649 11116 5713
rect 11274 5703 11308 5713
rect 11353 5753 11404 5769
rect 11353 5719 11370 5753
rect 11353 5703 11404 5719
rect 10898 5615 11116 5649
rect 11184 5645 11230 5679
rect 11150 5642 11230 5645
rect 11353 5643 11387 5703
rect 11438 5671 11473 5802
rect 12005 5845 12063 5939
rect 12005 5811 12017 5845
rect 12051 5811 12063 5845
rect 12005 5794 12063 5811
rect 12104 5861 12184 5905
rect 12233 5901 12299 5939
rect 12233 5867 12249 5901
rect 12283 5867 12299 5901
rect 12333 5889 12535 5905
rect 12104 5827 12150 5861
rect 12333 5855 12501 5889
rect 12333 5833 12367 5855
rect 12501 5837 12535 5855
rect 12602 5884 12636 5905
rect 12670 5901 12736 5939
rect 12670 5867 12686 5901
rect 12720 5867 12736 5901
rect 12770 5884 12804 5905
rect 12104 5794 12184 5827
rect 12219 5799 12367 5833
rect 12602 5833 12636 5850
rect 12838 5892 12904 5939
rect 12838 5858 12854 5892
rect 12888 5858 12904 5892
rect 12958 5884 12992 5905
rect 12770 5833 12804 5850
rect 10409 5614 10459 5615
rect 10157 5547 10290 5581
rect 10409 5580 10418 5614
rect 10452 5580 10459 5614
rect 11150 5608 11196 5642
rect 11150 5592 11230 5608
rect 10409 5577 10459 5580
rect 10042 5509 10088 5543
rect 10256 5543 10290 5547
rect 10540 5547 10742 5581
rect 10256 5525 10473 5543
rect 10042 5475 10122 5509
rect 10156 5479 10172 5513
rect 10206 5479 10222 5513
rect 10156 5441 10222 5479
rect 10256 5491 10439 5525
rect 10256 5475 10473 5491
rect 10540 5530 10574 5547
rect 10708 5530 10742 5547
rect 10540 5475 10574 5496
rect 10608 5479 10624 5513
rect 10658 5479 10674 5513
rect 10608 5441 10674 5479
rect 10883 5547 11098 5581
rect 11269 5579 11387 5643
rect 11421 5630 11473 5671
rect 11455 5606 11473 5630
rect 11269 5555 11303 5579
rect 10883 5530 10930 5547
rect 10708 5475 10742 5496
rect 10776 5483 10792 5517
rect 10826 5483 10842 5517
rect 10776 5441 10842 5483
rect 10883 5496 10896 5530
rect 11064 5530 11098 5547
rect 10883 5475 10930 5496
rect 10964 5479 10980 5513
rect 11014 5479 11030 5513
rect 10964 5441 11030 5479
rect 11064 5475 11098 5496
rect 11148 5530 11303 5555
rect 11421 5570 11426 5596
rect 11466 5570 11473 5606
rect 11182 5496 11303 5530
rect 11148 5475 11303 5496
rect 11337 5521 11387 5538
rect 11371 5487 11387 5521
rect 11337 5441 11387 5487
rect 11421 5536 11473 5570
rect 11455 5502 11473 5536
rect 11421 5475 11473 5502
rect 12005 5627 12063 5662
rect 12005 5593 12017 5627
rect 12051 5593 12063 5627
rect 12005 5534 12063 5593
rect 12005 5500 12017 5534
rect 12051 5500 12063 5534
rect 9327 5380 9379 5417
rect 9928 5407 9957 5441
rect 9991 5407 10047 5441
rect 10081 5407 10139 5441
rect 10173 5407 10231 5441
rect 10265 5407 10323 5441
rect 10357 5407 10415 5441
rect 10449 5407 10507 5441
rect 10541 5407 10599 5441
rect 10633 5407 10691 5441
rect 10725 5407 10783 5441
rect 10817 5407 10875 5441
rect 10909 5407 10967 5441
rect 11001 5407 11059 5441
rect 11093 5407 11151 5441
rect 11185 5407 11243 5441
rect 11277 5407 11335 5441
rect 11369 5407 11427 5441
rect 11461 5407 11490 5441
rect 12005 5429 12063 5500
rect 12104 5659 12170 5794
rect 12219 5757 12253 5799
rect 12204 5741 12253 5757
rect 12460 5769 12472 5803
rect 12506 5769 12559 5803
rect 12602 5799 12804 5833
rect 13026 5901 13092 5939
rect 13026 5867 13042 5901
rect 13076 5867 13092 5901
rect 13126 5884 13160 5905
rect 12958 5833 12992 5850
rect 13126 5833 13160 5850
rect 12958 5799 13160 5833
rect 13210 5884 13330 5905
rect 13244 5850 13330 5884
rect 13383 5897 13449 5939
rect 13383 5863 13399 5897
rect 13433 5863 13449 5897
rect 13210 5829 13330 5850
rect 13483 5861 13535 5905
rect 13210 5803 13449 5829
rect 13210 5769 13212 5803
rect 13246 5795 13449 5803
rect 13246 5769 13258 5795
rect 12460 5765 12559 5769
rect 12238 5707 12253 5741
rect 12204 5691 12253 5707
rect 12287 5735 12303 5749
rect 12287 5701 12288 5735
rect 12337 5715 12375 5749
rect 12460 5731 12543 5765
rect 12577 5731 12593 5765
rect 12627 5731 12643 5765
rect 12677 5735 12702 5765
rect 12322 5701 12375 5715
rect 12627 5701 12656 5731
rect 12690 5701 12702 5735
rect 12761 5706 12994 5763
rect 13415 5757 13449 5795
rect 13517 5827 13535 5861
rect 13483 5790 13535 5827
rect 13963 5853 14021 5947
rect 13963 5819 13975 5853
rect 14009 5819 14021 5853
rect 13963 5802 14021 5819
rect 14062 5869 14142 5913
rect 14191 5909 14257 5947
rect 14191 5875 14207 5909
rect 14241 5875 14257 5909
rect 14291 5897 14493 5913
rect 14062 5835 14108 5869
rect 14291 5863 14459 5897
rect 14291 5841 14325 5863
rect 14459 5845 14493 5863
rect 14560 5892 14594 5913
rect 14628 5909 14694 5947
rect 14628 5875 14644 5909
rect 14678 5875 14694 5909
rect 14728 5892 14762 5913
rect 14062 5802 14142 5835
rect 14177 5807 14325 5841
rect 14560 5841 14594 5858
rect 14796 5900 14862 5947
rect 14796 5866 14812 5900
rect 14846 5866 14862 5900
rect 14916 5892 14950 5913
rect 14728 5841 14762 5858
rect 12104 5621 12184 5659
rect 12104 5587 12150 5621
rect 12104 5531 12184 5587
rect 12219 5569 12253 5691
rect 12341 5637 12380 5667
rect 12341 5603 12375 5637
rect 12414 5633 12425 5667
rect 12761 5653 12795 5706
rect 12409 5603 12425 5633
rect 12471 5637 12728 5653
rect 12505 5619 12728 5637
rect 12762 5619 12795 5653
rect 12840 5667 12912 5669
rect 12874 5653 12912 5667
rect 12840 5619 12845 5633
rect 12879 5619 12912 5653
rect 12505 5603 12521 5619
rect 12840 5603 12912 5619
rect 12960 5637 12994 5706
rect 13028 5735 13106 5750
rect 13304 5741 13370 5757
rect 13304 5735 13336 5741
rect 13062 5734 13106 5735
rect 13062 5701 13072 5734
rect 13028 5700 13072 5701
rect 13028 5684 13106 5700
rect 13144 5701 13168 5735
rect 13202 5701 13218 5735
rect 13338 5701 13370 5707
rect 13144 5637 13178 5701
rect 13336 5691 13370 5701
rect 13415 5741 13466 5757
rect 13415 5707 13432 5741
rect 13415 5691 13466 5707
rect 12960 5603 13178 5637
rect 13246 5633 13292 5667
rect 13212 5630 13292 5633
rect 13415 5631 13449 5691
rect 13500 5659 13535 5790
rect 12471 5600 12521 5603
rect 12219 5535 12352 5569
rect 12471 5566 12478 5600
rect 12512 5566 12521 5600
rect 13212 5596 13258 5630
rect 13212 5580 13292 5596
rect 12471 5565 12521 5566
rect 12104 5497 12150 5531
rect 12318 5531 12352 5535
rect 12602 5535 12804 5569
rect 12318 5513 12535 5531
rect 12104 5463 12184 5497
rect 12218 5467 12234 5501
rect 12268 5467 12284 5501
rect 12218 5429 12284 5467
rect 12318 5479 12501 5513
rect 12318 5463 12535 5479
rect 12602 5518 12636 5535
rect 12770 5518 12804 5535
rect 12602 5463 12636 5484
rect 12670 5467 12686 5501
rect 12720 5467 12736 5501
rect 12670 5429 12736 5467
rect 12945 5535 13160 5569
rect 13331 5567 13449 5631
rect 13483 5618 13535 5659
rect 13517 5594 13535 5618
rect 13331 5543 13365 5567
rect 12945 5518 12992 5535
rect 12770 5463 12804 5484
rect 12838 5471 12854 5505
rect 12888 5471 12904 5505
rect 12838 5429 12904 5471
rect 12945 5484 12958 5518
rect 13126 5518 13160 5535
rect 12945 5463 12992 5484
rect 13026 5467 13042 5501
rect 13076 5467 13092 5501
rect 13026 5429 13092 5467
rect 13126 5463 13160 5484
rect 13210 5518 13365 5543
rect 13483 5558 13494 5584
rect 13528 5558 13535 5594
rect 13244 5484 13365 5518
rect 13210 5463 13365 5484
rect 13399 5509 13449 5526
rect 13433 5475 13449 5509
rect 13399 5429 13449 5475
rect 13483 5524 13535 5558
rect 13517 5490 13535 5524
rect 13483 5463 13535 5490
rect 13963 5635 14021 5670
rect 13963 5601 13975 5635
rect 14009 5601 14021 5635
rect 13963 5542 14021 5601
rect 13963 5508 13975 5542
rect 14009 5508 14021 5542
rect 13963 5437 14021 5508
rect 14062 5667 14128 5802
rect 14177 5765 14211 5807
rect 14162 5749 14211 5765
rect 14418 5777 14430 5811
rect 14464 5777 14517 5811
rect 14560 5807 14762 5841
rect 14984 5909 15050 5947
rect 14984 5875 15000 5909
rect 15034 5875 15050 5909
rect 15084 5892 15118 5913
rect 14916 5841 14950 5858
rect 15084 5841 15118 5858
rect 14916 5807 15118 5841
rect 15168 5892 15288 5913
rect 15202 5858 15288 5892
rect 15341 5905 15407 5947
rect 15341 5871 15357 5905
rect 15391 5871 15407 5905
rect 15168 5837 15288 5858
rect 15441 5869 15493 5913
rect 15168 5811 15407 5837
rect 15168 5777 15170 5811
rect 15204 5803 15407 5811
rect 15204 5777 15216 5803
rect 14418 5773 14517 5777
rect 14196 5715 14211 5749
rect 14162 5699 14211 5715
rect 14245 5743 14261 5757
rect 14245 5709 14246 5743
rect 14295 5723 14333 5757
rect 14418 5739 14501 5773
rect 14535 5739 14551 5773
rect 14585 5739 14601 5773
rect 14635 5743 14660 5773
rect 14280 5709 14333 5723
rect 14585 5709 14614 5739
rect 14648 5709 14660 5743
rect 14719 5714 14952 5771
rect 15373 5765 15407 5803
rect 15475 5835 15493 5869
rect 15441 5798 15493 5835
rect 15959 5859 16017 5953
rect 15959 5825 15971 5859
rect 16005 5825 16017 5859
rect 15959 5808 16017 5825
rect 16056 5875 16136 5919
rect 16185 5915 16251 5953
rect 16185 5881 16201 5915
rect 16235 5881 16251 5915
rect 16285 5903 16487 5919
rect 16056 5841 16102 5875
rect 16285 5869 16453 5903
rect 16285 5847 16319 5869
rect 16453 5851 16487 5869
rect 16554 5898 16588 5919
rect 16622 5915 16688 5953
rect 16622 5881 16638 5915
rect 16672 5881 16688 5915
rect 16722 5898 16756 5919
rect 16056 5808 16136 5841
rect 16171 5813 16319 5847
rect 16554 5847 16588 5864
rect 16790 5906 16856 5953
rect 16790 5872 16806 5906
rect 16840 5872 16856 5906
rect 16910 5898 16944 5919
rect 16722 5847 16756 5864
rect 14062 5629 14142 5667
rect 14062 5595 14108 5629
rect 14062 5539 14142 5595
rect 14177 5577 14211 5699
rect 14299 5645 14338 5675
rect 14299 5611 14333 5645
rect 14372 5641 14383 5675
rect 14719 5661 14753 5714
rect 14367 5611 14383 5641
rect 14429 5645 14686 5661
rect 14463 5627 14686 5645
rect 14720 5627 14753 5661
rect 14798 5675 14870 5677
rect 14832 5661 14870 5675
rect 14798 5627 14803 5641
rect 14837 5627 14870 5661
rect 14463 5611 14479 5627
rect 14798 5611 14870 5627
rect 14918 5645 14952 5714
rect 14986 5743 15064 5758
rect 15262 5749 15328 5765
rect 15262 5743 15294 5749
rect 15020 5742 15064 5743
rect 15020 5709 15030 5742
rect 14986 5708 15030 5709
rect 14986 5692 15064 5708
rect 15102 5709 15126 5743
rect 15160 5709 15176 5743
rect 15296 5709 15328 5715
rect 15102 5645 15136 5709
rect 15294 5699 15328 5709
rect 15373 5749 15424 5765
rect 15373 5715 15390 5749
rect 15373 5699 15424 5715
rect 14918 5611 15136 5645
rect 15204 5641 15250 5675
rect 15170 5638 15250 5641
rect 15373 5639 15407 5699
rect 15458 5667 15493 5798
rect 14429 5608 14479 5611
rect 14177 5543 14310 5577
rect 14429 5574 14436 5608
rect 14470 5574 14479 5608
rect 15170 5604 15216 5638
rect 15170 5588 15250 5604
rect 14429 5573 14479 5574
rect 14062 5505 14108 5539
rect 14276 5539 14310 5543
rect 14560 5543 14762 5577
rect 14276 5521 14493 5539
rect 14062 5471 14142 5505
rect 14176 5475 14192 5509
rect 14226 5475 14242 5509
rect 14176 5437 14242 5475
rect 14276 5487 14459 5521
rect 14276 5471 14493 5487
rect 14560 5526 14594 5543
rect 14728 5526 14762 5543
rect 14560 5471 14594 5492
rect 14628 5475 14644 5509
rect 14678 5475 14694 5509
rect 14628 5437 14694 5475
rect 14903 5543 15118 5577
rect 15289 5575 15407 5639
rect 15441 5626 15493 5667
rect 15475 5602 15493 5626
rect 15289 5551 15323 5575
rect 14903 5526 14950 5543
rect 14728 5471 14762 5492
rect 14796 5479 14812 5513
rect 14846 5479 14862 5513
rect 14796 5437 14862 5479
rect 14903 5492 14916 5526
rect 15084 5526 15118 5543
rect 14903 5471 14950 5492
rect 14984 5475 15000 5509
rect 15034 5475 15050 5509
rect 14984 5437 15050 5475
rect 15084 5471 15118 5492
rect 15168 5526 15323 5551
rect 15441 5566 15452 5592
rect 15486 5566 15493 5602
rect 15202 5492 15323 5526
rect 15168 5471 15323 5492
rect 15357 5517 15407 5534
rect 15391 5483 15407 5517
rect 15357 5437 15407 5483
rect 15441 5532 15493 5566
rect 15475 5498 15493 5532
rect 15441 5471 15493 5498
rect 15959 5641 16017 5676
rect 15959 5607 15971 5641
rect 16005 5607 16017 5641
rect 15959 5548 16017 5607
rect 15959 5514 15971 5548
rect 16005 5514 16017 5548
rect 15959 5443 16017 5514
rect 16056 5673 16122 5808
rect 16171 5771 16205 5813
rect 16156 5755 16205 5771
rect 16412 5783 16424 5817
rect 16458 5783 16511 5817
rect 16554 5813 16756 5847
rect 16978 5915 17044 5953
rect 16978 5881 16994 5915
rect 17028 5881 17044 5915
rect 17078 5898 17112 5919
rect 16910 5847 16944 5864
rect 17078 5847 17112 5864
rect 16910 5813 17112 5847
rect 17162 5898 17282 5919
rect 17196 5864 17282 5898
rect 17335 5911 17401 5953
rect 17335 5877 17351 5911
rect 17385 5877 17401 5911
rect 17162 5843 17282 5864
rect 17435 5875 17487 5919
rect 17162 5817 17401 5843
rect 17162 5783 17164 5817
rect 17198 5809 17401 5817
rect 17198 5783 17210 5809
rect 16412 5779 16511 5783
rect 16190 5721 16205 5755
rect 16156 5705 16205 5721
rect 16239 5749 16255 5763
rect 16239 5715 16240 5749
rect 16289 5729 16327 5763
rect 16412 5745 16495 5779
rect 16529 5745 16545 5779
rect 16579 5745 16595 5779
rect 16629 5749 16654 5779
rect 16274 5715 16327 5729
rect 16579 5715 16608 5745
rect 16642 5715 16654 5749
rect 16713 5720 16946 5777
rect 17367 5771 17401 5809
rect 17469 5841 17487 5875
rect 17435 5804 17487 5841
rect 16056 5635 16136 5673
rect 16056 5601 16102 5635
rect 16056 5545 16136 5601
rect 16171 5583 16205 5705
rect 16293 5651 16332 5681
rect 16293 5617 16327 5651
rect 16366 5647 16377 5681
rect 16713 5667 16747 5720
rect 16361 5617 16377 5647
rect 16423 5651 16680 5667
rect 16457 5633 16680 5651
rect 16714 5633 16747 5667
rect 16792 5681 16864 5683
rect 16826 5667 16864 5681
rect 16792 5633 16797 5647
rect 16831 5633 16864 5667
rect 16457 5617 16473 5633
rect 16792 5617 16864 5633
rect 16912 5651 16946 5720
rect 16980 5749 17058 5764
rect 17256 5755 17322 5771
rect 17256 5749 17288 5755
rect 17014 5748 17058 5749
rect 17014 5715 17024 5748
rect 16980 5714 17024 5715
rect 16980 5698 17058 5714
rect 17096 5715 17120 5749
rect 17154 5715 17170 5749
rect 17290 5715 17322 5721
rect 17096 5651 17130 5715
rect 17288 5705 17322 5715
rect 17367 5755 17418 5771
rect 17367 5721 17384 5755
rect 17367 5705 17418 5721
rect 16912 5617 17130 5651
rect 17198 5647 17244 5681
rect 17164 5644 17244 5647
rect 17367 5645 17401 5705
rect 17452 5673 17487 5804
rect 16423 5614 16473 5617
rect 16171 5549 16304 5583
rect 16423 5580 16430 5614
rect 16464 5580 16473 5614
rect 17164 5610 17210 5644
rect 17164 5594 17244 5610
rect 16423 5579 16473 5580
rect 16056 5511 16102 5545
rect 16270 5545 16304 5549
rect 16554 5549 16756 5583
rect 16270 5527 16487 5545
rect 16056 5477 16136 5511
rect 16170 5481 16186 5515
rect 16220 5481 16236 5515
rect 16170 5443 16236 5481
rect 16270 5493 16453 5527
rect 16270 5477 16487 5493
rect 16554 5532 16588 5549
rect 16722 5532 16756 5549
rect 16554 5477 16588 5498
rect 16622 5481 16638 5515
rect 16672 5481 16688 5515
rect 16622 5443 16688 5481
rect 16897 5549 17112 5583
rect 17283 5581 17401 5645
rect 17435 5632 17487 5673
rect 17469 5608 17487 5632
rect 17283 5557 17317 5581
rect 16897 5532 16944 5549
rect 16722 5477 16756 5498
rect 16790 5485 16806 5519
rect 16840 5485 16856 5519
rect 16790 5443 16856 5485
rect 16897 5498 16910 5532
rect 17078 5532 17112 5549
rect 16897 5477 16944 5498
rect 16978 5481 16994 5515
rect 17028 5481 17044 5515
rect 16978 5443 17044 5481
rect 17078 5477 17112 5498
rect 17162 5532 17317 5557
rect 17435 5572 17446 5598
rect 17480 5572 17487 5608
rect 17196 5498 17317 5532
rect 17162 5477 17317 5498
rect 17351 5523 17401 5540
rect 17385 5489 17401 5523
rect 17351 5443 17401 5489
rect 17435 5538 17487 5572
rect 17469 5504 17487 5538
rect 17435 5477 17487 5504
rect 11988 5395 12017 5429
rect 12051 5395 12109 5429
rect 12143 5395 12201 5429
rect 12235 5395 12293 5429
rect 12327 5395 12385 5429
rect 12419 5395 12477 5429
rect 12511 5395 12569 5429
rect 12603 5395 12661 5429
rect 12695 5395 12753 5429
rect 12787 5395 12845 5429
rect 12879 5395 12937 5429
rect 12971 5395 13029 5429
rect 13063 5395 13121 5429
rect 13155 5395 13213 5429
rect 13247 5395 13305 5429
rect 13339 5395 13397 5429
rect 13431 5395 13489 5429
rect 13523 5395 13552 5429
rect 13946 5403 13975 5437
rect 14009 5403 14067 5437
rect 14101 5403 14159 5437
rect 14193 5403 14251 5437
rect 14285 5403 14343 5437
rect 14377 5403 14435 5437
rect 14469 5403 14527 5437
rect 14561 5403 14619 5437
rect 14653 5403 14711 5437
rect 14745 5403 14803 5437
rect 14837 5403 14895 5437
rect 14929 5403 14987 5437
rect 15021 5403 15079 5437
rect 15113 5403 15171 5437
rect 15205 5403 15263 5437
rect 15297 5403 15355 5437
rect 15389 5403 15447 5437
rect 15481 5403 15510 5437
rect 15942 5409 15971 5443
rect 16005 5409 16061 5443
rect 16095 5409 16153 5443
rect 16187 5409 16245 5443
rect 16279 5409 16337 5443
rect 16371 5409 16429 5443
rect 16463 5409 16521 5443
rect 16555 5409 16613 5443
rect 16647 5409 16705 5443
rect 16739 5409 16797 5443
rect 16831 5409 16889 5443
rect 16923 5409 16981 5443
rect 17015 5409 17073 5443
rect 17107 5409 17165 5443
rect 17199 5409 17257 5443
rect 17291 5409 17349 5443
rect 17383 5409 17441 5443
rect 17475 5409 17504 5443
rect 7948 5211 8028 5249
rect 7948 5177 7994 5211
rect 7948 5121 8028 5177
rect 8063 5159 8097 5281
rect 8185 5227 8224 5257
rect 8185 5193 8219 5227
rect 8258 5223 8269 5257
rect 8605 5243 8639 5296
rect 8253 5193 8269 5223
rect 8315 5227 8572 5243
rect 8349 5209 8572 5227
rect 8606 5209 8639 5243
rect 8684 5257 8756 5259
rect 8718 5243 8756 5257
rect 8684 5209 8689 5223
rect 8723 5209 8756 5243
rect 8349 5193 8365 5209
rect 8684 5193 8756 5209
rect 8804 5227 8838 5296
rect 8872 5325 8950 5340
rect 9148 5331 9214 5347
rect 9148 5325 9180 5331
rect 8906 5324 8950 5325
rect 8906 5291 8916 5324
rect 8872 5290 8916 5291
rect 8872 5274 8950 5290
rect 8988 5291 9012 5325
rect 9046 5291 9062 5325
rect 9182 5291 9214 5297
rect 8988 5227 9022 5291
rect 9180 5281 9214 5291
rect 9259 5331 9310 5347
rect 9259 5297 9276 5331
rect 9259 5281 9310 5297
rect 8804 5193 9022 5227
rect 9090 5223 9136 5257
rect 9056 5220 9136 5223
rect 9259 5221 9293 5281
rect 9344 5249 9379 5380
rect 18302 5379 18331 5413
rect 18365 5379 18423 5413
rect 18457 5379 18515 5413
rect 18549 5379 18607 5413
rect 18641 5379 18699 5413
rect 18733 5379 18791 5413
rect 18825 5379 18883 5413
rect 18917 5379 18975 5413
rect 19009 5379 19067 5413
rect 19101 5379 19159 5413
rect 19193 5379 19222 5413
rect 8315 5190 8365 5193
rect 8063 5125 8196 5159
rect 8315 5156 8322 5190
rect 8356 5156 8365 5190
rect 9056 5186 9102 5220
rect 9056 5170 9136 5186
rect 8315 5155 8365 5156
rect 7948 5087 7994 5121
rect 8162 5121 8196 5125
rect 8446 5125 8648 5159
rect 8162 5103 8379 5121
rect 7948 5053 8028 5087
rect 8062 5057 8078 5091
rect 8112 5057 8128 5091
rect 8062 5019 8128 5057
rect 8162 5069 8345 5103
rect 8162 5053 8379 5069
rect 8446 5108 8480 5125
rect 8614 5108 8648 5125
rect 8446 5053 8480 5074
rect 8514 5057 8530 5091
rect 8564 5057 8580 5091
rect 8514 5019 8580 5057
rect 8789 5125 9004 5159
rect 9175 5157 9293 5221
rect 9327 5208 9379 5249
rect 18374 5322 18423 5338
rect 18374 5288 18383 5322
rect 18417 5288 18423 5322
rect 18374 5217 18423 5288
rect 18467 5322 18569 5379
rect 18501 5288 18535 5322
rect 18467 5272 18569 5288
rect 18605 5222 18643 5345
rect 9361 5184 9379 5208
rect 9175 5133 9209 5157
rect 8789 5108 8836 5125
rect 8614 5053 8648 5074
rect 8682 5061 8698 5095
rect 8732 5061 8748 5095
rect 8682 5019 8748 5061
rect 8789 5074 8802 5108
rect 8970 5108 9004 5125
rect 8789 5053 8836 5074
rect 8870 5057 8886 5091
rect 8920 5057 8936 5091
rect 8870 5019 8936 5057
rect 8970 5053 9004 5074
rect 9054 5108 9209 5133
rect 9327 5148 9338 5174
rect 9372 5148 9379 5184
rect 9088 5074 9209 5108
rect 9054 5053 9209 5074
rect 9243 5099 9293 5116
rect 9277 5065 9293 5099
rect 9243 5019 9293 5065
rect 9327 5114 9379 5148
rect 9361 5080 9379 5114
rect 18319 5183 18515 5217
rect 18549 5183 18565 5217
rect 18605 5188 18608 5222
rect 18642 5188 18643 5222
rect 9327 5053 9379 5080
rect 10046 5077 10075 5111
rect 10109 5077 10167 5111
rect 10201 5077 10259 5111
rect 10293 5077 10351 5111
rect 10385 5077 10443 5111
rect 10477 5077 10535 5111
rect 10569 5077 10627 5111
rect 10661 5077 10719 5111
rect 10753 5077 10811 5111
rect 10845 5077 10903 5111
rect 10937 5077 10995 5111
rect 11029 5077 11087 5111
rect 11121 5077 11179 5111
rect 11213 5077 11271 5111
rect 11305 5077 11363 5111
rect 11397 5077 11455 5111
rect 11489 5077 11547 5111
rect 11581 5077 11610 5111
rect 3880 4979 3909 5013
rect 3943 4979 3999 5013
rect 4033 4979 4091 5013
rect 4125 4979 4183 5013
rect 4217 4979 4275 5013
rect 4309 4979 4367 5013
rect 4401 4979 4459 5013
rect 4493 4979 4551 5013
rect 4585 4979 4643 5013
rect 4677 4979 4735 5013
rect 4769 4979 4827 5013
rect 4861 4979 4919 5013
rect 4953 4979 5011 5013
rect 5045 4979 5103 5013
rect 5137 4979 5195 5013
rect 5229 4979 5287 5013
rect 5321 4979 5379 5013
rect 5413 4979 5442 5013
rect 5830 4979 5859 5013
rect 5893 4979 5951 5013
rect 5985 4979 6043 5013
rect 6077 4979 6135 5013
rect 6169 4979 6227 5013
rect 6261 4979 6319 5013
rect 6353 4979 6411 5013
rect 6445 4979 6503 5013
rect 6537 4979 6595 5013
rect 6629 4979 6687 5013
rect 6721 4979 6779 5013
rect 6813 4979 6871 5013
rect 6905 4979 6963 5013
rect 6997 4979 7055 5013
rect 7089 4979 7147 5013
rect 7181 4979 7239 5013
rect 7273 4979 7331 5013
rect 7365 4979 7394 5013
rect 7832 4985 7861 5019
rect 7895 4985 7953 5019
rect 7987 4985 8045 5019
rect 8079 4985 8137 5019
rect 8171 4985 8229 5019
rect 8263 4985 8321 5019
rect 8355 4985 8413 5019
rect 8447 4985 8505 5019
rect 8539 4985 8597 5019
rect 8631 4985 8689 5019
rect 8723 4985 8781 5019
rect 8815 4985 8873 5019
rect 8907 4985 8965 5019
rect 8999 4985 9057 5019
rect 9091 4985 9149 5019
rect 9183 4985 9241 5019
rect 9275 4985 9333 5019
rect 9367 4985 9396 5019
rect 10070 4999 10150 5043
rect 10199 5039 10265 5077
rect 10199 5005 10215 5039
rect 10249 5005 10265 5039
rect 10299 5027 10501 5043
rect 10070 4965 10116 4999
rect 10299 4993 10467 5027
rect 10299 4971 10333 4993
rect 10467 4975 10501 4993
rect 10568 5022 10602 5043
rect 10636 5039 10702 5077
rect 10636 5005 10652 5039
rect 10686 5005 10702 5039
rect 10736 5022 10770 5043
rect 10070 4932 10150 4965
rect 10185 4937 10333 4971
rect 10568 4971 10602 4988
rect 10804 5030 10870 5077
rect 10804 4996 10820 5030
rect 10854 4996 10870 5030
rect 10924 5022 10958 5043
rect 10736 4971 10770 4988
rect 10070 4797 10136 4932
rect 10185 4895 10219 4937
rect 10170 4879 10219 4895
rect 10426 4907 10438 4941
rect 10472 4907 10525 4941
rect 10568 4937 10770 4971
rect 10992 5039 11058 5077
rect 10992 5005 11008 5039
rect 11042 5005 11058 5039
rect 11092 5022 11126 5043
rect 10924 4971 10958 4988
rect 11092 4971 11126 4988
rect 10924 4937 11126 4971
rect 11176 5022 11296 5043
rect 11210 4988 11296 5022
rect 11349 5035 11415 5077
rect 11349 5001 11365 5035
rect 11399 5001 11415 5035
rect 11176 4967 11296 4988
rect 11449 4999 11501 5043
rect 11176 4941 11415 4967
rect 11176 4907 11178 4941
rect 11212 4933 11415 4941
rect 11212 4907 11224 4933
rect 10426 4903 10525 4907
rect 10204 4845 10219 4879
rect 10170 4829 10219 4845
rect 10253 4873 10269 4887
rect 10253 4839 10254 4873
rect 10303 4853 10341 4887
rect 10426 4869 10509 4903
rect 10543 4869 10559 4903
rect 10593 4869 10609 4903
rect 10643 4873 10668 4903
rect 10288 4839 10341 4853
rect 10593 4839 10622 4869
rect 10656 4839 10668 4873
rect 10727 4844 10960 4901
rect 11381 4895 11415 4933
rect 11483 4965 11501 4999
rect 11449 4928 11501 4965
rect 11535 4983 11593 5077
rect 12228 5033 12257 5067
rect 12291 5033 12345 5067
rect 12379 5033 12437 5067
rect 12471 5033 12529 5067
rect 12563 5033 12621 5067
rect 12655 5033 12713 5067
rect 12747 5033 12805 5067
rect 12839 5033 12897 5067
rect 12931 5033 12989 5067
rect 13023 5033 13081 5067
rect 13115 5033 13173 5067
rect 13207 5033 13265 5067
rect 13299 5033 13357 5067
rect 13391 5033 13449 5067
rect 13483 5033 13541 5067
rect 13575 5033 13633 5067
rect 13667 5033 13725 5067
rect 13759 5033 13788 5067
rect 11535 4949 11547 4983
rect 11581 4949 11593 4983
rect 11535 4932 11593 4949
rect 12245 4939 12303 5033
rect 10070 4759 10150 4797
rect 10070 4725 10116 4759
rect 10070 4669 10150 4725
rect 10185 4707 10219 4829
rect 10307 4775 10346 4805
rect 10307 4741 10341 4775
rect 10380 4771 10391 4805
rect 10727 4791 10761 4844
rect 10375 4741 10391 4771
rect 10437 4775 10694 4791
rect 10471 4757 10694 4775
rect 10728 4757 10761 4791
rect 10806 4805 10878 4807
rect 10840 4791 10878 4805
rect 10806 4757 10811 4771
rect 10845 4757 10878 4791
rect 10471 4741 10487 4757
rect 10806 4741 10878 4757
rect 10926 4775 10960 4844
rect 10994 4873 11072 4888
rect 11270 4879 11336 4895
rect 11270 4873 11302 4879
rect 11028 4872 11072 4873
rect 11028 4839 11038 4872
rect 10994 4838 11038 4839
rect 10994 4822 11072 4838
rect 11110 4839 11134 4873
rect 11168 4839 11184 4873
rect 11304 4839 11336 4845
rect 11110 4775 11144 4839
rect 11302 4829 11336 4839
rect 11381 4879 11432 4895
rect 11381 4845 11398 4879
rect 11381 4829 11432 4845
rect 10926 4741 11144 4775
rect 11212 4771 11258 4805
rect 11178 4768 11258 4771
rect 11381 4769 11415 4829
rect 11466 4797 11501 4928
rect 12245 4905 12257 4939
rect 12291 4905 12303 4939
rect 12245 4888 12303 4905
rect 12340 4955 12420 4999
rect 12469 4995 12535 5033
rect 12469 4961 12485 4995
rect 12519 4961 12535 4995
rect 12569 4983 12771 4999
rect 12340 4921 12386 4955
rect 12569 4949 12737 4983
rect 12569 4927 12603 4949
rect 12737 4931 12771 4949
rect 12838 4978 12872 4999
rect 12906 4995 12972 5033
rect 12906 4961 12922 4995
rect 12956 4961 12972 4995
rect 13006 4978 13040 4999
rect 12340 4888 12420 4921
rect 12455 4893 12603 4927
rect 12838 4927 12872 4944
rect 13074 4986 13140 5033
rect 13074 4952 13090 4986
rect 13124 4952 13140 4986
rect 13194 4978 13228 4999
rect 13006 4927 13040 4944
rect 10437 4740 10487 4741
rect 10185 4673 10318 4707
rect 10437 4706 10446 4740
rect 10480 4706 10487 4740
rect 11178 4734 11224 4768
rect 11178 4718 11258 4734
rect 10437 4703 10487 4706
rect 10070 4635 10116 4669
rect 10284 4669 10318 4673
rect 10568 4673 10770 4707
rect 10284 4651 10501 4669
rect 10070 4601 10150 4635
rect 10184 4605 10200 4639
rect 10234 4605 10250 4639
rect 10184 4567 10250 4605
rect 10284 4617 10467 4651
rect 10284 4601 10501 4617
rect 10568 4656 10602 4673
rect 10736 4656 10770 4673
rect 10568 4601 10602 4622
rect 10636 4605 10652 4639
rect 10686 4605 10702 4639
rect 10636 4567 10702 4605
rect 10911 4673 11126 4707
rect 11297 4705 11415 4769
rect 11449 4756 11501 4797
rect 11483 4732 11501 4756
rect 11297 4681 11331 4705
rect 10911 4656 10958 4673
rect 10736 4601 10770 4622
rect 10804 4609 10820 4643
rect 10854 4609 10870 4643
rect 10804 4567 10870 4609
rect 10911 4622 10924 4656
rect 11092 4656 11126 4673
rect 10911 4601 10958 4622
rect 10992 4605 11008 4639
rect 11042 4605 11058 4639
rect 10992 4567 11058 4605
rect 11092 4601 11126 4622
rect 11176 4656 11331 4681
rect 11449 4696 11454 4722
rect 11494 4696 11501 4732
rect 11210 4622 11331 4656
rect 11176 4601 11331 4622
rect 11365 4647 11415 4664
rect 11399 4613 11415 4647
rect 11365 4567 11415 4613
rect 11449 4662 11501 4696
rect 11483 4628 11501 4662
rect 11449 4601 11501 4628
rect 11535 4765 11593 4800
rect 11535 4731 11547 4765
rect 11581 4731 11593 4765
rect 11535 4672 11593 4731
rect 11535 4638 11547 4672
rect 11581 4638 11593 4672
rect 11535 4567 11593 4638
rect 12245 4721 12303 4756
rect 12245 4687 12257 4721
rect 12291 4687 12303 4721
rect 12245 4628 12303 4687
rect 12245 4594 12257 4628
rect 12291 4594 12303 4628
rect 10046 4533 10075 4567
rect 10109 4533 10167 4567
rect 10201 4533 10259 4567
rect 10293 4533 10351 4567
rect 10385 4533 10443 4567
rect 10477 4533 10535 4567
rect 10569 4533 10627 4567
rect 10661 4533 10719 4567
rect 10753 4533 10811 4567
rect 10845 4533 10903 4567
rect 10937 4533 10995 4567
rect 11029 4533 11087 4567
rect 11121 4533 11179 4567
rect 11213 4533 11271 4567
rect 11305 4533 11363 4567
rect 11397 4533 11455 4567
rect 11489 4533 11547 4567
rect 11581 4533 11610 4567
rect 12245 4523 12303 4594
rect 12340 4753 12406 4888
rect 12455 4851 12489 4893
rect 12440 4835 12489 4851
rect 12696 4863 12708 4897
rect 12742 4863 12795 4897
rect 12838 4893 13040 4927
rect 13262 4995 13328 5033
rect 13262 4961 13278 4995
rect 13312 4961 13328 4995
rect 13362 4978 13396 4999
rect 13194 4927 13228 4944
rect 13362 4927 13396 4944
rect 13194 4893 13396 4927
rect 13446 4978 13566 4999
rect 13480 4944 13566 4978
rect 13619 4991 13685 5033
rect 14228 5027 14257 5061
rect 14291 5027 14347 5061
rect 14381 5027 14439 5061
rect 14473 5027 14531 5061
rect 14565 5027 14623 5061
rect 14657 5027 14715 5061
rect 14749 5027 14807 5061
rect 14841 5027 14899 5061
rect 14933 5027 14991 5061
rect 15025 5027 15083 5061
rect 15117 5027 15175 5061
rect 15209 5027 15267 5061
rect 15301 5027 15359 5061
rect 15393 5027 15451 5061
rect 15485 5027 15543 5061
rect 15577 5027 15635 5061
rect 15669 5027 15727 5061
rect 15761 5027 15790 5061
rect 13619 4957 13635 4991
rect 13669 4957 13685 4991
rect 13446 4923 13566 4944
rect 13719 4955 13771 4999
rect 13446 4897 13685 4923
rect 13446 4863 13448 4897
rect 13482 4889 13685 4897
rect 13482 4863 13494 4889
rect 12696 4859 12795 4863
rect 12474 4801 12489 4835
rect 12440 4785 12489 4801
rect 12523 4829 12539 4843
rect 12523 4795 12524 4829
rect 12573 4809 12611 4843
rect 12696 4825 12779 4859
rect 12813 4825 12829 4859
rect 12863 4825 12879 4859
rect 12913 4829 12938 4859
rect 12558 4795 12611 4809
rect 12863 4795 12892 4825
rect 12926 4795 12938 4829
rect 12997 4800 13230 4857
rect 13651 4851 13685 4889
rect 13753 4921 13771 4955
rect 13719 4884 13771 4921
rect 12340 4715 12420 4753
rect 12340 4681 12386 4715
rect 12340 4625 12420 4681
rect 12455 4663 12489 4785
rect 12577 4731 12616 4761
rect 12577 4697 12611 4731
rect 12650 4727 12661 4761
rect 12997 4747 13031 4800
rect 12645 4697 12661 4727
rect 12707 4731 12964 4747
rect 12741 4713 12964 4731
rect 12998 4713 13031 4747
rect 13076 4761 13148 4763
rect 13110 4747 13148 4761
rect 13076 4713 13081 4727
rect 13115 4713 13148 4747
rect 12741 4697 12757 4713
rect 13076 4697 13148 4713
rect 13196 4731 13230 4800
rect 13264 4829 13342 4844
rect 13540 4835 13606 4851
rect 13540 4829 13572 4835
rect 13298 4828 13342 4829
rect 13298 4795 13308 4828
rect 13264 4794 13308 4795
rect 13264 4778 13342 4794
rect 13380 4795 13404 4829
rect 13438 4795 13454 4829
rect 13574 4795 13606 4801
rect 13380 4731 13414 4795
rect 13572 4785 13606 4795
rect 13651 4835 13702 4851
rect 13651 4801 13668 4835
rect 13651 4785 13702 4801
rect 13196 4697 13414 4731
rect 13482 4727 13528 4761
rect 13448 4724 13528 4727
rect 13651 4725 13685 4785
rect 13736 4753 13771 4884
rect 14245 4933 14303 5027
rect 14245 4899 14257 4933
rect 14291 4899 14303 4933
rect 14245 4882 14303 4899
rect 14342 4949 14422 4993
rect 14471 4989 14537 5027
rect 14471 4955 14487 4989
rect 14521 4955 14537 4989
rect 14571 4977 14773 4993
rect 14342 4915 14388 4949
rect 14571 4943 14739 4977
rect 14571 4921 14605 4943
rect 14739 4925 14773 4943
rect 14840 4972 14874 4993
rect 14908 4989 14974 5027
rect 14908 4955 14924 4989
rect 14958 4955 14974 4989
rect 15008 4972 15042 4993
rect 14342 4882 14422 4915
rect 14457 4887 14605 4921
rect 14840 4921 14874 4938
rect 15076 4980 15142 5027
rect 15076 4946 15092 4980
rect 15126 4946 15142 4980
rect 15196 4972 15230 4993
rect 15008 4921 15042 4938
rect 12707 4694 12757 4697
rect 12455 4629 12588 4663
rect 12707 4660 12714 4694
rect 12748 4660 12757 4694
rect 13448 4690 13494 4724
rect 13448 4674 13528 4690
rect 12707 4659 12757 4660
rect 12340 4591 12386 4625
rect 12554 4625 12588 4629
rect 12838 4629 13040 4663
rect 12554 4607 12771 4625
rect 12340 4557 12420 4591
rect 12454 4561 12470 4595
rect 12504 4561 12520 4595
rect 12454 4523 12520 4561
rect 12554 4573 12737 4607
rect 12554 4557 12771 4573
rect 12838 4612 12872 4629
rect 13006 4612 13040 4629
rect 12838 4557 12872 4578
rect 12906 4561 12922 4595
rect 12956 4561 12972 4595
rect 12906 4523 12972 4561
rect 13181 4629 13396 4663
rect 13567 4661 13685 4725
rect 13719 4712 13771 4753
rect 13753 4688 13771 4712
rect 13567 4637 13601 4661
rect 13181 4612 13228 4629
rect 13006 4557 13040 4578
rect 13074 4565 13090 4599
rect 13124 4565 13140 4599
rect 13074 4523 13140 4565
rect 13181 4578 13194 4612
rect 13362 4612 13396 4629
rect 13181 4557 13228 4578
rect 13262 4561 13278 4595
rect 13312 4561 13328 4595
rect 13262 4523 13328 4561
rect 13362 4557 13396 4578
rect 13446 4612 13601 4637
rect 13719 4652 13730 4678
rect 13764 4652 13771 4688
rect 13480 4578 13601 4612
rect 13446 4557 13601 4578
rect 13635 4603 13685 4620
rect 13669 4569 13685 4603
rect 13635 4523 13685 4569
rect 13719 4618 13771 4652
rect 13753 4584 13771 4618
rect 13719 4557 13771 4584
rect 14245 4715 14303 4750
rect 14245 4681 14257 4715
rect 14291 4681 14303 4715
rect 14245 4622 14303 4681
rect 14245 4588 14257 4622
rect 14291 4588 14303 4622
rect 12228 4489 12257 4523
rect 12291 4489 12345 4523
rect 12379 4489 12437 4523
rect 12471 4489 12529 4523
rect 12563 4489 12621 4523
rect 12655 4489 12713 4523
rect 12747 4489 12805 4523
rect 12839 4489 12897 4523
rect 12931 4489 12989 4523
rect 13023 4489 13081 4523
rect 13115 4489 13173 4523
rect 13207 4489 13265 4523
rect 13299 4489 13357 4523
rect 13391 4489 13449 4523
rect 13483 4489 13541 4523
rect 13575 4489 13633 4523
rect 13667 4489 13725 4523
rect 13759 4489 13788 4523
rect 14245 4517 14303 4588
rect 14342 4747 14408 4882
rect 14457 4845 14491 4887
rect 14442 4829 14491 4845
rect 14698 4857 14710 4891
rect 14744 4857 14797 4891
rect 14840 4887 15042 4921
rect 15264 4989 15330 5027
rect 15264 4955 15280 4989
rect 15314 4955 15330 4989
rect 15364 4972 15398 4993
rect 15196 4921 15230 4938
rect 15364 4921 15398 4938
rect 15196 4887 15398 4921
rect 15448 4972 15568 4993
rect 15482 4938 15568 4972
rect 15621 4985 15687 5027
rect 16252 5009 16281 5043
rect 16315 5009 16369 5043
rect 16403 5009 16461 5043
rect 16495 5009 16553 5043
rect 16587 5009 16645 5043
rect 16679 5009 16737 5043
rect 16771 5009 16829 5043
rect 16863 5009 16921 5043
rect 16955 5009 17013 5043
rect 17047 5009 17105 5043
rect 17139 5009 17197 5043
rect 17231 5009 17289 5043
rect 17323 5009 17381 5043
rect 17415 5009 17473 5043
rect 17507 5009 17565 5043
rect 17599 5009 17657 5043
rect 17691 5009 17749 5043
rect 17783 5009 17812 5043
rect 18319 5021 18387 5183
rect 18421 5070 18432 5108
rect 18470 5104 18571 5108
rect 18471 5070 18571 5104
rect 15621 4951 15637 4985
rect 15671 4951 15687 4985
rect 15448 4917 15568 4938
rect 15721 4949 15773 4993
rect 15448 4891 15687 4917
rect 15448 4857 15450 4891
rect 15484 4883 15687 4891
rect 15484 4857 15496 4883
rect 14698 4853 14797 4857
rect 14476 4795 14491 4829
rect 14442 4779 14491 4795
rect 14525 4823 14541 4837
rect 14525 4789 14526 4823
rect 14575 4803 14613 4837
rect 14698 4819 14781 4853
rect 14815 4819 14831 4853
rect 14865 4819 14881 4853
rect 14915 4823 14940 4853
rect 14560 4789 14613 4803
rect 14865 4789 14894 4819
rect 14928 4789 14940 4823
rect 14999 4794 15232 4851
rect 15653 4845 15687 4883
rect 15755 4915 15773 4949
rect 15721 4878 15773 4915
rect 14342 4709 14422 4747
rect 14342 4675 14388 4709
rect 14342 4619 14422 4675
rect 14457 4657 14491 4779
rect 14579 4725 14618 4755
rect 14579 4691 14613 4725
rect 14652 4721 14663 4755
rect 14999 4741 15033 4794
rect 14647 4691 14663 4721
rect 14709 4725 14966 4741
rect 14743 4707 14966 4725
rect 15000 4707 15033 4741
rect 15078 4755 15150 4757
rect 15112 4741 15150 4755
rect 15078 4707 15083 4721
rect 15117 4707 15150 4741
rect 14743 4691 14759 4707
rect 15078 4691 15150 4707
rect 15198 4725 15232 4794
rect 15266 4823 15344 4838
rect 15542 4829 15608 4845
rect 15542 4823 15574 4829
rect 15300 4822 15344 4823
rect 15300 4789 15310 4822
rect 15266 4788 15310 4789
rect 15266 4772 15344 4788
rect 15382 4789 15406 4823
rect 15440 4789 15456 4823
rect 15576 4789 15608 4795
rect 15382 4725 15416 4789
rect 15574 4779 15608 4789
rect 15653 4829 15704 4845
rect 15653 4795 15670 4829
rect 15653 4779 15704 4795
rect 15198 4691 15416 4725
rect 15484 4721 15530 4755
rect 15450 4718 15530 4721
rect 15653 4719 15687 4779
rect 15738 4747 15773 4878
rect 16269 4915 16327 5009
rect 16269 4881 16281 4915
rect 16315 4881 16327 4915
rect 16269 4864 16327 4881
rect 16364 4931 16444 4975
rect 16493 4971 16559 5009
rect 16493 4937 16509 4971
rect 16543 4937 16559 4971
rect 16593 4959 16795 4975
rect 16364 4897 16410 4931
rect 16593 4925 16761 4959
rect 16593 4903 16627 4925
rect 16761 4907 16795 4925
rect 16862 4954 16896 4975
rect 16930 4971 16996 5009
rect 16930 4937 16946 4971
rect 16980 4937 16996 4971
rect 17030 4954 17064 4975
rect 16364 4864 16444 4897
rect 16479 4869 16627 4903
rect 16862 4903 16896 4920
rect 17098 4962 17164 5009
rect 17098 4928 17114 4962
rect 17148 4928 17164 4962
rect 17218 4954 17252 4975
rect 17030 4903 17064 4920
rect 14709 4688 14759 4691
rect 14457 4623 14590 4657
rect 14709 4654 14716 4688
rect 14750 4654 14759 4688
rect 15450 4684 15496 4718
rect 15450 4668 15530 4684
rect 14709 4653 14759 4654
rect 14342 4585 14388 4619
rect 14556 4619 14590 4623
rect 14840 4623 15042 4657
rect 14556 4601 14773 4619
rect 14342 4551 14422 4585
rect 14456 4555 14472 4589
rect 14506 4555 14522 4589
rect 14456 4517 14522 4555
rect 14556 4567 14739 4601
rect 14556 4551 14773 4567
rect 14840 4606 14874 4623
rect 15008 4606 15042 4623
rect 14840 4551 14874 4572
rect 14908 4555 14924 4589
rect 14958 4555 14974 4589
rect 14908 4517 14974 4555
rect 15183 4623 15398 4657
rect 15569 4655 15687 4719
rect 15721 4706 15773 4747
rect 15755 4682 15773 4706
rect 15569 4631 15603 4655
rect 15183 4606 15230 4623
rect 15008 4551 15042 4572
rect 15076 4559 15092 4593
rect 15126 4559 15142 4593
rect 15076 4517 15142 4559
rect 15183 4572 15196 4606
rect 15364 4606 15398 4623
rect 15183 4551 15230 4572
rect 15264 4555 15280 4589
rect 15314 4555 15330 4589
rect 15264 4517 15330 4555
rect 15364 4551 15398 4572
rect 15448 4606 15603 4631
rect 15721 4646 15732 4672
rect 15766 4646 15773 4682
rect 15482 4572 15603 4606
rect 15448 4551 15603 4572
rect 15637 4597 15687 4614
rect 15671 4563 15687 4597
rect 15637 4517 15687 4563
rect 15721 4612 15773 4646
rect 15755 4578 15773 4612
rect 15721 4551 15773 4578
rect 16269 4697 16327 4732
rect 16269 4663 16281 4697
rect 16315 4663 16327 4697
rect 16269 4604 16327 4663
rect 16269 4570 16281 4604
rect 16315 4570 16327 4604
rect 14228 4483 14257 4517
rect 14291 4483 14347 4517
rect 14381 4483 14439 4517
rect 14473 4483 14531 4517
rect 14565 4483 14623 4517
rect 14657 4483 14715 4517
rect 14749 4483 14807 4517
rect 14841 4483 14899 4517
rect 14933 4483 14991 4517
rect 15025 4483 15083 4517
rect 15117 4483 15175 4517
rect 15209 4483 15267 4517
rect 15301 4483 15359 4517
rect 15393 4483 15451 4517
rect 15485 4483 15543 4517
rect 15577 4483 15635 4517
rect 15669 4483 15727 4517
rect 15761 4483 15790 4517
rect 16269 4499 16327 4570
rect 16364 4729 16430 4864
rect 16479 4827 16513 4869
rect 16464 4811 16513 4827
rect 16720 4839 16732 4873
rect 16766 4839 16819 4873
rect 16862 4869 17064 4903
rect 17286 4971 17352 5009
rect 17286 4937 17302 4971
rect 17336 4937 17352 4971
rect 17386 4954 17420 4975
rect 17218 4903 17252 4920
rect 17386 4903 17420 4920
rect 17218 4869 17420 4903
rect 17470 4954 17590 4975
rect 17504 4920 17590 4954
rect 17643 4967 17709 5009
rect 18319 5005 18422 5021
rect 17643 4933 17659 4967
rect 17693 4933 17709 4967
rect 17470 4899 17590 4920
rect 17743 4931 17795 4975
rect 18319 4971 18383 5005
rect 18417 4971 18422 5005
rect 18319 4939 18422 4971
rect 18469 5005 18503 5021
rect 17470 4873 17709 4899
rect 17470 4839 17472 4873
rect 17506 4865 17709 4873
rect 17506 4839 17518 4865
rect 16720 4835 16819 4839
rect 16498 4777 16513 4811
rect 16464 4761 16513 4777
rect 16547 4805 16563 4819
rect 16547 4771 16548 4805
rect 16597 4785 16635 4819
rect 16720 4801 16803 4835
rect 16837 4801 16853 4835
rect 16887 4801 16903 4835
rect 16937 4805 16962 4835
rect 16582 4771 16635 4785
rect 16887 4771 16916 4801
rect 16950 4771 16962 4805
rect 17021 4776 17254 4833
rect 17675 4827 17709 4865
rect 17777 4897 17795 4931
rect 17743 4860 17795 4897
rect 18469 4869 18503 4971
rect 18537 4937 18571 5070
rect 18605 5104 18643 5188
rect 18677 5217 18732 5345
rect 18770 5322 18876 5345
rect 18804 5288 18876 5322
rect 18961 5337 19027 5379
rect 18961 5303 18977 5337
rect 19011 5303 19027 5337
rect 18961 5299 19027 5303
rect 19061 5318 19112 5345
rect 18770 5272 18876 5288
rect 18841 5265 18876 5272
rect 19095 5284 19112 5318
rect 18711 5194 18732 5217
rect 18677 5160 18690 5183
rect 18724 5160 18732 5194
rect 18677 5113 18732 5160
rect 18773 5217 18807 5233
rect 18639 5073 18643 5104
rect 18773 5073 18807 5183
rect 18639 5070 18807 5073
rect 18605 5039 18807 5070
rect 18841 5231 19027 5265
rect 19061 5231 19112 5284
rect 19147 5285 19205 5379
rect 19147 5251 19159 5285
rect 19193 5251 19205 5285
rect 19147 5234 19205 5251
rect 18841 5005 18875 5231
rect 18993 5197 19027 5231
rect 18650 4971 18666 5005
rect 18700 4971 18741 5005
rect 18775 4971 18875 5005
rect 18909 5181 18948 5197
rect 18909 5147 18914 5181
rect 18909 5131 18948 5147
rect 18993 5181 19044 5197
rect 18993 5147 19010 5181
rect 18993 5131 19044 5147
rect 18909 4937 18943 5131
rect 19078 5097 19112 5231
rect 18537 4903 18943 4937
rect 18977 5081 19011 5097
rect 18977 5013 19011 5047
rect 18977 4945 19011 4979
rect 18977 4869 19011 4911
rect 19045 5081 19112 5097
rect 19045 5047 19061 5081
rect 19095 5047 19112 5081
rect 19045 5042 19112 5047
rect 19045 5013 19064 5042
rect 19045 4979 19061 5013
rect 19102 5004 19112 5042
rect 19095 4979 19112 5004
rect 19045 4945 19112 4979
rect 19045 4911 19061 4945
rect 19095 4911 19112 4945
rect 19045 4903 19112 4911
rect 19147 5067 19205 5102
rect 19147 5033 19159 5067
rect 19193 5033 19205 5067
rect 19147 4974 19205 5033
rect 19147 4940 19159 4974
rect 19193 4940 19205 4974
rect 19147 4869 19205 4940
rect 16364 4691 16444 4729
rect 16364 4657 16410 4691
rect 16364 4601 16444 4657
rect 16479 4639 16513 4761
rect 16601 4707 16640 4737
rect 16601 4673 16635 4707
rect 16674 4703 16685 4737
rect 17021 4723 17055 4776
rect 16669 4673 16685 4703
rect 16731 4707 16988 4723
rect 16765 4689 16988 4707
rect 17022 4689 17055 4723
rect 17100 4737 17172 4739
rect 17134 4723 17172 4737
rect 17100 4689 17105 4703
rect 17139 4689 17172 4723
rect 16765 4673 16781 4689
rect 17100 4673 17172 4689
rect 17220 4707 17254 4776
rect 17288 4805 17366 4820
rect 17564 4811 17630 4827
rect 17564 4805 17596 4811
rect 17322 4804 17366 4805
rect 17322 4771 17332 4804
rect 17288 4770 17332 4771
rect 17288 4754 17366 4770
rect 17404 4771 17428 4805
rect 17462 4771 17478 4805
rect 17598 4771 17630 4777
rect 17404 4707 17438 4771
rect 17596 4761 17630 4771
rect 17675 4811 17726 4827
rect 17675 4777 17692 4811
rect 17675 4761 17726 4777
rect 17220 4673 17438 4707
rect 17506 4703 17552 4737
rect 17472 4700 17552 4703
rect 17675 4701 17709 4761
rect 17760 4729 17795 4860
rect 18302 4835 18331 4869
rect 18365 4835 18423 4869
rect 18457 4835 18515 4869
rect 18549 4835 18607 4869
rect 18641 4835 18699 4869
rect 18733 4835 18791 4869
rect 18825 4835 18883 4869
rect 18917 4835 18975 4869
rect 19009 4835 19067 4869
rect 19101 4835 19159 4869
rect 19193 4835 19222 4869
rect 16731 4670 16781 4673
rect 16479 4605 16612 4639
rect 16731 4636 16738 4670
rect 16772 4636 16781 4670
rect 17472 4666 17518 4700
rect 17472 4650 17552 4666
rect 16731 4635 16781 4636
rect 16364 4567 16410 4601
rect 16578 4601 16612 4605
rect 16862 4605 17064 4639
rect 16578 4583 16795 4601
rect 16364 4533 16444 4567
rect 16478 4537 16494 4571
rect 16528 4537 16544 4571
rect 16478 4499 16544 4537
rect 16578 4549 16761 4583
rect 16578 4533 16795 4549
rect 16862 4588 16896 4605
rect 17030 4588 17064 4605
rect 16862 4533 16896 4554
rect 16930 4537 16946 4571
rect 16980 4537 16996 4571
rect 16930 4499 16996 4537
rect 17205 4605 17420 4639
rect 17591 4637 17709 4701
rect 17743 4688 17795 4729
rect 17777 4664 17795 4688
rect 17591 4613 17625 4637
rect 17205 4588 17252 4605
rect 17030 4533 17064 4554
rect 17098 4541 17114 4575
rect 17148 4541 17164 4575
rect 17098 4499 17164 4541
rect 17205 4554 17218 4588
rect 17386 4588 17420 4605
rect 17205 4533 17252 4554
rect 17286 4537 17302 4571
rect 17336 4537 17352 4571
rect 17286 4499 17352 4537
rect 17386 4533 17420 4554
rect 17470 4588 17625 4613
rect 17743 4628 17754 4654
rect 17788 4628 17795 4664
rect 17504 4554 17625 4588
rect 17470 4533 17625 4554
rect 17659 4579 17709 4596
rect 17693 4545 17709 4579
rect 17659 4499 17709 4545
rect 17743 4594 17795 4628
rect 17777 4560 17795 4594
rect 17743 4533 17795 4560
rect 16252 4465 16281 4499
rect 16315 4465 16369 4499
rect 16403 4465 16461 4499
rect 16495 4465 16553 4499
rect 16587 4465 16645 4499
rect 16679 4465 16737 4499
rect 16771 4465 16829 4499
rect 16863 4465 16921 4499
rect 16955 4465 17013 4499
rect 17047 4465 17105 4499
rect 17139 4465 17197 4499
rect 17231 4465 17289 4499
rect 17323 4465 17381 4499
rect 17415 4465 17473 4499
rect 17507 4465 17565 4499
rect 17599 4465 17657 4499
rect 17691 4465 17749 4499
rect 17783 4465 17812 4499
rect 5994 3323 6023 3357
rect 6057 3323 6111 3357
rect 6145 3323 6203 3357
rect 6237 3323 6295 3357
rect 6329 3323 6358 3357
rect 6011 3229 6069 3323
rect 6011 3195 6023 3229
rect 6057 3195 6069 3229
rect 6011 3178 6069 3195
rect 6148 3277 6214 3289
rect 6148 3243 6164 3277
rect 6198 3243 6214 3277
rect 6148 3209 6214 3243
rect 6148 3175 6164 3209
rect 6198 3175 6214 3209
rect 6148 3163 6214 3175
rect 6248 3277 6294 3323
rect 6282 3243 6294 3277
rect 6248 3209 6294 3243
rect 6282 3175 6294 3209
rect 6148 3122 6194 3163
rect 6248 3159 6294 3175
rect 6182 3088 6194 3122
rect 6011 3011 6069 3046
rect 6011 2977 6023 3011
rect 6057 2977 6069 3011
rect 6011 2918 6069 2977
rect 6011 2884 6023 2918
rect 6057 2884 6069 2918
rect 6011 2813 6069 2884
rect 6148 3043 6194 3088
rect 6228 3090 6244 3125
rect 6278 3090 6294 3125
rect 6228 3077 6294 3090
rect 6148 3025 6214 3043
rect 6148 2991 6164 3025
rect 6198 2991 6214 3025
rect 6148 2957 6214 2991
rect 6148 2923 6164 2957
rect 6198 2923 6214 2957
rect 6148 2889 6214 2923
rect 6148 2855 6164 2889
rect 6198 2855 6214 2889
rect 6148 2847 6214 2855
rect 6248 3025 6290 3041
rect 6282 2991 6290 3025
rect 6248 2957 6290 2991
rect 6282 2923 6290 2957
rect 6248 2889 6290 2923
rect 6282 2855 6290 2889
rect 6248 2813 6290 2855
rect 5994 2779 6023 2813
rect 6057 2779 6111 2813
rect 6145 2779 6203 2813
rect 6237 2779 6295 2813
rect 6329 2779 6358 2813
rect 1716 2271 1745 2305
rect 1779 2271 1835 2305
rect 1869 2271 1927 2305
rect 1961 2271 2019 2305
rect 2053 2271 2111 2305
rect 2145 2271 2203 2305
rect 2237 2271 2295 2305
rect 2329 2271 2387 2305
rect 2421 2271 2479 2305
rect 2513 2271 2571 2305
rect 2605 2271 2663 2305
rect 2697 2271 2755 2305
rect 2789 2271 2847 2305
rect 2881 2271 2939 2305
rect 2973 2271 3031 2305
rect 3065 2271 3123 2305
rect 3157 2271 3215 2305
rect 3249 2271 3278 2305
rect 1733 2177 1791 2271
rect 1733 2143 1745 2177
rect 1779 2143 1791 2177
rect 1733 2126 1791 2143
rect 1830 2193 1910 2237
rect 1959 2233 2025 2271
rect 1959 2199 1975 2233
rect 2009 2199 2025 2233
rect 2059 2221 2261 2237
rect 1830 2159 1876 2193
rect 2059 2187 2227 2221
rect 2059 2165 2093 2187
rect 2227 2169 2261 2187
rect 2328 2216 2362 2237
rect 2396 2233 2462 2271
rect 2396 2199 2412 2233
rect 2446 2199 2462 2233
rect 2496 2216 2530 2237
rect 1830 2126 1910 2159
rect 1945 2131 2093 2165
rect 2328 2165 2362 2182
rect 2564 2224 2630 2271
rect 2564 2190 2580 2224
rect 2614 2190 2630 2224
rect 2684 2216 2718 2237
rect 2496 2165 2530 2182
rect 1733 1959 1791 1994
rect 1733 1925 1745 1959
rect 1779 1925 1791 1959
rect 1733 1866 1791 1925
rect 1733 1832 1745 1866
rect 1779 1832 1791 1866
rect 1733 1761 1791 1832
rect 1830 1991 1896 2126
rect 1945 2089 1979 2131
rect 1930 2073 1979 2089
rect 2186 2101 2198 2135
rect 2232 2101 2285 2135
rect 2328 2131 2530 2165
rect 2752 2233 2818 2271
rect 2752 2199 2768 2233
rect 2802 2199 2818 2233
rect 2852 2216 2886 2237
rect 2684 2165 2718 2182
rect 2852 2165 2886 2182
rect 2684 2131 2886 2165
rect 2936 2216 3056 2237
rect 2970 2182 3056 2216
rect 3109 2229 3175 2271
rect 3786 2267 3815 2301
rect 3849 2267 3905 2301
rect 3939 2267 3997 2301
rect 4031 2267 4089 2301
rect 4123 2267 4181 2301
rect 4215 2267 4273 2301
rect 4307 2267 4365 2301
rect 4399 2267 4457 2301
rect 4491 2267 4549 2301
rect 4583 2267 4641 2301
rect 4675 2267 4733 2301
rect 4767 2267 4825 2301
rect 4859 2267 4917 2301
rect 4951 2267 5009 2301
rect 5043 2267 5101 2301
rect 5135 2267 5193 2301
rect 5227 2267 5285 2301
rect 5319 2267 5348 2301
rect 5742 2267 5771 2301
rect 5805 2267 5857 2301
rect 5891 2267 5949 2301
rect 5983 2267 6041 2301
rect 6075 2267 6133 2301
rect 6167 2267 6225 2301
rect 6259 2267 6317 2301
rect 6351 2267 6409 2301
rect 6443 2267 6501 2301
rect 6535 2267 6593 2301
rect 6627 2267 6685 2301
rect 6719 2267 6777 2301
rect 6811 2267 6869 2301
rect 6903 2267 6961 2301
rect 6995 2267 7053 2301
rect 7087 2267 7145 2301
rect 7179 2267 7237 2301
rect 7271 2267 7300 2301
rect 7740 2273 7769 2307
rect 7803 2273 7859 2307
rect 7893 2273 7951 2307
rect 7985 2273 8043 2307
rect 8077 2273 8135 2307
rect 8169 2273 8227 2307
rect 8261 2273 8319 2307
rect 8353 2273 8411 2307
rect 8445 2273 8503 2307
rect 8537 2273 8595 2307
rect 8629 2273 8687 2307
rect 8721 2273 8779 2307
rect 8813 2273 8871 2307
rect 8905 2273 8963 2307
rect 8997 2273 9055 2307
rect 9089 2273 9147 2307
rect 9181 2273 9239 2307
rect 9273 2273 9302 2307
rect 9696 2273 9725 2307
rect 9759 2273 9811 2307
rect 9845 2273 9903 2307
rect 9937 2273 9995 2307
rect 10029 2273 10087 2307
rect 10121 2273 10179 2307
rect 10213 2273 10271 2307
rect 10305 2273 10363 2307
rect 10397 2273 10455 2307
rect 10489 2273 10547 2307
rect 10581 2273 10639 2307
rect 10673 2273 10731 2307
rect 10765 2273 10823 2307
rect 10857 2273 10915 2307
rect 10949 2273 11007 2307
rect 11041 2273 11099 2307
rect 11133 2273 11191 2307
rect 11225 2273 11254 2307
rect 11684 2273 11713 2307
rect 11747 2273 11803 2307
rect 11837 2273 11895 2307
rect 11929 2273 11987 2307
rect 12021 2273 12079 2307
rect 12113 2273 12171 2307
rect 12205 2273 12263 2307
rect 12297 2273 12355 2307
rect 12389 2273 12447 2307
rect 12481 2273 12539 2307
rect 12573 2273 12631 2307
rect 12665 2273 12723 2307
rect 12757 2273 12815 2307
rect 12849 2273 12907 2307
rect 12941 2273 12999 2307
rect 13033 2273 13091 2307
rect 13125 2273 13183 2307
rect 13217 2273 13246 2307
rect 13638 2273 13667 2307
rect 13701 2273 13755 2307
rect 13789 2273 13847 2307
rect 13881 2273 13939 2307
rect 13973 2273 14031 2307
rect 14065 2273 14123 2307
rect 14157 2273 14215 2307
rect 14249 2273 14307 2307
rect 14341 2273 14399 2307
rect 14433 2273 14491 2307
rect 14525 2273 14583 2307
rect 14617 2273 14675 2307
rect 14709 2273 14767 2307
rect 14801 2273 14859 2307
rect 14893 2273 14951 2307
rect 14985 2273 15043 2307
rect 15077 2273 15135 2307
rect 15169 2273 15198 2307
rect 15700 2273 15729 2307
rect 15763 2273 15819 2307
rect 15853 2273 15911 2307
rect 15945 2273 16003 2307
rect 16037 2273 16095 2307
rect 16129 2273 16187 2307
rect 16221 2273 16279 2307
rect 16313 2273 16371 2307
rect 16405 2273 16463 2307
rect 16497 2273 16555 2307
rect 16589 2273 16647 2307
rect 16681 2273 16739 2307
rect 16773 2273 16831 2307
rect 16865 2273 16923 2307
rect 16957 2273 17015 2307
rect 17049 2273 17107 2307
rect 17141 2273 17199 2307
rect 17233 2273 17262 2307
rect 3109 2195 3125 2229
rect 3159 2195 3175 2229
rect 2936 2161 3056 2182
rect 3209 2193 3261 2237
rect 2936 2135 3175 2161
rect 2936 2101 2938 2135
rect 2972 2127 3175 2135
rect 2972 2101 2984 2127
rect 2186 2097 2285 2101
rect 1964 2039 1979 2073
rect 1930 2023 1979 2039
rect 2013 2067 2029 2081
rect 2013 2033 2014 2067
rect 2063 2047 2101 2081
rect 2186 2063 2269 2097
rect 2303 2063 2319 2097
rect 2353 2063 2369 2097
rect 2403 2067 2428 2097
rect 2048 2033 2101 2047
rect 2353 2033 2382 2063
rect 2416 2033 2428 2067
rect 2487 2038 2720 2095
rect 3141 2089 3175 2127
rect 3243 2159 3261 2193
rect 3209 2122 3261 2159
rect 3803 2173 3861 2267
rect 3803 2139 3815 2173
rect 3849 2139 3861 2173
rect 3803 2122 3861 2139
rect 3900 2189 3980 2233
rect 4029 2229 4095 2267
rect 4029 2195 4045 2229
rect 4079 2195 4095 2229
rect 4129 2217 4331 2233
rect 3900 2155 3946 2189
rect 4129 2183 4297 2217
rect 4129 2161 4163 2183
rect 4297 2165 4331 2183
rect 4398 2212 4432 2233
rect 4466 2229 4532 2267
rect 4466 2195 4482 2229
rect 4516 2195 4532 2229
rect 4566 2212 4600 2233
rect 3900 2122 3980 2155
rect 4015 2127 4163 2161
rect 4398 2161 4432 2178
rect 4634 2220 4700 2267
rect 4634 2186 4650 2220
rect 4684 2186 4700 2220
rect 4754 2212 4788 2233
rect 4566 2161 4600 2178
rect 1830 1953 1910 1991
rect 1830 1919 1876 1953
rect 1830 1863 1910 1919
rect 1945 1901 1979 2023
rect 2067 1969 2106 1999
rect 2067 1935 2101 1969
rect 2140 1965 2151 1999
rect 2487 1985 2521 2038
rect 2135 1935 2151 1965
rect 2197 1969 2454 1985
rect 2231 1951 2454 1969
rect 2488 1951 2521 1985
rect 2566 1999 2638 2001
rect 2600 1985 2638 1999
rect 2566 1951 2571 1965
rect 2605 1951 2638 1985
rect 2231 1935 2247 1951
rect 2566 1935 2638 1951
rect 2686 1969 2720 2038
rect 2754 2067 2832 2082
rect 3030 2073 3096 2089
rect 3030 2067 3062 2073
rect 2788 2066 2832 2067
rect 2788 2033 2798 2066
rect 2754 2032 2798 2033
rect 2754 2016 2832 2032
rect 2870 2033 2894 2067
rect 2928 2033 2944 2067
rect 3064 2033 3096 2039
rect 2870 1969 2904 2033
rect 3062 2023 3096 2033
rect 3141 2073 3192 2089
rect 3141 2039 3158 2073
rect 3141 2023 3192 2039
rect 2686 1935 2904 1969
rect 2972 1965 3018 1999
rect 2938 1962 3018 1965
rect 3141 1963 3175 2023
rect 3226 1991 3261 2122
rect 2197 1934 2247 1935
rect 1945 1867 2078 1901
rect 2197 1900 2206 1934
rect 2240 1900 2247 1934
rect 2938 1928 2984 1962
rect 2938 1912 3018 1928
rect 2197 1897 2247 1900
rect 1830 1829 1876 1863
rect 2044 1863 2078 1867
rect 2328 1867 2530 1901
rect 2044 1845 2261 1863
rect 1830 1795 1910 1829
rect 1944 1799 1960 1833
rect 1994 1799 2010 1833
rect 1944 1761 2010 1799
rect 2044 1811 2227 1845
rect 2044 1795 2261 1811
rect 2328 1850 2362 1867
rect 2496 1850 2530 1867
rect 2328 1795 2362 1816
rect 2396 1799 2412 1833
rect 2446 1799 2462 1833
rect 2396 1761 2462 1799
rect 2671 1867 2886 1901
rect 3057 1899 3175 1963
rect 3209 1950 3261 1991
rect 3243 1926 3261 1950
rect 3057 1875 3091 1899
rect 2671 1850 2718 1867
rect 2496 1795 2530 1816
rect 2564 1803 2580 1837
rect 2614 1803 2630 1837
rect 2564 1761 2630 1803
rect 2671 1816 2684 1850
rect 2852 1850 2886 1867
rect 2671 1795 2718 1816
rect 2752 1799 2768 1833
rect 2802 1799 2818 1833
rect 2752 1761 2818 1799
rect 2852 1795 2886 1816
rect 2936 1850 3091 1875
rect 3209 1890 3214 1916
rect 3254 1890 3261 1926
rect 2970 1816 3091 1850
rect 2936 1795 3091 1816
rect 3125 1841 3175 1858
rect 3159 1807 3175 1841
rect 3125 1761 3175 1807
rect 3209 1856 3261 1890
rect 3243 1822 3261 1856
rect 3209 1795 3261 1822
rect 3803 1955 3861 1990
rect 3803 1921 3815 1955
rect 3849 1921 3861 1955
rect 3803 1862 3861 1921
rect 3803 1828 3815 1862
rect 3849 1828 3861 1862
rect 1716 1727 1745 1761
rect 1779 1727 1835 1761
rect 1869 1727 1927 1761
rect 1961 1727 2019 1761
rect 2053 1727 2111 1761
rect 2145 1727 2203 1761
rect 2237 1727 2295 1761
rect 2329 1727 2387 1761
rect 2421 1727 2479 1761
rect 2513 1727 2571 1761
rect 2605 1727 2663 1761
rect 2697 1727 2755 1761
rect 2789 1727 2847 1761
rect 2881 1727 2939 1761
rect 2973 1727 3031 1761
rect 3065 1727 3123 1761
rect 3157 1727 3215 1761
rect 3249 1727 3278 1761
rect 3803 1757 3861 1828
rect 3900 1987 3966 2122
rect 4015 2085 4049 2127
rect 4000 2069 4049 2085
rect 4256 2097 4268 2131
rect 4302 2097 4355 2131
rect 4398 2127 4600 2161
rect 4822 2229 4888 2267
rect 4822 2195 4838 2229
rect 4872 2195 4888 2229
rect 4922 2212 4956 2233
rect 4754 2161 4788 2178
rect 4922 2161 4956 2178
rect 4754 2127 4956 2161
rect 5006 2212 5126 2233
rect 5040 2178 5126 2212
rect 5179 2225 5245 2267
rect 5179 2191 5195 2225
rect 5229 2191 5245 2225
rect 5006 2157 5126 2178
rect 5279 2189 5331 2233
rect 5006 2131 5245 2157
rect 5006 2097 5008 2131
rect 5042 2123 5245 2131
rect 5042 2097 5054 2123
rect 4256 2093 4355 2097
rect 4034 2035 4049 2069
rect 4000 2019 4049 2035
rect 4083 2063 4099 2077
rect 4083 2029 4084 2063
rect 4133 2043 4171 2077
rect 4256 2059 4339 2093
rect 4373 2059 4389 2093
rect 4423 2059 4439 2093
rect 4473 2063 4498 2093
rect 4118 2029 4171 2043
rect 4423 2029 4452 2059
rect 4486 2029 4498 2063
rect 4557 2034 4790 2091
rect 5211 2085 5245 2123
rect 5313 2155 5331 2189
rect 5279 2118 5331 2155
rect 5759 2173 5817 2267
rect 5759 2139 5771 2173
rect 5805 2139 5817 2173
rect 5759 2122 5817 2139
rect 5852 2189 5932 2233
rect 5981 2229 6047 2267
rect 5981 2195 5997 2229
rect 6031 2195 6047 2229
rect 6081 2217 6283 2233
rect 5852 2155 5898 2189
rect 6081 2183 6249 2217
rect 6081 2161 6115 2183
rect 6249 2165 6283 2183
rect 6350 2212 6384 2233
rect 6418 2229 6484 2267
rect 6418 2195 6434 2229
rect 6468 2195 6484 2229
rect 6518 2212 6552 2233
rect 5852 2122 5932 2155
rect 5967 2127 6115 2161
rect 6350 2161 6384 2178
rect 6586 2220 6652 2267
rect 6586 2186 6602 2220
rect 6636 2186 6652 2220
rect 6706 2212 6740 2233
rect 6518 2161 6552 2178
rect 3900 1949 3980 1987
rect 3900 1915 3946 1949
rect 3900 1859 3980 1915
rect 4015 1897 4049 2019
rect 4137 1965 4176 1995
rect 4137 1931 4171 1965
rect 4210 1961 4221 1995
rect 4557 1981 4591 2034
rect 4205 1931 4221 1961
rect 4267 1965 4524 1981
rect 4301 1947 4524 1965
rect 4558 1947 4591 1981
rect 4636 1995 4708 1997
rect 4670 1981 4708 1995
rect 4636 1947 4641 1961
rect 4675 1947 4708 1981
rect 4301 1931 4317 1947
rect 4636 1931 4708 1947
rect 4756 1965 4790 2034
rect 4824 2063 4902 2078
rect 5100 2069 5166 2085
rect 5100 2063 5132 2069
rect 4858 2062 4902 2063
rect 4858 2029 4868 2062
rect 4824 2028 4868 2029
rect 4824 2012 4902 2028
rect 4940 2029 4964 2063
rect 4998 2029 5014 2063
rect 5134 2029 5166 2035
rect 4940 1965 4974 2029
rect 5132 2019 5166 2029
rect 5211 2069 5262 2085
rect 5211 2035 5228 2069
rect 5211 2019 5262 2035
rect 4756 1931 4974 1965
rect 5042 1961 5088 1995
rect 5008 1958 5088 1961
rect 5211 1959 5245 2019
rect 5296 1987 5331 2118
rect 4267 1928 4317 1931
rect 4015 1863 4148 1897
rect 4267 1894 4274 1928
rect 4308 1894 4317 1928
rect 5008 1924 5054 1958
rect 5008 1908 5088 1924
rect 4267 1893 4317 1894
rect 3900 1825 3946 1859
rect 4114 1859 4148 1863
rect 4398 1863 4600 1897
rect 4114 1841 4331 1859
rect 3900 1791 3980 1825
rect 4014 1795 4030 1829
rect 4064 1795 4080 1829
rect 4014 1757 4080 1795
rect 4114 1807 4297 1841
rect 4114 1791 4331 1807
rect 4398 1846 4432 1863
rect 4566 1846 4600 1863
rect 4398 1791 4432 1812
rect 4466 1795 4482 1829
rect 4516 1795 4532 1829
rect 4466 1757 4532 1795
rect 4741 1863 4956 1897
rect 5127 1895 5245 1959
rect 5279 1946 5331 1987
rect 5313 1922 5331 1946
rect 5127 1871 5161 1895
rect 4741 1846 4788 1863
rect 4566 1791 4600 1812
rect 4634 1799 4650 1833
rect 4684 1799 4700 1833
rect 4634 1757 4700 1799
rect 4741 1812 4754 1846
rect 4922 1846 4956 1863
rect 4741 1791 4788 1812
rect 4822 1795 4838 1829
rect 4872 1795 4888 1829
rect 4822 1757 4888 1795
rect 4922 1791 4956 1812
rect 5006 1846 5161 1871
rect 5279 1886 5290 1912
rect 5324 1886 5331 1922
rect 5040 1812 5161 1846
rect 5006 1791 5161 1812
rect 5195 1837 5245 1854
rect 5229 1803 5245 1837
rect 5195 1757 5245 1803
rect 5279 1852 5331 1886
rect 5313 1818 5331 1852
rect 5279 1791 5331 1818
rect 5759 1955 5817 1990
rect 5759 1921 5771 1955
rect 5805 1921 5817 1955
rect 5759 1862 5817 1921
rect 5759 1828 5771 1862
rect 5805 1828 5817 1862
rect 5759 1757 5817 1828
rect 5852 1987 5918 2122
rect 5967 2085 6001 2127
rect 5952 2069 6001 2085
rect 6208 2097 6220 2131
rect 6254 2097 6307 2131
rect 6350 2127 6552 2161
rect 6774 2229 6840 2267
rect 6774 2195 6790 2229
rect 6824 2195 6840 2229
rect 6874 2212 6908 2233
rect 6706 2161 6740 2178
rect 6874 2161 6908 2178
rect 6706 2127 6908 2161
rect 6958 2212 7078 2233
rect 6992 2178 7078 2212
rect 7131 2225 7197 2267
rect 7131 2191 7147 2225
rect 7181 2191 7197 2225
rect 6958 2157 7078 2178
rect 7231 2189 7283 2233
rect 6958 2131 7197 2157
rect 6958 2097 6960 2131
rect 6994 2123 7197 2131
rect 6994 2097 7006 2123
rect 6208 2093 6307 2097
rect 5986 2035 6001 2069
rect 5952 2019 6001 2035
rect 6035 2063 6051 2077
rect 6035 2029 6036 2063
rect 6085 2043 6123 2077
rect 6208 2059 6291 2093
rect 6325 2059 6341 2093
rect 6375 2059 6391 2093
rect 6425 2063 6450 2093
rect 6070 2029 6123 2043
rect 6375 2029 6404 2059
rect 6438 2029 6450 2063
rect 6509 2034 6742 2091
rect 7163 2085 7197 2123
rect 7265 2155 7283 2189
rect 7231 2118 7283 2155
rect 7757 2179 7815 2273
rect 7757 2145 7769 2179
rect 7803 2145 7815 2179
rect 7757 2128 7815 2145
rect 7854 2195 7934 2239
rect 7983 2235 8049 2273
rect 7983 2201 7999 2235
rect 8033 2201 8049 2235
rect 8083 2223 8285 2239
rect 7854 2161 7900 2195
rect 8083 2189 8251 2223
rect 8083 2167 8117 2189
rect 8251 2171 8285 2189
rect 8352 2218 8386 2239
rect 8420 2235 8486 2273
rect 8420 2201 8436 2235
rect 8470 2201 8486 2235
rect 8520 2218 8554 2239
rect 7854 2128 7934 2161
rect 7969 2133 8117 2167
rect 8352 2167 8386 2184
rect 8588 2226 8654 2273
rect 8588 2192 8604 2226
rect 8638 2192 8654 2226
rect 8708 2218 8742 2239
rect 8520 2167 8554 2184
rect 5852 1949 5932 1987
rect 5852 1915 5898 1949
rect 5852 1859 5932 1915
rect 5967 1897 6001 2019
rect 6089 1965 6128 1995
rect 6089 1931 6123 1965
rect 6162 1961 6173 1995
rect 6509 1981 6543 2034
rect 6157 1931 6173 1961
rect 6219 1965 6476 1981
rect 6253 1947 6476 1965
rect 6510 1947 6543 1981
rect 6588 1995 6660 1997
rect 6622 1981 6660 1995
rect 6588 1947 6593 1961
rect 6627 1947 6660 1981
rect 6253 1931 6269 1947
rect 6588 1931 6660 1947
rect 6708 1965 6742 2034
rect 6776 2063 6854 2078
rect 7052 2069 7118 2085
rect 7052 2063 7084 2069
rect 6810 2062 6854 2063
rect 6810 2029 6820 2062
rect 6776 2028 6820 2029
rect 6776 2012 6854 2028
rect 6892 2029 6916 2063
rect 6950 2029 6966 2063
rect 7086 2029 7118 2035
rect 6892 1965 6926 2029
rect 7084 2019 7118 2029
rect 7163 2069 7214 2085
rect 7163 2035 7180 2069
rect 7163 2019 7214 2035
rect 6708 1931 6926 1965
rect 6994 1961 7040 1995
rect 6960 1958 7040 1961
rect 7163 1959 7197 2019
rect 7248 1987 7283 2118
rect 6219 1928 6269 1931
rect 5967 1863 6100 1897
rect 6219 1894 6226 1928
rect 6260 1894 6269 1928
rect 6960 1924 7006 1958
rect 6960 1908 7040 1924
rect 6219 1893 6269 1894
rect 5852 1825 5898 1859
rect 6066 1859 6100 1863
rect 6350 1863 6552 1897
rect 6066 1841 6283 1859
rect 5852 1791 5932 1825
rect 5966 1795 5982 1829
rect 6016 1795 6032 1829
rect 5966 1757 6032 1795
rect 6066 1807 6249 1841
rect 6066 1791 6283 1807
rect 6350 1846 6384 1863
rect 6518 1846 6552 1863
rect 6350 1791 6384 1812
rect 6418 1795 6434 1829
rect 6468 1795 6484 1829
rect 6418 1757 6484 1795
rect 6693 1863 6908 1897
rect 7079 1895 7197 1959
rect 7231 1946 7283 1987
rect 7265 1922 7283 1946
rect 7079 1871 7113 1895
rect 6693 1846 6740 1863
rect 6518 1791 6552 1812
rect 6586 1799 6602 1833
rect 6636 1799 6652 1833
rect 6586 1757 6652 1799
rect 6693 1812 6706 1846
rect 6874 1846 6908 1863
rect 6693 1791 6740 1812
rect 6774 1795 6790 1829
rect 6824 1795 6840 1829
rect 6774 1757 6840 1795
rect 6874 1791 6908 1812
rect 6958 1846 7113 1871
rect 7231 1886 7242 1912
rect 7276 1886 7283 1922
rect 6992 1812 7113 1846
rect 6958 1791 7113 1812
rect 7147 1837 7197 1854
rect 7181 1803 7197 1837
rect 7147 1757 7197 1803
rect 7231 1852 7283 1886
rect 7265 1818 7283 1852
rect 7231 1791 7283 1818
rect 7757 1961 7815 1996
rect 7757 1927 7769 1961
rect 7803 1927 7815 1961
rect 7757 1868 7815 1927
rect 7757 1834 7769 1868
rect 7803 1834 7815 1868
rect 7757 1763 7815 1834
rect 7854 1993 7920 2128
rect 7969 2091 8003 2133
rect 7954 2075 8003 2091
rect 8210 2103 8222 2137
rect 8256 2103 8309 2137
rect 8352 2133 8554 2167
rect 8776 2235 8842 2273
rect 8776 2201 8792 2235
rect 8826 2201 8842 2235
rect 8876 2218 8910 2239
rect 8708 2167 8742 2184
rect 8876 2167 8910 2184
rect 8708 2133 8910 2167
rect 8960 2218 9080 2239
rect 8994 2184 9080 2218
rect 9133 2231 9199 2273
rect 9133 2197 9149 2231
rect 9183 2197 9199 2231
rect 8960 2163 9080 2184
rect 9233 2195 9285 2239
rect 8960 2137 9199 2163
rect 8960 2103 8962 2137
rect 8996 2129 9199 2137
rect 8996 2103 9008 2129
rect 8210 2099 8309 2103
rect 7988 2041 8003 2075
rect 7954 2025 8003 2041
rect 8037 2069 8053 2083
rect 8037 2035 8038 2069
rect 8087 2049 8125 2083
rect 8210 2065 8293 2099
rect 8327 2065 8343 2099
rect 8377 2065 8393 2099
rect 8427 2069 8452 2099
rect 8072 2035 8125 2049
rect 8377 2035 8406 2065
rect 8440 2035 8452 2069
rect 8511 2040 8744 2097
rect 9165 2091 9199 2129
rect 9267 2161 9285 2195
rect 9233 2124 9285 2161
rect 9713 2179 9771 2273
rect 9713 2145 9725 2179
rect 9759 2145 9771 2179
rect 9713 2128 9771 2145
rect 9806 2195 9886 2239
rect 9935 2235 10001 2273
rect 9935 2201 9951 2235
rect 9985 2201 10001 2235
rect 10035 2223 10237 2239
rect 9806 2161 9852 2195
rect 10035 2189 10203 2223
rect 10035 2167 10069 2189
rect 10203 2171 10237 2189
rect 10304 2218 10338 2239
rect 10372 2235 10438 2273
rect 10372 2201 10388 2235
rect 10422 2201 10438 2235
rect 10472 2218 10506 2239
rect 9806 2128 9886 2161
rect 9921 2133 10069 2167
rect 10304 2167 10338 2184
rect 10540 2226 10606 2273
rect 10540 2192 10556 2226
rect 10590 2192 10606 2226
rect 10660 2218 10694 2239
rect 10472 2167 10506 2184
rect 7854 1955 7934 1993
rect 7854 1921 7900 1955
rect 7854 1865 7934 1921
rect 7969 1903 8003 2025
rect 8091 1971 8130 2001
rect 8091 1937 8125 1971
rect 8164 1967 8175 2001
rect 8511 1987 8545 2040
rect 8159 1937 8175 1967
rect 8221 1971 8478 1987
rect 8255 1953 8478 1971
rect 8512 1953 8545 1987
rect 8590 2001 8662 2003
rect 8624 1987 8662 2001
rect 8590 1953 8595 1967
rect 8629 1953 8662 1987
rect 8255 1937 8271 1953
rect 8590 1937 8662 1953
rect 8710 1971 8744 2040
rect 8778 2069 8856 2084
rect 9054 2075 9120 2091
rect 9054 2069 9086 2075
rect 8812 2068 8856 2069
rect 8812 2035 8822 2068
rect 8778 2034 8822 2035
rect 8778 2018 8856 2034
rect 8894 2035 8918 2069
rect 8952 2035 8968 2069
rect 9088 2035 9120 2041
rect 8894 1971 8928 2035
rect 9086 2025 9120 2035
rect 9165 2075 9216 2091
rect 9165 2041 9182 2075
rect 9165 2025 9216 2041
rect 8710 1937 8928 1971
rect 8996 1967 9042 2001
rect 8962 1964 9042 1967
rect 9165 1965 9199 2025
rect 9250 1993 9285 2124
rect 8221 1934 8271 1937
rect 7969 1869 8102 1903
rect 8221 1900 8228 1934
rect 8262 1900 8271 1934
rect 8962 1930 9008 1964
rect 8962 1914 9042 1930
rect 8221 1899 8271 1900
rect 7854 1831 7900 1865
rect 8068 1865 8102 1869
rect 8352 1869 8554 1903
rect 8068 1847 8285 1865
rect 7854 1797 7934 1831
rect 7968 1801 7984 1835
rect 8018 1801 8034 1835
rect 7968 1763 8034 1801
rect 8068 1813 8251 1847
rect 8068 1797 8285 1813
rect 8352 1852 8386 1869
rect 8520 1852 8554 1869
rect 8352 1797 8386 1818
rect 8420 1801 8436 1835
rect 8470 1801 8486 1835
rect 8420 1763 8486 1801
rect 8695 1869 8910 1903
rect 9081 1901 9199 1965
rect 9233 1952 9285 1993
rect 9267 1928 9285 1952
rect 9081 1877 9115 1901
rect 8695 1852 8742 1869
rect 8520 1797 8554 1818
rect 8588 1805 8604 1839
rect 8638 1805 8654 1839
rect 8588 1763 8654 1805
rect 8695 1818 8708 1852
rect 8876 1852 8910 1869
rect 8695 1797 8742 1818
rect 8776 1801 8792 1835
rect 8826 1801 8842 1835
rect 8776 1763 8842 1801
rect 8876 1797 8910 1818
rect 8960 1852 9115 1877
rect 9233 1892 9244 1918
rect 9278 1892 9285 1928
rect 8994 1818 9115 1852
rect 8960 1797 9115 1818
rect 9149 1843 9199 1860
rect 9183 1809 9199 1843
rect 9149 1763 9199 1809
rect 9233 1858 9285 1892
rect 9267 1824 9285 1858
rect 9233 1797 9285 1824
rect 9713 1961 9771 1996
rect 9713 1927 9725 1961
rect 9759 1927 9771 1961
rect 9713 1868 9771 1927
rect 9713 1834 9725 1868
rect 9759 1834 9771 1868
rect 9713 1763 9771 1834
rect 9806 1993 9872 2128
rect 9921 2091 9955 2133
rect 9906 2075 9955 2091
rect 10162 2103 10174 2137
rect 10208 2103 10261 2137
rect 10304 2133 10506 2167
rect 10728 2235 10794 2273
rect 10728 2201 10744 2235
rect 10778 2201 10794 2235
rect 10828 2218 10862 2239
rect 10660 2167 10694 2184
rect 10828 2167 10862 2184
rect 10660 2133 10862 2167
rect 10912 2218 11032 2239
rect 10946 2184 11032 2218
rect 11085 2231 11151 2273
rect 11085 2197 11101 2231
rect 11135 2197 11151 2231
rect 10912 2163 11032 2184
rect 11185 2195 11237 2239
rect 10912 2137 11151 2163
rect 10912 2103 10914 2137
rect 10948 2129 11151 2137
rect 10948 2103 10960 2129
rect 10162 2099 10261 2103
rect 9940 2041 9955 2075
rect 9906 2025 9955 2041
rect 9989 2069 10005 2083
rect 9989 2035 9990 2069
rect 10039 2049 10077 2083
rect 10162 2065 10245 2099
rect 10279 2065 10295 2099
rect 10329 2065 10345 2099
rect 10379 2069 10404 2099
rect 10024 2035 10077 2049
rect 10329 2035 10358 2065
rect 10392 2035 10404 2069
rect 10463 2040 10696 2097
rect 11117 2091 11151 2129
rect 11219 2161 11237 2195
rect 11185 2124 11237 2161
rect 11701 2179 11759 2273
rect 11701 2145 11713 2179
rect 11747 2145 11759 2179
rect 11701 2128 11759 2145
rect 11798 2195 11878 2239
rect 11927 2235 11993 2273
rect 11927 2201 11943 2235
rect 11977 2201 11993 2235
rect 12027 2223 12229 2239
rect 11798 2161 11844 2195
rect 12027 2189 12195 2223
rect 12027 2167 12061 2189
rect 12195 2171 12229 2189
rect 12296 2218 12330 2239
rect 12364 2235 12430 2273
rect 12364 2201 12380 2235
rect 12414 2201 12430 2235
rect 12464 2218 12498 2239
rect 11798 2128 11878 2161
rect 11913 2133 12061 2167
rect 12296 2167 12330 2184
rect 12532 2226 12598 2273
rect 12532 2192 12548 2226
rect 12582 2192 12598 2226
rect 12652 2218 12686 2239
rect 12464 2167 12498 2184
rect 9806 1955 9886 1993
rect 9806 1921 9852 1955
rect 9806 1865 9886 1921
rect 9921 1903 9955 2025
rect 10043 1971 10082 2001
rect 10043 1937 10077 1971
rect 10116 1967 10127 2001
rect 10463 1987 10497 2040
rect 10111 1937 10127 1967
rect 10173 1971 10430 1987
rect 10207 1953 10430 1971
rect 10464 1953 10497 1987
rect 10542 2001 10614 2003
rect 10576 1987 10614 2001
rect 10542 1953 10547 1967
rect 10581 1953 10614 1987
rect 10207 1937 10223 1953
rect 10542 1937 10614 1953
rect 10662 1971 10696 2040
rect 10730 2069 10808 2084
rect 11006 2075 11072 2091
rect 11006 2069 11038 2075
rect 10764 2068 10808 2069
rect 10764 2035 10774 2068
rect 10730 2034 10774 2035
rect 10730 2018 10808 2034
rect 10846 2035 10870 2069
rect 10904 2035 10920 2069
rect 11040 2035 11072 2041
rect 10846 1971 10880 2035
rect 11038 2025 11072 2035
rect 11117 2075 11168 2091
rect 11117 2041 11134 2075
rect 11117 2025 11168 2041
rect 10662 1937 10880 1971
rect 10948 1967 10994 2001
rect 10914 1964 10994 1967
rect 11117 1965 11151 2025
rect 11202 1993 11237 2124
rect 10173 1934 10223 1937
rect 9921 1869 10054 1903
rect 10173 1900 10180 1934
rect 10214 1900 10223 1934
rect 10914 1930 10960 1964
rect 10914 1914 10994 1930
rect 10173 1899 10223 1900
rect 9806 1831 9852 1865
rect 10020 1865 10054 1869
rect 10304 1869 10506 1903
rect 10020 1847 10237 1865
rect 9806 1797 9886 1831
rect 9920 1801 9936 1835
rect 9970 1801 9986 1835
rect 9920 1763 9986 1801
rect 10020 1813 10203 1847
rect 10020 1797 10237 1813
rect 10304 1852 10338 1869
rect 10472 1852 10506 1869
rect 10304 1797 10338 1818
rect 10372 1801 10388 1835
rect 10422 1801 10438 1835
rect 10372 1763 10438 1801
rect 10647 1869 10862 1903
rect 11033 1901 11151 1965
rect 11185 1952 11237 1993
rect 11219 1928 11237 1952
rect 11033 1877 11067 1901
rect 10647 1852 10694 1869
rect 10472 1797 10506 1818
rect 10540 1805 10556 1839
rect 10590 1805 10606 1839
rect 10540 1763 10606 1805
rect 10647 1818 10660 1852
rect 10828 1852 10862 1869
rect 10647 1797 10694 1818
rect 10728 1801 10744 1835
rect 10778 1801 10794 1835
rect 10728 1763 10794 1801
rect 10828 1797 10862 1818
rect 10912 1852 11067 1877
rect 11185 1892 11196 1918
rect 11230 1892 11237 1928
rect 10946 1818 11067 1852
rect 10912 1797 11067 1818
rect 11101 1843 11151 1860
rect 11135 1809 11151 1843
rect 11101 1763 11151 1809
rect 11185 1858 11237 1892
rect 11219 1824 11237 1858
rect 11185 1797 11237 1824
rect 11701 1961 11759 1996
rect 11701 1927 11713 1961
rect 11747 1927 11759 1961
rect 11701 1868 11759 1927
rect 11701 1834 11713 1868
rect 11747 1834 11759 1868
rect 11701 1763 11759 1834
rect 11798 1993 11864 2128
rect 11913 2091 11947 2133
rect 11898 2075 11947 2091
rect 12154 2103 12166 2137
rect 12200 2103 12253 2137
rect 12296 2133 12498 2167
rect 12720 2235 12786 2273
rect 12720 2201 12736 2235
rect 12770 2201 12786 2235
rect 12820 2218 12854 2239
rect 12652 2167 12686 2184
rect 12820 2167 12854 2184
rect 12652 2133 12854 2167
rect 12904 2218 13024 2239
rect 12938 2184 13024 2218
rect 13077 2231 13143 2273
rect 13077 2197 13093 2231
rect 13127 2197 13143 2231
rect 12904 2163 13024 2184
rect 13177 2195 13229 2239
rect 12904 2137 13143 2163
rect 12904 2103 12906 2137
rect 12940 2129 13143 2137
rect 12940 2103 12952 2129
rect 12154 2099 12253 2103
rect 11932 2041 11947 2075
rect 11898 2025 11947 2041
rect 11981 2069 11997 2083
rect 11981 2035 11982 2069
rect 12031 2049 12069 2083
rect 12154 2065 12237 2099
rect 12271 2065 12287 2099
rect 12321 2065 12337 2099
rect 12371 2069 12396 2099
rect 12016 2035 12069 2049
rect 12321 2035 12350 2065
rect 12384 2035 12396 2069
rect 12455 2040 12688 2097
rect 13109 2091 13143 2129
rect 13211 2161 13229 2195
rect 13177 2124 13229 2161
rect 13655 2179 13713 2273
rect 13655 2145 13667 2179
rect 13701 2145 13713 2179
rect 13655 2128 13713 2145
rect 13750 2195 13830 2239
rect 13879 2235 13945 2273
rect 13879 2201 13895 2235
rect 13929 2201 13945 2235
rect 13979 2223 14181 2239
rect 13750 2161 13796 2195
rect 13979 2189 14147 2223
rect 13979 2167 14013 2189
rect 14147 2171 14181 2189
rect 14248 2218 14282 2239
rect 14316 2235 14382 2273
rect 14316 2201 14332 2235
rect 14366 2201 14382 2235
rect 14416 2218 14450 2239
rect 13750 2128 13830 2161
rect 13865 2133 14013 2167
rect 14248 2167 14282 2184
rect 14484 2226 14550 2273
rect 14484 2192 14500 2226
rect 14534 2192 14550 2226
rect 14604 2218 14638 2239
rect 14416 2167 14450 2184
rect 11798 1955 11878 1993
rect 11798 1921 11844 1955
rect 11798 1865 11878 1921
rect 11913 1903 11947 2025
rect 12035 1971 12074 2001
rect 12035 1937 12069 1971
rect 12108 1967 12119 2001
rect 12455 1987 12489 2040
rect 12103 1937 12119 1967
rect 12165 1971 12422 1987
rect 12199 1953 12422 1971
rect 12456 1953 12489 1987
rect 12534 2001 12606 2003
rect 12568 1987 12606 2001
rect 12534 1953 12539 1967
rect 12573 1953 12606 1987
rect 12199 1937 12215 1953
rect 12534 1937 12606 1953
rect 12654 1971 12688 2040
rect 12722 2069 12800 2084
rect 12998 2075 13064 2091
rect 12998 2069 13030 2075
rect 12756 2068 12800 2069
rect 12756 2035 12766 2068
rect 12722 2034 12766 2035
rect 12722 2018 12800 2034
rect 12838 2035 12862 2069
rect 12896 2035 12912 2069
rect 13032 2035 13064 2041
rect 12838 1971 12872 2035
rect 13030 2025 13064 2035
rect 13109 2075 13160 2091
rect 13109 2041 13126 2075
rect 13109 2025 13160 2041
rect 12654 1937 12872 1971
rect 12940 1967 12986 2001
rect 12906 1964 12986 1967
rect 13109 1965 13143 2025
rect 13194 1993 13229 2124
rect 12165 1934 12215 1937
rect 11913 1869 12046 1903
rect 12165 1900 12172 1934
rect 12206 1900 12215 1934
rect 12906 1930 12952 1964
rect 12906 1914 12986 1930
rect 12165 1899 12215 1900
rect 11798 1831 11844 1865
rect 12012 1865 12046 1869
rect 12296 1869 12498 1903
rect 12012 1847 12229 1865
rect 11798 1797 11878 1831
rect 11912 1801 11928 1835
rect 11962 1801 11978 1835
rect 11912 1763 11978 1801
rect 12012 1813 12195 1847
rect 12012 1797 12229 1813
rect 12296 1852 12330 1869
rect 12464 1852 12498 1869
rect 12296 1797 12330 1818
rect 12364 1801 12380 1835
rect 12414 1801 12430 1835
rect 12364 1763 12430 1801
rect 12639 1869 12854 1903
rect 13025 1901 13143 1965
rect 13177 1952 13229 1993
rect 13211 1928 13229 1952
rect 13025 1877 13059 1901
rect 12639 1852 12686 1869
rect 12464 1797 12498 1818
rect 12532 1805 12548 1839
rect 12582 1805 12598 1839
rect 12532 1763 12598 1805
rect 12639 1818 12652 1852
rect 12820 1852 12854 1869
rect 12639 1797 12686 1818
rect 12720 1801 12736 1835
rect 12770 1801 12786 1835
rect 12720 1763 12786 1801
rect 12820 1797 12854 1818
rect 12904 1852 13059 1877
rect 13177 1892 13188 1918
rect 13222 1892 13229 1928
rect 12938 1818 13059 1852
rect 12904 1797 13059 1818
rect 13093 1843 13143 1860
rect 13127 1809 13143 1843
rect 13093 1763 13143 1809
rect 13177 1858 13229 1892
rect 13211 1824 13229 1858
rect 13177 1797 13229 1824
rect 13655 1961 13713 1996
rect 13655 1927 13667 1961
rect 13701 1927 13713 1961
rect 13655 1868 13713 1927
rect 13655 1834 13667 1868
rect 13701 1834 13713 1868
rect 13655 1763 13713 1834
rect 13750 1993 13816 2128
rect 13865 2091 13899 2133
rect 13850 2075 13899 2091
rect 14106 2103 14118 2137
rect 14152 2103 14205 2137
rect 14248 2133 14450 2167
rect 14672 2235 14738 2273
rect 14672 2201 14688 2235
rect 14722 2201 14738 2235
rect 14772 2218 14806 2239
rect 14604 2167 14638 2184
rect 14772 2167 14806 2184
rect 14604 2133 14806 2167
rect 14856 2218 14976 2239
rect 14890 2184 14976 2218
rect 15029 2231 15095 2273
rect 15029 2197 15045 2231
rect 15079 2197 15095 2231
rect 14856 2163 14976 2184
rect 15129 2195 15181 2239
rect 14856 2137 15095 2163
rect 14856 2103 14858 2137
rect 14892 2129 15095 2137
rect 14892 2103 14904 2129
rect 14106 2099 14205 2103
rect 13884 2041 13899 2075
rect 13850 2025 13899 2041
rect 13933 2069 13949 2083
rect 13933 2035 13934 2069
rect 13983 2049 14021 2083
rect 14106 2065 14189 2099
rect 14223 2065 14239 2099
rect 14273 2065 14289 2099
rect 14323 2069 14348 2099
rect 13968 2035 14021 2049
rect 14273 2035 14302 2065
rect 14336 2035 14348 2069
rect 14407 2040 14640 2097
rect 15061 2091 15095 2129
rect 15163 2161 15181 2195
rect 15129 2124 15181 2161
rect 15717 2179 15775 2273
rect 15717 2145 15729 2179
rect 15763 2145 15775 2179
rect 15717 2128 15775 2145
rect 15814 2195 15894 2239
rect 15943 2235 16009 2273
rect 15943 2201 15959 2235
rect 15993 2201 16009 2235
rect 16043 2223 16245 2239
rect 15814 2161 15860 2195
rect 16043 2189 16211 2223
rect 16043 2167 16077 2189
rect 16211 2171 16245 2189
rect 16312 2218 16346 2239
rect 16380 2235 16446 2273
rect 16380 2201 16396 2235
rect 16430 2201 16446 2235
rect 16480 2218 16514 2239
rect 15814 2128 15894 2161
rect 15929 2133 16077 2167
rect 16312 2167 16346 2184
rect 16548 2226 16614 2273
rect 16548 2192 16564 2226
rect 16598 2192 16614 2226
rect 16668 2218 16702 2239
rect 16480 2167 16514 2184
rect 13750 1955 13830 1993
rect 13750 1921 13796 1955
rect 13750 1865 13830 1921
rect 13865 1903 13899 2025
rect 13987 1971 14026 2001
rect 13987 1937 14021 1971
rect 14060 1967 14071 2001
rect 14407 1987 14441 2040
rect 14055 1937 14071 1967
rect 14117 1971 14374 1987
rect 14151 1953 14374 1971
rect 14408 1953 14441 1987
rect 14486 2001 14558 2003
rect 14520 1987 14558 2001
rect 14486 1953 14491 1967
rect 14525 1953 14558 1987
rect 14151 1937 14167 1953
rect 14486 1937 14558 1953
rect 14606 1971 14640 2040
rect 14674 2069 14752 2084
rect 14950 2075 15016 2091
rect 14950 2069 14982 2075
rect 14708 2068 14752 2069
rect 14708 2035 14718 2068
rect 14674 2034 14718 2035
rect 14674 2018 14752 2034
rect 14790 2035 14814 2069
rect 14848 2035 14864 2069
rect 14984 2035 15016 2041
rect 14790 1971 14824 2035
rect 14982 2025 15016 2035
rect 15061 2075 15112 2091
rect 15061 2041 15078 2075
rect 15061 2025 15112 2041
rect 14606 1937 14824 1971
rect 14892 1967 14938 2001
rect 14858 1964 14938 1967
rect 15061 1965 15095 2025
rect 15146 1993 15181 2124
rect 14117 1934 14167 1937
rect 13865 1869 13998 1903
rect 14117 1900 14124 1934
rect 14158 1900 14167 1934
rect 14858 1930 14904 1964
rect 14858 1914 14938 1930
rect 14117 1899 14167 1900
rect 13750 1831 13796 1865
rect 13964 1865 13998 1869
rect 14248 1869 14450 1903
rect 13964 1847 14181 1865
rect 13750 1797 13830 1831
rect 13864 1801 13880 1835
rect 13914 1801 13930 1835
rect 13864 1763 13930 1801
rect 13964 1813 14147 1847
rect 13964 1797 14181 1813
rect 14248 1852 14282 1869
rect 14416 1852 14450 1869
rect 14248 1797 14282 1818
rect 14316 1801 14332 1835
rect 14366 1801 14382 1835
rect 14316 1763 14382 1801
rect 14591 1869 14806 1903
rect 14977 1901 15095 1965
rect 15129 1952 15181 1993
rect 15163 1928 15181 1952
rect 14977 1877 15011 1901
rect 14591 1852 14638 1869
rect 14416 1797 14450 1818
rect 14484 1805 14500 1839
rect 14534 1805 14550 1839
rect 14484 1763 14550 1805
rect 14591 1818 14604 1852
rect 14772 1852 14806 1869
rect 14591 1797 14638 1818
rect 14672 1801 14688 1835
rect 14722 1801 14738 1835
rect 14672 1763 14738 1801
rect 14772 1797 14806 1818
rect 14856 1852 15011 1877
rect 15129 1892 15140 1918
rect 15174 1892 15181 1928
rect 14890 1818 15011 1852
rect 14856 1797 15011 1818
rect 15045 1843 15095 1860
rect 15079 1809 15095 1843
rect 15045 1763 15095 1809
rect 15129 1858 15181 1892
rect 15163 1824 15181 1858
rect 15129 1797 15181 1824
rect 15717 1961 15775 1996
rect 15717 1927 15729 1961
rect 15763 1927 15775 1961
rect 15717 1868 15775 1927
rect 15717 1834 15729 1868
rect 15763 1834 15775 1868
rect 15717 1763 15775 1834
rect 15814 1993 15880 2128
rect 15929 2091 15963 2133
rect 15914 2075 15963 2091
rect 16170 2103 16182 2137
rect 16216 2103 16269 2137
rect 16312 2133 16514 2167
rect 16736 2235 16802 2273
rect 16736 2201 16752 2235
rect 16786 2201 16802 2235
rect 16836 2218 16870 2239
rect 16668 2167 16702 2184
rect 16836 2167 16870 2184
rect 16668 2133 16870 2167
rect 16920 2218 17040 2239
rect 16954 2184 17040 2218
rect 17093 2231 17159 2273
rect 17093 2197 17109 2231
rect 17143 2197 17159 2231
rect 16920 2163 17040 2184
rect 17193 2195 17245 2239
rect 16920 2137 17159 2163
rect 16920 2103 16922 2137
rect 16956 2129 17159 2137
rect 16956 2103 16968 2129
rect 16170 2099 16269 2103
rect 15948 2041 15963 2075
rect 15914 2025 15963 2041
rect 15997 2069 16013 2083
rect 15997 2035 15998 2069
rect 16047 2049 16085 2083
rect 16170 2065 16253 2099
rect 16287 2065 16303 2099
rect 16337 2065 16353 2099
rect 16387 2069 16412 2099
rect 16032 2035 16085 2049
rect 16337 2035 16366 2065
rect 16400 2035 16412 2069
rect 16471 2040 16704 2097
rect 17125 2091 17159 2129
rect 17227 2161 17245 2195
rect 17193 2124 17245 2161
rect 15814 1955 15894 1993
rect 15814 1921 15860 1955
rect 15814 1865 15894 1921
rect 15929 1903 15963 2025
rect 16051 1971 16090 2001
rect 16051 1937 16085 1971
rect 16124 1967 16135 2001
rect 16471 1987 16505 2040
rect 16119 1937 16135 1967
rect 16181 1971 16438 1987
rect 16215 1953 16438 1971
rect 16472 1953 16505 1987
rect 16550 2001 16622 2003
rect 16584 1987 16622 2001
rect 16550 1953 16555 1967
rect 16589 1953 16622 1987
rect 16215 1937 16231 1953
rect 16550 1937 16622 1953
rect 16670 1971 16704 2040
rect 16738 2069 16816 2084
rect 17014 2075 17080 2091
rect 17014 2069 17046 2075
rect 16772 2068 16816 2069
rect 16772 2035 16782 2068
rect 16738 2034 16782 2035
rect 16738 2018 16816 2034
rect 16854 2035 16878 2069
rect 16912 2035 16928 2069
rect 17048 2035 17080 2041
rect 16854 1971 16888 2035
rect 17046 2025 17080 2035
rect 17125 2075 17176 2091
rect 17125 2041 17142 2075
rect 17125 2025 17176 2041
rect 16670 1937 16888 1971
rect 16956 1967 17002 2001
rect 16922 1964 17002 1967
rect 17125 1965 17159 2025
rect 17210 1993 17245 2124
rect 16181 1934 16231 1937
rect 15929 1869 16062 1903
rect 16181 1900 16188 1934
rect 16222 1900 16231 1934
rect 16922 1930 16968 1964
rect 16922 1914 17002 1930
rect 16181 1899 16231 1900
rect 15814 1831 15860 1865
rect 16028 1865 16062 1869
rect 16312 1869 16514 1903
rect 16028 1847 16245 1865
rect 15814 1797 15894 1831
rect 15928 1801 15944 1835
rect 15978 1801 15994 1835
rect 15928 1763 15994 1801
rect 16028 1813 16211 1847
rect 16028 1797 16245 1813
rect 16312 1852 16346 1869
rect 16480 1852 16514 1869
rect 16312 1797 16346 1818
rect 16380 1801 16396 1835
rect 16430 1801 16446 1835
rect 16380 1763 16446 1801
rect 16655 1869 16870 1903
rect 17041 1901 17159 1965
rect 17193 1952 17245 1993
rect 17227 1928 17245 1952
rect 17041 1877 17075 1901
rect 16655 1852 16702 1869
rect 16480 1797 16514 1818
rect 16548 1805 16564 1839
rect 16598 1805 16614 1839
rect 16548 1763 16614 1805
rect 16655 1818 16668 1852
rect 16836 1852 16870 1869
rect 16655 1797 16702 1818
rect 16736 1801 16752 1835
rect 16786 1801 16802 1835
rect 16736 1763 16802 1801
rect 16836 1797 16870 1818
rect 16920 1852 17075 1877
rect 17193 1892 17204 1918
rect 17238 1892 17245 1928
rect 16954 1818 17075 1852
rect 16920 1797 17075 1818
rect 17109 1843 17159 1860
rect 17143 1809 17159 1843
rect 17109 1763 17159 1809
rect 17193 1858 17245 1892
rect 17227 1824 17245 1858
rect 17193 1797 17245 1824
rect 3786 1723 3815 1757
rect 3849 1723 3905 1757
rect 3939 1723 3997 1757
rect 4031 1723 4089 1757
rect 4123 1723 4181 1757
rect 4215 1723 4273 1757
rect 4307 1723 4365 1757
rect 4399 1723 4457 1757
rect 4491 1723 4549 1757
rect 4583 1723 4641 1757
rect 4675 1723 4733 1757
rect 4767 1723 4825 1757
rect 4859 1723 4917 1757
rect 4951 1723 5009 1757
rect 5043 1723 5101 1757
rect 5135 1723 5193 1757
rect 5227 1723 5285 1757
rect 5319 1723 5348 1757
rect 5742 1723 5771 1757
rect 5805 1723 5857 1757
rect 5891 1723 5949 1757
rect 5983 1723 6041 1757
rect 6075 1723 6133 1757
rect 6167 1723 6225 1757
rect 6259 1723 6317 1757
rect 6351 1723 6409 1757
rect 6443 1723 6501 1757
rect 6535 1723 6593 1757
rect 6627 1723 6685 1757
rect 6719 1723 6777 1757
rect 6811 1723 6869 1757
rect 6903 1723 6961 1757
rect 6995 1723 7053 1757
rect 7087 1723 7145 1757
rect 7179 1723 7237 1757
rect 7271 1723 7300 1757
rect 7740 1729 7769 1763
rect 7803 1729 7859 1763
rect 7893 1729 7951 1763
rect 7985 1729 8043 1763
rect 8077 1729 8135 1763
rect 8169 1729 8227 1763
rect 8261 1729 8319 1763
rect 8353 1729 8411 1763
rect 8445 1729 8503 1763
rect 8537 1729 8595 1763
rect 8629 1729 8687 1763
rect 8721 1729 8779 1763
rect 8813 1729 8871 1763
rect 8905 1729 8963 1763
rect 8997 1729 9055 1763
rect 9089 1729 9147 1763
rect 9181 1729 9239 1763
rect 9273 1729 9302 1763
rect 9696 1729 9725 1763
rect 9759 1729 9811 1763
rect 9845 1729 9903 1763
rect 9937 1729 9995 1763
rect 10029 1729 10087 1763
rect 10121 1729 10179 1763
rect 10213 1729 10271 1763
rect 10305 1729 10363 1763
rect 10397 1729 10455 1763
rect 10489 1729 10547 1763
rect 10581 1729 10639 1763
rect 10673 1729 10731 1763
rect 10765 1729 10823 1763
rect 10857 1729 10915 1763
rect 10949 1729 11007 1763
rect 11041 1729 11099 1763
rect 11133 1729 11191 1763
rect 11225 1729 11254 1763
rect 11684 1729 11713 1763
rect 11747 1729 11803 1763
rect 11837 1729 11895 1763
rect 11929 1729 11987 1763
rect 12021 1729 12079 1763
rect 12113 1729 12171 1763
rect 12205 1729 12263 1763
rect 12297 1729 12355 1763
rect 12389 1729 12447 1763
rect 12481 1729 12539 1763
rect 12573 1729 12631 1763
rect 12665 1729 12723 1763
rect 12757 1729 12815 1763
rect 12849 1729 12907 1763
rect 12941 1729 12999 1763
rect 13033 1729 13091 1763
rect 13125 1729 13183 1763
rect 13217 1729 13246 1763
rect 13638 1729 13667 1763
rect 13701 1729 13755 1763
rect 13789 1729 13847 1763
rect 13881 1729 13939 1763
rect 13973 1729 14031 1763
rect 14065 1729 14123 1763
rect 14157 1729 14215 1763
rect 14249 1729 14307 1763
rect 14341 1729 14399 1763
rect 14433 1729 14491 1763
rect 14525 1729 14583 1763
rect 14617 1729 14675 1763
rect 14709 1729 14767 1763
rect 14801 1729 14859 1763
rect 14893 1729 14951 1763
rect 14985 1729 15043 1763
rect 15077 1729 15135 1763
rect 15169 1729 15198 1763
rect 15700 1729 15729 1763
rect 15763 1729 15819 1763
rect 15853 1729 15911 1763
rect 15945 1729 16003 1763
rect 16037 1729 16095 1763
rect 16129 1729 16187 1763
rect 16221 1729 16279 1763
rect 16313 1729 16371 1763
rect 16405 1729 16463 1763
rect 16497 1729 16555 1763
rect 16589 1729 16647 1763
rect 16681 1729 16739 1763
rect 16773 1729 16831 1763
rect 16865 1729 16923 1763
rect 16957 1729 17015 1763
rect 17049 1729 17107 1763
rect 17141 1729 17199 1763
rect 17233 1729 17262 1763
<< viali >>
rect 18579 43447 18613 43481
rect 19123 43447 19157 43481
rect 18579 43357 18613 43391
rect 19123 43357 19157 43391
rect 18579 43265 18613 43299
rect 18882 43258 18916 43294
rect 19123 43265 19157 43299
rect 18579 43173 18613 43207
rect 18579 43081 18613 43115
rect 18579 42989 18613 43023
rect 19123 43173 19157 43207
rect 19123 43081 19157 43115
rect 18579 42897 18613 42931
rect 18579 42805 18613 42839
rect 18579 42713 18613 42747
rect 18579 42621 18613 42655
rect 18579 42529 18613 42563
rect 18579 42437 18613 42471
rect 18579 42345 18613 42379
rect 18579 42253 18613 42287
rect 18579 42161 18613 42195
rect 18579 42069 18613 42103
rect 18579 41977 18613 42011
rect 19123 42989 19157 43023
rect 19123 42897 19157 42931
rect 19123 42805 19157 42839
rect 19123 42713 19157 42747
rect 19123 42621 19157 42655
rect 19123 42529 19157 42563
rect 19123 42437 19157 42471
rect 19123 42345 19157 42379
rect 19123 42253 19157 42287
rect 19123 42161 19157 42195
rect 19123 42069 19157 42103
rect 18886 41990 18891 42024
rect 18891 41990 18920 42024
rect 19123 41977 19157 42011
rect 18563 41461 18597 41495
rect 19107 41461 19141 41495
rect 18563 41369 18597 41403
rect 18868 41364 18902 41398
rect 18563 41277 18597 41311
rect 19107 41369 19141 41403
rect 18563 41185 18597 41219
rect 18563 41093 18597 41127
rect 18563 41001 18597 41035
rect 18563 40909 18597 40943
rect 18563 40817 18597 40851
rect 18563 40725 18597 40759
rect 18563 40633 18597 40667
rect 18563 40541 18597 40575
rect 18563 40449 18597 40483
rect 18563 40357 18597 40391
rect 18870 40434 18904 40468
rect 19107 41277 19141 41311
rect 19107 41185 19141 41219
rect 19107 41093 19141 41127
rect 19107 41001 19141 41035
rect 19107 40909 19141 40943
rect 19107 40817 19141 40851
rect 19107 40725 19141 40759
rect 19107 40633 19141 40667
rect 19107 40541 19141 40575
rect 19107 40449 19141 40483
rect 19107 40357 19141 40391
rect 18563 40265 18597 40299
rect 19107 40265 19141 40299
rect 18571 39665 18605 39699
rect 19115 39665 19149 39699
rect 18571 39573 18605 39607
rect 18862 39570 18896 39606
rect 18571 39481 18605 39515
rect 18571 39389 18605 39423
rect 18571 39297 18605 39331
rect 18571 39205 18605 39239
rect 18571 39113 18605 39147
rect 18571 39021 18605 39055
rect 18571 38929 18605 38963
rect 18876 39078 18910 39090
rect 18876 39056 18883 39078
rect 18883 39056 18910 39078
rect 19115 39573 19149 39607
rect 19115 39481 19149 39515
rect 19115 39389 19149 39423
rect 19115 39297 19149 39331
rect 19115 39205 19149 39239
rect 19115 39113 19149 39147
rect 19115 39021 19149 39055
rect 18571 38837 18605 38871
rect 19115 38929 19149 38963
rect 19115 38837 19149 38871
rect 18585 38403 18619 38437
rect 19129 38403 19163 38437
rect 18585 38311 18619 38345
rect 18886 38306 18920 38340
rect 19129 38311 19163 38345
rect 18585 38219 18619 38253
rect 18585 38127 18619 38161
rect 18585 38035 18619 38069
rect 18585 37943 18619 37977
rect 18585 37851 18619 37885
rect 18585 37759 18619 37793
rect 19129 38219 19163 38253
rect 19129 38127 19163 38161
rect 19129 38035 19163 38069
rect 19129 37943 19163 37977
rect 19129 37851 19163 37885
rect 18888 37767 18897 37794
rect 18897 37767 18922 37794
rect 18888 37760 18922 37767
rect 19129 37759 19163 37793
rect 18597 37249 18631 37283
rect 19141 37249 19175 37283
rect 18597 37161 18631 37195
rect 18892 37158 18926 37192
rect 19141 37161 19175 37195
rect 18597 37069 18631 37103
rect 18597 36977 18631 37011
rect 18597 36885 18631 36919
rect 18900 36893 18909 36920
rect 18909 36893 18934 36920
rect 18900 36884 18934 36893
rect 18597 36793 18631 36827
rect 19141 37069 19175 37103
rect 19141 36977 19175 37011
rect 19141 36885 19175 36919
rect 19141 36793 19175 36827
rect 18605 36365 18639 36399
rect 19149 36365 19183 36399
rect 18605 36273 18639 36307
rect 19149 36273 19183 36307
rect 18605 36181 18639 36215
rect 18904 36190 18940 36226
rect 19149 36181 19183 36215
rect 18605 36089 18639 36123
rect 18904 36097 18917 36130
rect 18917 36097 18948 36130
rect 18904 36094 18948 36097
rect 19149 36089 19183 36123
rect 18629 34977 18663 35011
rect 19173 34977 19207 35011
rect 18629 34885 18663 34919
rect 18836 34913 18870 34914
rect 18836 34880 18847 34913
rect 18847 34880 18870 34913
rect 19173 34885 19207 34919
rect 18629 34793 18663 34827
rect 19173 34793 19207 34827
rect 18629 34701 18663 34735
rect 19173 34701 19207 34735
rect 18629 34609 18663 34643
rect 19058 34630 19092 34634
rect 19058 34600 19060 34630
rect 19060 34600 19092 34630
rect 18629 34517 18663 34551
rect 19173 34609 19207 34643
rect 19173 34517 19207 34551
rect 18629 34425 18663 34459
rect 19173 34425 19207 34459
rect 18629 34333 18663 34367
rect 18629 34241 18663 34275
rect 19173 34333 19207 34367
rect 18629 34149 18663 34183
rect 18629 34057 18663 34091
rect 18867 34147 18901 34181
rect 19173 34241 19207 34275
rect 19173 34149 19207 34183
rect 18799 34060 18833 34094
rect 18629 33965 18663 33999
rect 19173 34057 19207 34091
rect 18629 33873 18663 33907
rect 19173 33965 19207 33999
rect 18629 33781 18663 33815
rect 18629 33689 18663 33723
rect 19173 33873 19207 33907
rect 18799 33748 18825 33780
rect 18825 33748 18833 33780
rect 18799 33746 18833 33748
rect 18867 33643 18901 33677
rect 19173 33781 19207 33815
rect 19173 33689 19207 33723
rect 18629 33597 18663 33631
rect 19173 33597 19207 33631
rect 18629 33505 18663 33539
rect 18988 33484 19028 33524
rect 19173 33505 19207 33539
rect 18629 33413 18663 33447
rect 18867 33405 18901 33439
rect 19173 33413 19207 33447
rect 18629 33321 18663 33355
rect 18799 33326 18833 33360
rect 18629 33229 18663 33263
rect 18940 33232 18941 33266
rect 18941 33232 18975 33266
rect 18975 33232 18976 33266
rect 19173 33321 19207 33355
rect 19173 33229 19207 33263
rect 18629 32695 18663 32729
rect 19173 32695 19207 32729
rect 18629 32603 18663 32637
rect 18836 32631 18870 32632
rect 18836 32598 18847 32631
rect 18847 32598 18870 32631
rect 19173 32603 19207 32637
rect 18629 32511 18663 32545
rect 19173 32511 19207 32545
rect 18629 32419 18663 32453
rect 19173 32419 19207 32453
rect 18629 32327 18663 32361
rect 19058 32348 19092 32352
rect 19058 32318 19060 32348
rect 19060 32318 19092 32348
rect 18629 32235 18663 32269
rect 19173 32327 19207 32361
rect 19173 32235 19207 32269
rect 18629 32143 18663 32177
rect 19173 32143 19207 32177
rect 18629 32051 18663 32085
rect 18629 31959 18663 31993
rect 19173 32051 19207 32085
rect 18629 31867 18663 31901
rect 18629 31775 18663 31809
rect 18867 31865 18901 31899
rect 19173 31959 19207 31993
rect 19173 31867 19207 31901
rect 18799 31778 18833 31812
rect 18629 31683 18663 31717
rect 19173 31775 19207 31809
rect 18629 31591 18663 31625
rect 19173 31683 19207 31717
rect 18629 31499 18663 31533
rect 18629 31407 18663 31441
rect 19173 31591 19207 31625
rect 18799 31466 18825 31498
rect 18825 31466 18833 31498
rect 18799 31464 18833 31466
rect 18867 31361 18901 31395
rect 19173 31499 19207 31533
rect 19173 31407 19207 31441
rect 18629 31315 18663 31349
rect 19173 31315 19207 31349
rect 18629 31223 18663 31257
rect 18988 31202 19028 31242
rect 19173 31223 19207 31257
rect 18629 31131 18663 31165
rect 18867 31123 18901 31157
rect 19173 31131 19207 31165
rect 18629 31039 18663 31073
rect 18799 31044 18833 31078
rect 18629 30947 18663 30981
rect 18940 30950 18941 30984
rect 18941 30950 18975 30984
rect 18975 30950 18976 30984
rect 19173 31039 19207 31073
rect 19173 30947 19207 30981
rect 18633 30449 18667 30483
rect 19177 30449 19211 30483
rect 18633 30357 18667 30391
rect 18840 30385 18874 30386
rect 18840 30352 18851 30385
rect 18851 30352 18874 30385
rect 19177 30357 19211 30391
rect 18633 30265 18667 30299
rect 19177 30265 19211 30299
rect 18633 30173 18667 30207
rect 19177 30173 19211 30207
rect 18633 30081 18667 30115
rect 19062 30102 19096 30106
rect 19062 30072 19064 30102
rect 19064 30072 19096 30102
rect 18633 29989 18667 30023
rect 19177 30081 19211 30115
rect 19177 29989 19211 30023
rect 18633 29897 18667 29931
rect 19177 29897 19211 29931
rect 18633 29805 18667 29839
rect 18633 29713 18667 29747
rect 19177 29805 19211 29839
rect 18633 29621 18667 29655
rect 18633 29529 18667 29563
rect 18871 29619 18905 29653
rect 19177 29713 19211 29747
rect 19177 29621 19211 29655
rect 18803 29532 18837 29566
rect 18633 29437 18667 29471
rect 19177 29529 19211 29563
rect 18633 29345 18667 29379
rect 19177 29437 19211 29471
rect 18633 29253 18667 29287
rect 18633 29161 18667 29195
rect 19177 29345 19211 29379
rect 18803 29220 18829 29252
rect 18829 29220 18837 29252
rect 18803 29218 18837 29220
rect 18871 29115 18905 29149
rect 19177 29253 19211 29287
rect 19177 29161 19211 29195
rect 18633 29069 18667 29103
rect 19177 29069 19211 29103
rect 18633 28977 18667 29011
rect 18992 28956 19032 28996
rect 19177 28977 19211 29011
rect 18633 28885 18667 28919
rect 18871 28877 18905 28911
rect 19177 28885 19211 28919
rect 18633 28793 18667 28827
rect 18803 28798 18837 28832
rect 18633 28701 18667 28735
rect 18944 28704 18945 28738
rect 18945 28704 18979 28738
rect 18979 28704 18980 28738
rect 19177 28793 19211 28827
rect 19177 28701 19211 28735
rect 18625 28263 18659 28297
rect 19169 28263 19203 28297
rect 18625 28171 18659 28205
rect 18832 28199 18866 28200
rect 18832 28166 18843 28199
rect 18843 28166 18866 28199
rect 19169 28171 19203 28205
rect 18625 28079 18659 28113
rect 19169 28079 19203 28113
rect 18625 27987 18659 28021
rect 19169 27987 19203 28021
rect 18625 27895 18659 27929
rect 19054 27916 19088 27920
rect 19054 27886 19056 27916
rect 19056 27886 19088 27916
rect 18625 27803 18659 27837
rect 19169 27895 19203 27929
rect 19169 27803 19203 27837
rect 18625 27711 18659 27745
rect 19169 27711 19203 27745
rect 18625 27619 18659 27653
rect 18625 27527 18659 27561
rect 19169 27619 19203 27653
rect 18625 27435 18659 27469
rect 18625 27343 18659 27377
rect 18863 27433 18897 27467
rect 19169 27527 19203 27561
rect 19169 27435 19203 27469
rect 18795 27346 18829 27380
rect 18625 27251 18659 27285
rect 19169 27343 19203 27377
rect 18625 27159 18659 27193
rect 19169 27251 19203 27285
rect 18625 27067 18659 27101
rect 18625 26975 18659 27009
rect 19169 27159 19203 27193
rect 18795 27034 18821 27066
rect 18821 27034 18829 27066
rect 18795 27032 18829 27034
rect 18863 26929 18897 26963
rect 19169 27067 19203 27101
rect 19169 26975 19203 27009
rect 18625 26883 18659 26917
rect 19169 26883 19203 26917
rect 18625 26791 18659 26825
rect 18984 26770 19024 26810
rect 19169 26791 19203 26825
rect 18625 26699 18659 26733
rect 18863 26691 18897 26725
rect 19169 26699 19203 26733
rect 18625 26607 18659 26641
rect 18795 26612 18829 26646
rect 18625 26515 18659 26549
rect 18936 26518 18937 26552
rect 18937 26518 18971 26552
rect 18971 26518 18972 26552
rect 19169 26607 19203 26641
rect 19169 26515 19203 26549
rect 18629 26017 18663 26051
rect 19173 26017 19207 26051
rect 18629 25925 18663 25959
rect 18836 25953 18870 25954
rect 18836 25920 18847 25953
rect 18847 25920 18870 25953
rect 19173 25925 19207 25959
rect 18629 25833 18663 25867
rect 19173 25833 19207 25867
rect 18629 25741 18663 25775
rect 19173 25741 19207 25775
rect 18629 25649 18663 25683
rect 19058 25670 19092 25674
rect 19058 25640 19060 25670
rect 19060 25640 19092 25670
rect 18629 25557 18663 25591
rect 19173 25649 19207 25683
rect 19173 25557 19207 25591
rect 18629 25465 18663 25499
rect 19173 25465 19207 25499
rect 18629 25373 18663 25407
rect 18629 25281 18663 25315
rect 19173 25373 19207 25407
rect 18629 25189 18663 25223
rect 18629 25097 18663 25131
rect 18867 25187 18901 25221
rect 19173 25281 19207 25315
rect 19173 25189 19207 25223
rect 18799 25100 18833 25134
rect 18629 25005 18663 25039
rect 19173 25097 19207 25131
rect 18629 24913 18663 24947
rect 19173 25005 19207 25039
rect 18629 24821 18663 24855
rect 18629 24729 18663 24763
rect 19173 24913 19207 24947
rect 18799 24788 18825 24820
rect 18825 24788 18833 24820
rect 18799 24786 18833 24788
rect 18867 24683 18901 24717
rect 19173 24821 19207 24855
rect 19173 24729 19207 24763
rect 18629 24637 18663 24671
rect 19173 24637 19207 24671
rect 18629 24545 18663 24579
rect 18988 24524 19028 24564
rect 19173 24545 19207 24579
rect 18629 24453 18663 24487
rect 18867 24445 18901 24479
rect 19173 24453 19207 24487
rect 18629 24361 18663 24395
rect 18799 24366 18833 24400
rect 18629 24269 18663 24303
rect 18940 24272 18941 24306
rect 18941 24272 18975 24306
rect 18975 24272 18976 24306
rect 19173 24361 19207 24395
rect 19173 24269 19207 24303
rect 7699 23355 7733 23389
rect 7791 23355 7825 23389
rect 7883 23355 7917 23389
rect 7975 23355 8009 23389
rect 8067 23355 8101 23389
rect 8159 23355 8193 23389
rect 8251 23355 8285 23389
rect 8343 23355 8377 23389
rect 8435 23355 8469 23389
rect 8527 23355 8561 23389
rect 8619 23355 8653 23389
rect 8711 23355 8745 23389
rect 8803 23355 8837 23389
rect 8895 23355 8929 23389
rect 8987 23355 9021 23389
rect 9079 23355 9113 23389
rect 9171 23355 9205 23389
rect 9263 23355 9297 23389
rect 9355 23355 9389 23389
rect 9447 23355 9481 23389
rect 9945 23359 9979 23393
rect 10037 23359 10071 23393
rect 10129 23359 10163 23393
rect 10221 23359 10255 23393
rect 10313 23359 10347 23393
rect 10405 23359 10439 23393
rect 10497 23359 10531 23393
rect 10589 23359 10623 23393
rect 10681 23359 10715 23393
rect 10773 23359 10807 23393
rect 10865 23359 10899 23393
rect 10957 23359 10991 23393
rect 11049 23359 11083 23393
rect 11141 23359 11175 23393
rect 11233 23359 11267 23393
rect 11325 23359 11359 23393
rect 11417 23359 11451 23393
rect 11509 23359 11543 23393
rect 11601 23359 11635 23393
rect 11693 23359 11727 23393
rect 7796 23185 7830 23219
rect 7702 23077 7736 23078
rect 7702 23043 7736 23077
rect 7702 23042 7736 23043
rect 7875 23117 7909 23151
rect 7954 22990 7994 23030
rect 8216 23193 8250 23219
rect 8216 23185 8218 23193
rect 8218 23185 8250 23193
rect 8113 23117 8147 23151
rect 8530 23185 8564 23219
rect 8617 23117 8651 23151
rect 9350 23171 9384 23182
rect 9350 23148 9383 23171
rect 9383 23148 9384 23171
rect 9070 22958 9100 22960
rect 9100 22958 9104 22960
rect 9070 22926 9104 22958
rect 10042 23189 10076 23223
rect 9948 23081 9982 23082
rect 9948 23047 9982 23081
rect 9948 23046 9982 23047
rect 10121 23121 10155 23155
rect 10200 22994 10240 23034
rect 10462 23197 10496 23223
rect 10462 23189 10464 23197
rect 10464 23189 10496 23197
rect 10359 23121 10393 23155
rect 10776 23189 10810 23223
rect 10863 23121 10897 23155
rect 11596 23175 11630 23186
rect 11596 23152 11629 23175
rect 11629 23152 11630 23175
rect 11316 22962 11346 22964
rect 11346 22962 11350 22964
rect 11316 22930 11350 22962
rect 12131 23351 12165 23385
rect 12223 23351 12257 23385
rect 12315 23351 12349 23385
rect 12407 23351 12441 23385
rect 12499 23351 12533 23385
rect 12591 23351 12625 23385
rect 12683 23351 12717 23385
rect 12775 23351 12809 23385
rect 12867 23351 12901 23385
rect 12959 23351 12993 23385
rect 13051 23351 13085 23385
rect 13143 23351 13177 23385
rect 13235 23351 13269 23385
rect 13327 23351 13361 23385
rect 13419 23351 13453 23385
rect 13511 23351 13545 23385
rect 13603 23351 13637 23385
rect 13695 23351 13729 23385
rect 13787 23351 13821 23385
rect 13879 23351 13913 23385
rect 14377 23355 14411 23389
rect 14469 23355 14503 23389
rect 14561 23355 14595 23389
rect 14653 23355 14687 23389
rect 14745 23355 14779 23389
rect 14837 23355 14871 23389
rect 14929 23355 14963 23389
rect 15021 23355 15055 23389
rect 15113 23355 15147 23389
rect 15205 23355 15239 23389
rect 15297 23355 15331 23389
rect 15389 23355 15423 23389
rect 15481 23355 15515 23389
rect 15573 23355 15607 23389
rect 15665 23355 15699 23389
rect 15757 23355 15791 23389
rect 15849 23355 15883 23389
rect 15941 23355 15975 23389
rect 16033 23355 16067 23389
rect 16125 23355 16159 23389
rect 16659 23355 16693 23389
rect 16751 23355 16785 23389
rect 16843 23355 16877 23389
rect 16935 23355 16969 23389
rect 17027 23355 17061 23389
rect 17119 23355 17153 23389
rect 17211 23355 17245 23389
rect 17303 23355 17337 23389
rect 17395 23355 17429 23389
rect 17487 23355 17521 23389
rect 17579 23355 17613 23389
rect 17671 23355 17705 23389
rect 17763 23355 17797 23389
rect 17855 23355 17889 23389
rect 17947 23355 17981 23389
rect 18039 23355 18073 23389
rect 18131 23355 18165 23389
rect 18223 23355 18257 23389
rect 18315 23355 18349 23389
rect 18407 23355 18441 23389
rect 12228 23181 12262 23215
rect 12134 23073 12168 23074
rect 12134 23039 12168 23073
rect 12134 23038 12168 23039
rect 12307 23113 12341 23147
rect 12386 22986 12426 23026
rect 12648 23189 12682 23215
rect 12648 23181 12650 23189
rect 12650 23181 12682 23189
rect 12545 23113 12579 23147
rect 7699 22811 7733 22845
rect 7791 22811 7825 22845
rect 7883 22811 7917 22845
rect 7975 22811 8009 22845
rect 8067 22811 8101 22845
rect 8159 22811 8193 22845
rect 8251 22811 8285 22845
rect 8343 22811 8377 22845
rect 8435 22811 8469 22845
rect 8527 22811 8561 22845
rect 8619 22811 8653 22845
rect 8711 22811 8745 22845
rect 8803 22811 8837 22845
rect 8895 22811 8929 22845
rect 8987 22811 9021 22845
rect 9079 22811 9113 22845
rect 9171 22811 9205 22845
rect 9263 22811 9297 22845
rect 9355 22811 9389 22845
rect 9447 22811 9481 22845
rect 9945 22815 9979 22849
rect 10037 22815 10071 22849
rect 10129 22815 10163 22849
rect 10221 22815 10255 22849
rect 10313 22815 10347 22849
rect 10405 22815 10439 22849
rect 10497 22815 10531 22849
rect 10589 22815 10623 22849
rect 10681 22815 10715 22849
rect 10773 22815 10807 22849
rect 10865 22815 10899 22849
rect 10957 22815 10991 22849
rect 11049 22815 11083 22849
rect 11141 22815 11175 22849
rect 11233 22815 11267 22849
rect 11325 22815 11359 22849
rect 11417 22815 11451 22849
rect 11509 22815 11543 22849
rect 11601 22815 11635 22849
rect 11693 22815 11727 22849
rect 12962 23181 12996 23215
rect 13049 23113 13083 23147
rect 13782 23167 13816 23178
rect 13782 23144 13815 23167
rect 13815 23144 13816 23167
rect 13502 22954 13532 22956
rect 13532 22954 13536 22956
rect 13502 22922 13536 22954
rect 14474 23185 14508 23219
rect 14380 23077 14414 23078
rect 14380 23043 14414 23077
rect 14380 23042 14414 23043
rect 14553 23117 14587 23151
rect 14632 22990 14672 23030
rect 14894 23193 14928 23219
rect 14894 23185 14896 23193
rect 14896 23185 14928 23193
rect 14791 23117 14825 23151
rect 15208 23185 15242 23219
rect 15295 23117 15329 23151
rect 16028 23171 16062 23182
rect 16028 23148 16061 23171
rect 16061 23148 16062 23171
rect 15748 22958 15778 22960
rect 15778 22958 15782 22960
rect 15748 22926 15782 22958
rect 16756 23185 16790 23219
rect 16662 23077 16696 23078
rect 16662 23043 16696 23077
rect 16662 23042 16696 23043
rect 16835 23117 16869 23151
rect 16914 22990 16954 23030
rect 17176 23193 17210 23219
rect 17176 23185 17178 23193
rect 17178 23185 17210 23193
rect 17073 23117 17107 23151
rect 17490 23185 17524 23219
rect 17577 23117 17611 23151
rect 18310 23171 18344 23182
rect 18310 23148 18343 23171
rect 18343 23148 18344 23171
rect 18030 22958 18060 22960
rect 18060 22958 18064 22960
rect 18030 22926 18064 22958
rect 12131 22807 12165 22841
rect 12223 22807 12257 22841
rect 12315 22807 12349 22841
rect 12407 22807 12441 22841
rect 12499 22807 12533 22841
rect 12591 22807 12625 22841
rect 12683 22807 12717 22841
rect 12775 22807 12809 22841
rect 12867 22807 12901 22841
rect 12959 22807 12993 22841
rect 13051 22807 13085 22841
rect 13143 22807 13177 22841
rect 13235 22807 13269 22841
rect 13327 22807 13361 22841
rect 13419 22807 13453 22841
rect 13511 22807 13545 22841
rect 13603 22807 13637 22841
rect 13695 22807 13729 22841
rect 13787 22807 13821 22841
rect 13879 22807 13913 22841
rect 14377 22811 14411 22845
rect 14469 22811 14503 22845
rect 14561 22811 14595 22845
rect 14653 22811 14687 22845
rect 14745 22811 14779 22845
rect 14837 22811 14871 22845
rect 14929 22811 14963 22845
rect 15021 22811 15055 22845
rect 15113 22811 15147 22845
rect 15205 22811 15239 22845
rect 15297 22811 15331 22845
rect 15389 22811 15423 22845
rect 15481 22811 15515 22845
rect 15573 22811 15607 22845
rect 15665 22811 15699 22845
rect 15757 22811 15791 22845
rect 15849 22811 15883 22845
rect 15941 22811 15975 22845
rect 16033 22811 16067 22845
rect 16125 22811 16159 22845
rect 16659 22811 16693 22845
rect 16751 22811 16785 22845
rect 16843 22811 16877 22845
rect 16935 22811 16969 22845
rect 17027 22811 17061 22845
rect 17119 22811 17153 22845
rect 17211 22811 17245 22845
rect 17303 22811 17337 22845
rect 17395 22811 17429 22845
rect 17487 22811 17521 22845
rect 17579 22811 17613 22845
rect 17671 22811 17705 22845
rect 17763 22811 17797 22845
rect 17855 22811 17889 22845
rect 17947 22811 17981 22845
rect 18039 22811 18073 22845
rect 18131 22811 18165 22845
rect 18223 22811 18257 22845
rect 18315 22811 18349 22845
rect 18407 22811 18441 22845
rect 9459 17777 9493 17811
rect 9551 17777 9585 17811
rect 9643 17777 9677 17811
rect 9719 17777 9753 17811
rect 16296 17667 16330 17701
rect 16374 17667 16408 17701
rect 16466 17667 16500 17701
rect 16558 17667 16592 17701
rect 17162 17669 17196 17703
rect 17248 17669 17282 17703
rect 17340 17669 17374 17703
rect 17432 17669 17466 17703
rect 15510 17629 15544 17663
rect 15596 17629 15630 17663
rect 15688 17629 15722 17663
rect 15780 17629 15814 17663
rect 9496 17532 9532 17568
rect 9596 17545 9626 17572
rect 9626 17545 9632 17572
rect 9596 17536 9632 17545
rect 17940 17659 17974 17693
rect 18016 17659 18050 17693
rect 18108 17659 18142 17693
rect 18200 17659 18234 17693
rect 19056 17661 19090 17695
rect 19138 17661 19172 17695
rect 19230 17661 19264 17695
rect 19322 17661 19356 17695
rect 19922 17663 19956 17697
rect 20012 17663 20046 17697
rect 20104 17663 20138 17697
rect 20196 17663 20230 17697
rect 15635 17402 15669 17436
rect 16413 17434 16449 17468
rect 9459 17233 9493 17267
rect 9551 17233 9585 17267
rect 9643 17233 9677 17267
rect 9719 17233 9753 17267
rect 15725 17397 15729 17428
rect 15729 17397 15763 17428
rect 15725 17394 15763 17397
rect 16517 17435 16541 17464
rect 16541 17435 16551 17464
rect 16517 17430 16551 17435
rect 17287 17442 17321 17476
rect 17377 17437 17381 17468
rect 17381 17437 17415 17468
rect 17377 17434 17415 17437
rect 18059 17438 18097 17472
rect 20692 17653 20726 17687
rect 20780 17653 20814 17687
rect 20872 17653 20906 17687
rect 20964 17653 20998 17687
rect 16296 17123 16330 17157
rect 16374 17123 16408 17157
rect 16466 17123 16500 17157
rect 16558 17123 16592 17157
rect 17162 17125 17196 17159
rect 17248 17125 17282 17159
rect 17340 17125 17374 17159
rect 17432 17125 17466 17159
rect 18147 17427 18149 17460
rect 18149 17427 18183 17460
rect 18147 17426 18183 17427
rect 19177 17428 19213 17462
rect 19281 17429 19305 17458
rect 19305 17429 19315 17458
rect 19281 17424 19315 17429
rect 20051 17436 20085 17470
rect 21394 17651 21428 17685
rect 21486 17651 21520 17685
rect 21578 17651 21612 17685
rect 21670 17651 21704 17685
rect 22178 17653 22212 17687
rect 22268 17653 22302 17687
rect 22360 17653 22394 17687
rect 22452 17653 22486 17687
rect 20141 17431 20145 17462
rect 20145 17431 20179 17462
rect 20141 17428 20179 17431
rect 20823 17432 20861 17466
rect 15510 17085 15544 17119
rect 15596 17085 15630 17119
rect 15688 17085 15722 17119
rect 15780 17085 15814 17119
rect 17940 17115 17974 17149
rect 18016 17115 18050 17149
rect 18108 17115 18142 17149
rect 18200 17115 18234 17149
rect 19056 17117 19090 17151
rect 19138 17117 19172 17151
rect 19230 17117 19264 17151
rect 19322 17117 19356 17151
rect 19922 17119 19956 17153
rect 20012 17119 20046 17153
rect 20104 17119 20138 17153
rect 20196 17119 20230 17153
rect 20911 17421 20913 17454
rect 20913 17421 20947 17454
rect 20911 17420 20947 17421
rect 23036 17643 23070 17677
rect 23128 17643 23162 17677
rect 23220 17643 23254 17677
rect 23310 17643 23344 17677
rect 21433 17418 21469 17452
rect 21537 17419 21561 17448
rect 21561 17419 21571 17448
rect 21537 17414 21571 17419
rect 22307 17426 22341 17460
rect 20692 17109 20726 17143
rect 20780 17109 20814 17143
rect 20872 17109 20906 17143
rect 20964 17109 20998 17143
rect 22397 17421 22401 17452
rect 22401 17421 22435 17452
rect 22397 17418 22435 17421
rect 23079 17422 23117 17456
rect 23167 17411 23169 17444
rect 23169 17411 23203 17444
rect 23167 17410 23203 17411
rect 21394 17107 21428 17141
rect 21486 17107 21520 17141
rect 21578 17107 21612 17141
rect 21670 17107 21704 17141
rect 22178 17109 22212 17143
rect 22268 17109 22302 17143
rect 22360 17109 22394 17143
rect 22452 17109 22486 17143
rect 23036 17099 23070 17133
rect 23128 17099 23162 17133
rect 23220 17099 23254 17133
rect 23310 17099 23344 17133
rect 16275 16677 16309 16711
rect 16365 16677 16399 16711
rect 16457 16677 16491 16711
rect 16549 16677 16583 16711
rect 4405 16569 4439 16603
rect 4497 16569 4531 16603
rect 4589 16569 4623 16603
rect 4681 16569 4715 16603
rect 4773 16569 4807 16603
rect 4865 16569 4899 16603
rect 4957 16569 4991 16603
rect 5049 16569 5083 16603
rect 9271 16573 9305 16607
rect 9363 16573 9397 16607
rect 9455 16573 9489 16607
rect 9547 16573 9581 16607
rect 9639 16573 9673 16607
rect 9731 16573 9765 16607
rect 9823 16573 9857 16607
rect 9915 16573 9949 16607
rect 5044 16383 5078 16390
rect 5044 16352 5069 16383
rect 5069 16352 5078 16383
rect 4554 16291 4588 16292
rect 4554 16258 4587 16291
rect 4587 16258 4588 16291
rect 4674 16291 4708 16294
rect 4674 16260 4704 16291
rect 4704 16260 4708 16291
rect 17133 16667 17167 16701
rect 17225 16667 17259 16701
rect 17317 16667 17351 16701
rect 17407 16667 17441 16701
rect 17915 16669 17949 16703
rect 18007 16669 18041 16703
rect 18099 16669 18133 16703
rect 18191 16669 18225 16703
rect 9910 16387 9944 16394
rect 9910 16356 9935 16387
rect 9935 16356 9944 16387
rect 16416 16399 16452 16400
rect 16416 16366 16450 16399
rect 16450 16366 16452 16399
rect 9420 16295 9454 16296
rect 9420 16262 9453 16295
rect 9453 16262 9454 16295
rect 9540 16295 9574 16298
rect 9540 16264 9570 16295
rect 9570 16264 9574 16295
rect 16502 16354 16540 16388
rect 17184 16389 17222 16392
rect 17184 16358 17218 16389
rect 17218 16358 17222 16389
rect 18621 16667 18655 16701
rect 18713 16667 18747 16701
rect 18805 16667 18839 16701
rect 18893 16667 18927 16701
rect 17278 16350 17312 16384
rect 18048 16391 18082 16396
rect 18048 16362 18058 16391
rect 18058 16362 18082 16391
rect 18150 16358 18186 16392
rect 16275 16133 16309 16167
rect 16365 16133 16399 16167
rect 16457 16133 16491 16167
rect 16549 16133 16583 16167
rect 18672 16389 18708 16390
rect 18672 16356 18706 16389
rect 18706 16356 18708 16389
rect 19389 16657 19423 16691
rect 19481 16657 19515 16691
rect 19573 16657 19607 16691
rect 19663 16657 19697 16691
rect 20263 16659 20297 16693
rect 20355 16659 20389 16693
rect 20447 16659 20481 16693
rect 20529 16659 20563 16693
rect 21385 16661 21419 16695
rect 21477 16661 21511 16695
rect 21569 16661 21603 16695
rect 21645 16661 21679 16695
rect 18758 16344 18796 16378
rect 19440 16379 19478 16382
rect 19440 16348 19474 16379
rect 19474 16348 19478 16379
rect 17133 16123 17167 16157
rect 17225 16123 17259 16157
rect 17317 16123 17351 16157
rect 17407 16123 17441 16157
rect 17915 16125 17949 16159
rect 18007 16125 18041 16159
rect 18099 16125 18133 16159
rect 18191 16125 18225 16159
rect 19534 16340 19568 16374
rect 20304 16381 20338 16386
rect 20304 16352 20314 16381
rect 20314 16352 20338 16381
rect 20406 16348 20442 16382
rect 21436 16383 21472 16384
rect 21436 16350 21470 16383
rect 21470 16350 21472 16383
rect 22153 16651 22187 16685
rect 22245 16651 22279 16685
rect 22337 16651 22371 16685
rect 22423 16651 22457 16685
rect 23027 16653 23061 16687
rect 23119 16653 23153 16687
rect 23211 16653 23245 16687
rect 23289 16653 23323 16687
rect 18621 16123 18655 16157
rect 18713 16123 18747 16157
rect 18805 16123 18839 16157
rect 18893 16123 18927 16157
rect 21522 16338 21560 16372
rect 22204 16373 22242 16376
rect 22204 16342 22238 16373
rect 22238 16342 22242 16373
rect 22298 16334 22332 16368
rect 23068 16375 23102 16380
rect 23068 16346 23078 16375
rect 23078 16346 23102 16375
rect 23170 16342 23206 16376
rect 19389 16113 19423 16147
rect 19481 16113 19515 16147
rect 19573 16113 19607 16147
rect 19663 16113 19697 16147
rect 20263 16115 20297 16149
rect 20355 16115 20389 16149
rect 20447 16115 20481 16149
rect 20529 16115 20563 16149
rect 21385 16117 21419 16151
rect 21477 16117 21511 16151
rect 21569 16117 21603 16151
rect 21645 16117 21679 16151
rect 22153 16107 22187 16141
rect 22245 16107 22279 16141
rect 22337 16107 22371 16141
rect 22423 16107 22457 16141
rect 23027 16109 23061 16143
rect 23119 16109 23153 16143
rect 23211 16109 23245 16143
rect 23289 16109 23323 16143
rect 4405 16025 4439 16059
rect 4497 16025 4531 16059
rect 4589 16025 4623 16059
rect 4681 16025 4715 16059
rect 4773 16025 4807 16059
rect 4865 16025 4899 16059
rect 4957 16025 4991 16059
rect 5049 16025 5083 16059
rect 9271 16029 9305 16063
rect 9363 16029 9397 16063
rect 9455 16029 9489 16063
rect 9547 16029 9581 16063
rect 9639 16029 9673 16063
rect 9731 16029 9765 16063
rect 9823 16029 9857 16063
rect 9915 16029 9949 16063
rect 4505 15825 4539 15859
rect 4595 15825 4629 15859
rect 4687 15825 4721 15859
rect 4779 15825 4813 15859
rect 4871 15825 4905 15859
rect 4963 15825 4997 15859
rect 9371 15829 9405 15863
rect 9461 15829 9495 15863
rect 9553 15829 9587 15863
rect 9645 15829 9679 15863
rect 9737 15829 9771 15863
rect 9829 15829 9863 15863
rect 6637 15715 6671 15749
rect 6729 15715 6763 15749
rect 6821 15715 6855 15749
rect 6913 15715 6947 15749
rect 7005 15715 7039 15749
rect 7097 15715 7131 15749
rect 7189 15715 7223 15749
rect 7281 15715 7315 15749
rect 4588 15530 4630 15570
rect 4778 15547 4820 15560
rect 4778 15520 4781 15547
rect 4781 15520 4815 15547
rect 4815 15520 4820 15547
rect 4970 15456 5006 15490
rect 6632 15364 6668 15400
rect 4505 15281 4539 15315
rect 4595 15281 4629 15315
rect 4687 15281 4721 15315
rect 4779 15281 4813 15315
rect 4871 15281 4905 15315
rect 4963 15281 4997 15315
rect 6804 15403 6819 15434
rect 6819 15403 6838 15434
rect 6804 15398 6838 15403
rect 6902 15276 6936 15310
rect 11503 15719 11537 15753
rect 11595 15719 11629 15753
rect 11687 15719 11721 15753
rect 11779 15719 11813 15753
rect 11871 15719 11905 15753
rect 11963 15719 11997 15753
rect 12055 15719 12089 15753
rect 12147 15719 12181 15753
rect 9454 15534 9496 15574
rect 9644 15551 9686 15564
rect 9644 15524 9647 15551
rect 9647 15524 9681 15551
rect 9681 15524 9686 15551
rect 6998 15344 7032 15380
rect 7190 15398 7224 15432
rect 5779 15215 5813 15249
rect 5871 15215 5905 15249
rect 5963 15215 5997 15249
rect 6055 15215 6089 15249
rect 6147 15215 6181 15249
rect 6239 15215 6273 15249
rect 9836 15460 9872 15494
rect 11498 15368 11534 15404
rect 4415 15005 4449 15039
rect 4507 15005 4541 15039
rect 4599 15005 4633 15039
rect 4691 15005 4725 15039
rect 4783 15005 4817 15039
rect 4875 15005 4909 15039
rect 4967 15005 5001 15039
rect 5059 15005 5093 15039
rect 6144 15139 6151 15148
rect 6151 15139 6184 15148
rect 6144 15112 6184 15139
rect 5056 14921 5079 14930
rect 5079 14921 5090 14930
rect 5056 14896 5090 14921
rect 5824 14937 5858 14938
rect 5824 14904 5858 14937
rect 5964 14937 6000 14938
rect 5964 14904 5965 14937
rect 5965 14904 5999 14937
rect 5999 14904 6000 14937
rect 4564 14727 4598 14728
rect 4564 14694 4597 14727
rect 4597 14694 4598 14727
rect 4684 14727 4718 14730
rect 4684 14696 4714 14727
rect 4714 14696 4718 14727
rect 9371 15285 9405 15319
rect 9461 15285 9495 15319
rect 9553 15285 9587 15319
rect 9645 15285 9679 15319
rect 9737 15285 9771 15319
rect 9829 15285 9863 15319
rect 11670 15407 11685 15438
rect 11685 15407 11704 15438
rect 11670 15402 11704 15407
rect 11768 15280 11802 15314
rect 11864 15348 11898 15384
rect 12056 15402 12090 15436
rect 10645 15219 10679 15253
rect 10737 15219 10771 15253
rect 10829 15219 10863 15253
rect 10921 15219 10955 15253
rect 11013 15219 11047 15253
rect 11105 15219 11139 15253
rect 6637 15171 6671 15205
rect 6729 15171 6763 15205
rect 6821 15171 6855 15205
rect 6913 15171 6947 15205
rect 7005 15171 7039 15205
rect 7097 15171 7131 15205
rect 7189 15171 7223 15205
rect 7281 15171 7315 15205
rect 9281 15009 9315 15043
rect 9373 15009 9407 15043
rect 9465 15009 9499 15043
rect 9557 15009 9591 15043
rect 9649 15009 9683 15043
rect 9741 15009 9775 15043
rect 9833 15009 9867 15043
rect 9925 15009 9959 15043
rect 11010 15143 11017 15152
rect 11017 15143 11050 15152
rect 11010 15116 11050 15143
rect 9922 14925 9945 14934
rect 9945 14925 9956 14934
rect 9922 14900 9956 14925
rect 10690 14941 10724 14942
rect 10690 14908 10724 14941
rect 10830 14941 10866 14942
rect 10830 14908 10831 14941
rect 10831 14908 10865 14941
rect 10865 14908 10866 14941
rect 5779 14671 5813 14705
rect 5871 14671 5905 14705
rect 5963 14671 5997 14705
rect 6055 14671 6089 14705
rect 6147 14671 6181 14705
rect 6239 14671 6273 14705
rect 9430 14731 9464 14732
rect 9430 14698 9463 14731
rect 9463 14698 9464 14731
rect 9550 14731 9584 14734
rect 9550 14700 9580 14731
rect 9580 14700 9584 14731
rect 11503 15175 11537 15209
rect 11595 15175 11629 15209
rect 11687 15175 11721 15209
rect 11779 15175 11813 15209
rect 11871 15175 11905 15209
rect 11963 15175 11997 15209
rect 12055 15175 12089 15209
rect 12147 15175 12181 15209
rect 23513 14815 23547 14849
rect 23605 14815 23639 14849
rect 23697 14815 23731 14849
rect 23789 14815 23823 14849
rect 23881 14815 23915 14849
rect 23973 14815 24007 14849
rect 24065 14815 24099 14849
rect 24157 14815 24191 14849
rect 24249 14815 24283 14849
rect 24341 14815 24375 14849
rect 24433 14815 24467 14849
rect 24525 14815 24559 14849
rect 24617 14815 24651 14849
rect 24709 14815 24743 14849
rect 24801 14815 24835 14849
rect 24893 14815 24927 14849
rect 24985 14815 25019 14849
rect 25077 14815 25111 14849
rect 25169 14815 25203 14849
rect 25261 14815 25295 14849
rect 25353 14815 25387 14849
rect 25445 14815 25479 14849
rect 10645 14675 10679 14709
rect 10737 14675 10771 14709
rect 10829 14675 10863 14709
rect 10921 14675 10955 14709
rect 11013 14675 11047 14709
rect 11105 14675 11139 14709
rect 23530 14546 23568 14580
rect 4415 14461 4449 14495
rect 4507 14461 4541 14495
rect 4599 14461 4633 14495
rect 4691 14461 4725 14495
rect 4783 14461 4817 14495
rect 4875 14461 4909 14495
rect 4967 14461 5001 14495
rect 5059 14461 5093 14495
rect 9281 14465 9315 14499
rect 9373 14465 9407 14499
rect 9465 14465 9499 14499
rect 9557 14465 9591 14499
rect 9649 14465 9683 14499
rect 9741 14465 9775 14499
rect 9833 14465 9867 14499
rect 9925 14465 9959 14499
rect 23672 14537 23708 14562
rect 23672 14528 23679 14537
rect 23679 14528 23708 14537
rect 24150 14616 24186 14650
rect 24349 14645 24383 14679
rect 23974 14509 24008 14543
rect 23790 14441 23824 14475
rect 24342 14541 24376 14543
rect 24342 14509 24349 14541
rect 24349 14509 24376 14541
rect 24456 14549 24492 14552
rect 24456 14518 24459 14549
rect 24459 14518 24492 14549
rect 24556 14554 24592 14588
rect 24712 14537 24746 14562
rect 24712 14528 24729 14537
rect 24729 14528 24746 14537
rect 24811 14509 24845 14543
rect 24995 14645 25029 14679
rect 24894 14441 24928 14475
rect 25179 14509 25213 14543
rect 25078 14441 25112 14475
rect 25356 14560 25390 14594
rect 4515 14261 4549 14295
rect 4605 14261 4639 14295
rect 4697 14261 4731 14295
rect 4789 14261 4823 14295
rect 4881 14261 4915 14295
rect 4973 14261 5007 14295
rect 5761 14249 5795 14283
rect 5853 14249 5887 14283
rect 5945 14249 5979 14283
rect 6037 14249 6071 14283
rect 6129 14249 6163 14283
rect 6221 14249 6255 14283
rect 6313 14249 6347 14283
rect 6405 14249 6439 14283
rect 4598 13966 4640 14006
rect 4788 13983 4830 13996
rect 4788 13956 4791 13983
rect 4791 13956 4825 13983
rect 4825 13956 4830 13983
rect 7751 14233 7785 14267
rect 7843 14233 7877 14267
rect 7935 14233 7969 14267
rect 8027 14233 8061 14267
rect 8119 14233 8153 14267
rect 8211 14233 8245 14267
rect 8303 14233 8337 14267
rect 9379 14265 9413 14299
rect 9471 14265 9505 14299
rect 9563 14265 9597 14299
rect 9655 14265 9689 14299
rect 9747 14265 9781 14299
rect 9839 14265 9873 14299
rect 7896 14132 7932 14166
rect 5850 13971 5884 13976
rect 5850 13942 5855 13971
rect 5855 13942 5884 13971
rect 4978 13850 5014 13884
rect 4515 13717 4549 13751
rect 4605 13717 4639 13751
rect 4697 13717 4731 13751
rect 4789 13717 4823 13751
rect 4881 13717 4915 13751
rect 4973 13717 5007 13751
rect 6020 13846 6054 13880
rect 6118 13886 6152 13920
rect 6212 13937 6237 13970
rect 6237 13937 6248 13970
rect 6212 13932 6248 13937
rect 8212 14058 8237 14076
rect 8237 14058 8254 14076
rect 6394 13849 6399 13852
rect 6399 13849 6432 13852
rect 6823 13875 6857 13909
rect 6915 13875 6949 13909
rect 7007 13875 7041 13909
rect 7099 13875 7133 13909
rect 7191 13875 7225 13909
rect 7279 13875 7313 13909
rect 7752 13921 7757 13938
rect 7757 13921 7791 13938
rect 7791 13921 7792 13938
rect 7752 13904 7792 13921
rect 8212 14036 8254 14058
rect 7880 13955 7930 13960
rect 7880 13921 7883 13955
rect 7883 13921 7917 13955
rect 7917 13921 7930 13955
rect 7880 13918 7930 13921
rect 8052 13955 8090 13956
rect 8052 13921 8059 13955
rect 8059 13921 8090 13955
rect 8052 13920 8090 13921
rect 6394 13815 6432 13849
rect 6394 13814 6399 13815
rect 6399 13814 6432 13815
rect 5761 13705 5795 13739
rect 5853 13705 5887 13739
rect 5945 13705 5979 13739
rect 6037 13705 6071 13739
rect 6129 13705 6163 13739
rect 6221 13705 6255 13739
rect 6313 13705 6347 13739
rect 6405 13705 6439 13739
rect 7162 13731 7173 13764
rect 7173 13731 7196 13764
rect 7162 13730 7196 13731
rect 6834 13520 6868 13554
rect 7012 13597 7046 13604
rect 7012 13570 7030 13597
rect 7030 13570 7046 13597
rect 10627 14253 10661 14287
rect 10719 14253 10753 14287
rect 10811 14253 10845 14287
rect 10903 14253 10937 14287
rect 10995 14253 11029 14287
rect 11087 14253 11121 14287
rect 11179 14253 11213 14287
rect 11271 14253 11305 14287
rect 23513 14271 23547 14305
rect 23605 14271 23639 14305
rect 23697 14271 23731 14305
rect 23789 14271 23823 14305
rect 23881 14271 23915 14305
rect 23973 14271 24007 14305
rect 24065 14271 24099 14305
rect 24157 14271 24191 14305
rect 24249 14271 24283 14305
rect 24341 14271 24375 14305
rect 24433 14271 24467 14305
rect 24525 14271 24559 14305
rect 24617 14271 24651 14305
rect 24709 14271 24743 14305
rect 24801 14271 24835 14305
rect 24893 14271 24927 14305
rect 24985 14271 25019 14305
rect 25077 14271 25111 14305
rect 25169 14271 25203 14305
rect 25261 14271 25295 14305
rect 25353 14271 25387 14305
rect 25445 14271 25479 14305
rect 9464 13970 9506 14010
rect 9654 13987 9696 14000
rect 9654 13960 9657 13987
rect 9657 13960 9691 13987
rect 9691 13960 9696 13987
rect 12617 14237 12651 14271
rect 12709 14237 12743 14271
rect 12801 14237 12835 14271
rect 12893 14237 12927 14271
rect 12985 14237 13019 14271
rect 13077 14237 13111 14271
rect 13169 14237 13203 14271
rect 12762 14136 12798 14170
rect 10716 13975 10750 13980
rect 10716 13946 10721 13975
rect 10721 13946 10750 13975
rect 9844 13854 9880 13888
rect 7751 13689 7785 13723
rect 7843 13689 7877 13723
rect 7935 13689 7969 13723
rect 8027 13689 8061 13723
rect 8119 13689 8153 13723
rect 8211 13689 8245 13723
rect 8303 13689 8337 13723
rect 9379 13721 9413 13755
rect 9471 13721 9505 13755
rect 9563 13721 9597 13755
rect 9655 13721 9689 13755
rect 9747 13721 9781 13755
rect 9839 13721 9873 13755
rect 10886 13850 10920 13884
rect 10984 13890 11018 13924
rect 11078 13941 11103 13974
rect 11103 13941 11114 13974
rect 11078 13936 11114 13941
rect 13078 14062 13103 14080
rect 13103 14062 13120 14080
rect 11260 13853 11265 13856
rect 11265 13853 11298 13856
rect 11689 13879 11723 13913
rect 11781 13879 11815 13913
rect 11873 13879 11907 13913
rect 11965 13879 11999 13913
rect 12057 13879 12091 13913
rect 12147 13879 12181 13913
rect 12618 13925 12623 13942
rect 12623 13925 12657 13942
rect 12657 13925 12658 13942
rect 12618 13908 12658 13925
rect 13078 14040 13120 14062
rect 12746 13959 12796 13964
rect 12746 13925 12749 13959
rect 12749 13925 12783 13959
rect 12783 13925 12796 13959
rect 12746 13922 12796 13925
rect 12918 13959 12956 13960
rect 12918 13925 12925 13959
rect 12925 13925 12956 13959
rect 12918 13924 12956 13925
rect 11260 13819 11298 13853
rect 11260 13818 11265 13819
rect 11265 13818 11298 13819
rect 10627 13709 10661 13743
rect 10719 13709 10753 13743
rect 10811 13709 10845 13743
rect 10903 13709 10937 13743
rect 10995 13709 11029 13743
rect 11087 13709 11121 13743
rect 11179 13709 11213 13743
rect 11271 13709 11305 13743
rect 12028 13735 12039 13768
rect 12039 13735 12062 13768
rect 12028 13734 12062 13735
rect 11700 13524 11734 13558
rect 5885 13407 5919 13441
rect 5977 13407 6011 13441
rect 6069 13407 6103 13441
rect 6161 13407 6195 13441
rect 6253 13407 6287 13441
rect 6345 13407 6379 13441
rect 4407 13337 4441 13371
rect 4499 13337 4533 13371
rect 4591 13337 4625 13371
rect 4683 13337 4717 13371
rect 4775 13337 4809 13371
rect 4867 13337 4901 13371
rect 4959 13337 4993 13371
rect 5051 13337 5085 13371
rect 5048 13219 5082 13220
rect 5048 13186 5071 13219
rect 5071 13186 5082 13219
rect 6146 13322 6155 13334
rect 6155 13322 6182 13334
rect 6146 13298 6182 13322
rect 11878 13601 11912 13608
rect 11878 13574 11896 13601
rect 11896 13574 11912 13601
rect 12617 13693 12651 13727
rect 12709 13693 12743 13727
rect 12801 13693 12835 13727
rect 12893 13693 12927 13727
rect 12985 13693 13019 13727
rect 13077 13693 13111 13727
rect 13169 13693 13203 13727
rect 10751 13411 10785 13445
rect 10843 13411 10877 13445
rect 10935 13411 10969 13445
rect 11027 13411 11061 13445
rect 11119 13411 11153 13445
rect 11211 13411 11245 13445
rect 6823 13331 6857 13365
rect 6915 13331 6949 13365
rect 7007 13331 7041 13365
rect 7099 13331 7133 13365
rect 7191 13331 7225 13365
rect 7279 13331 7313 13365
rect 9273 13341 9307 13375
rect 9365 13341 9399 13375
rect 9457 13341 9491 13375
rect 9549 13341 9583 13375
rect 9641 13341 9675 13375
rect 9733 13341 9767 13375
rect 9825 13341 9859 13375
rect 9917 13341 9951 13375
rect 6342 13249 6373 13278
rect 6373 13249 6380 13278
rect 6342 13240 6380 13249
rect 4556 13059 4590 13060
rect 4556 13026 4589 13059
rect 4589 13026 4590 13059
rect 4676 13059 4710 13062
rect 4676 13028 4706 13059
rect 4706 13028 4710 13059
rect 5994 13049 6017 13060
rect 6017 13049 6028 13060
rect 5994 13026 6028 13049
rect 6196 13032 6232 13066
rect 9914 13223 9948 13224
rect 9914 13190 9937 13223
rect 9937 13190 9948 13223
rect 11012 13326 11021 13338
rect 11021 13326 11048 13338
rect 11012 13302 11048 13326
rect 11689 13335 11723 13369
rect 11781 13335 11815 13369
rect 11873 13335 11907 13369
rect 11965 13335 11999 13369
rect 12057 13335 12091 13369
rect 12147 13335 12181 13369
rect 11208 13253 11239 13282
rect 11239 13253 11246 13282
rect 11208 13244 11246 13253
rect 9422 13063 9456 13064
rect 9422 13030 9455 13063
rect 9455 13030 9456 13063
rect 9542 13063 9576 13066
rect 9542 13032 9572 13063
rect 9572 13032 9576 13063
rect 5885 12863 5919 12897
rect 5977 12863 6011 12897
rect 6069 12863 6103 12897
rect 6161 12863 6195 12897
rect 6253 12863 6287 12897
rect 6345 12863 6379 12897
rect 10860 13053 10883 13064
rect 10883 13053 10894 13064
rect 10860 13030 10894 13053
rect 11062 13036 11098 13070
rect 10751 12867 10785 12901
rect 10843 12867 10877 12901
rect 10935 12867 10969 12901
rect 11027 12867 11061 12901
rect 11119 12867 11153 12901
rect 11211 12867 11245 12901
rect 4407 12793 4441 12827
rect 4499 12793 4533 12827
rect 4591 12793 4625 12827
rect 4683 12793 4717 12827
rect 4775 12793 4809 12827
rect 4867 12793 4901 12827
rect 4959 12793 4993 12827
rect 5051 12793 5085 12827
rect 9273 12797 9307 12831
rect 9365 12797 9399 12831
rect 9457 12797 9491 12831
rect 9549 12797 9583 12831
rect 9641 12797 9675 12831
rect 9733 12797 9767 12831
rect 9825 12797 9859 12831
rect 9917 12797 9951 12831
rect 4507 12593 4541 12627
rect 4597 12593 4631 12627
rect 4689 12593 4723 12627
rect 4781 12593 4815 12627
rect 4873 12593 4907 12627
rect 4965 12593 4999 12627
rect 9371 12597 9405 12631
rect 9463 12597 9497 12631
rect 9555 12597 9589 12631
rect 9647 12597 9681 12631
rect 9739 12597 9773 12631
rect 9831 12597 9865 12631
rect 4590 12298 4632 12338
rect 5881 12387 5915 12421
rect 5973 12387 6007 12421
rect 6065 12387 6099 12421
rect 6157 12387 6191 12421
rect 6249 12387 6283 12421
rect 6341 12387 6375 12421
rect 4970 12336 5006 12370
rect 4780 12315 4822 12328
rect 4780 12288 4783 12315
rect 4783 12288 4817 12315
rect 4817 12288 4822 12315
rect 9456 12302 9498 12342
rect 10747 12391 10781 12425
rect 10839 12391 10873 12425
rect 10931 12391 10965 12425
rect 11023 12391 11057 12425
rect 11115 12391 11149 12425
rect 11207 12391 11241 12425
rect 9836 12340 9872 12374
rect 9646 12319 9688 12332
rect 9646 12292 9649 12319
rect 9649 12292 9683 12319
rect 9683 12292 9688 12319
rect 6346 12162 6380 12196
rect 4507 12049 4541 12083
rect 4597 12049 4631 12083
rect 4689 12049 4723 12083
rect 4781 12049 4815 12083
rect 4873 12049 4907 12083
rect 4965 12049 4999 12083
rect 6018 12109 6054 12112
rect 6018 12078 6052 12109
rect 6052 12078 6054 12109
rect 6158 12109 6194 12110
rect 6158 12076 6159 12109
rect 6159 12076 6193 12109
rect 6193 12076 6194 12109
rect 11212 12166 11246 12200
rect 9371 12053 9405 12087
rect 9463 12053 9497 12087
rect 9555 12053 9589 12087
rect 9647 12053 9681 12087
rect 9739 12053 9773 12087
rect 9831 12053 9865 12087
rect 10884 12113 10920 12116
rect 10884 12082 10918 12113
rect 10918 12082 10920 12113
rect 11024 12113 11060 12114
rect 11024 12080 11025 12113
rect 11025 12080 11059 12113
rect 11059 12080 11060 12113
rect 5881 11843 5915 11877
rect 5973 11843 6007 11877
rect 6065 11843 6099 11877
rect 6157 11843 6191 11877
rect 6249 11843 6283 11877
rect 6341 11843 6375 11877
rect 10747 11847 10781 11881
rect 10839 11847 10873 11881
rect 10931 11847 10965 11881
rect 11023 11847 11057 11881
rect 11115 11847 11149 11881
rect 11207 11847 11241 11881
rect 4417 11773 4451 11807
rect 4509 11773 4543 11807
rect 4601 11773 4635 11807
rect 4693 11773 4727 11807
rect 4785 11773 4819 11807
rect 4877 11773 4911 11807
rect 4969 11773 5003 11807
rect 5061 11773 5095 11807
rect 9283 11777 9317 11811
rect 9375 11777 9409 11811
rect 9467 11777 9501 11811
rect 9559 11777 9593 11811
rect 9651 11777 9685 11811
rect 9743 11777 9777 11811
rect 9835 11777 9869 11811
rect 9927 11777 9961 11811
rect 5048 11655 5084 11656
rect 5048 11622 5081 11655
rect 5081 11622 5084 11655
rect 4566 11495 4600 11496
rect 4566 11462 4599 11495
rect 4599 11462 4600 11495
rect 4686 11495 4720 11498
rect 4686 11464 4716 11495
rect 4716 11464 4720 11495
rect 9914 11659 9950 11660
rect 9914 11626 9947 11659
rect 9947 11626 9950 11659
rect 9432 11499 9466 11500
rect 9432 11466 9465 11499
rect 9465 11466 9466 11499
rect 9552 11499 9586 11502
rect 9552 11468 9582 11499
rect 9582 11468 9586 11499
rect 4417 11229 4451 11263
rect 4509 11229 4543 11263
rect 4601 11229 4635 11263
rect 4693 11229 4727 11263
rect 4785 11229 4819 11263
rect 4877 11229 4911 11263
rect 4969 11229 5003 11263
rect 5061 11229 5095 11263
rect 9283 11233 9317 11267
rect 9375 11233 9409 11267
rect 9467 11233 9501 11267
rect 9559 11233 9593 11267
rect 9651 11233 9685 11267
rect 9743 11233 9777 11267
rect 9835 11233 9869 11267
rect 9927 11233 9961 11267
rect 4515 11029 4549 11063
rect 4607 11029 4641 11063
rect 4699 11029 4733 11063
rect 4791 11029 4825 11063
rect 4883 11029 4917 11063
rect 4975 11029 5009 11063
rect 9381 11033 9415 11067
rect 9473 11033 9507 11067
rect 9565 11033 9599 11067
rect 9657 11033 9691 11067
rect 9749 11033 9783 11067
rect 9841 11033 9875 11067
rect 4600 10734 4642 10774
rect 4790 10751 4832 10764
rect 4790 10724 4793 10751
rect 4793 10724 4827 10751
rect 4827 10724 4832 10751
rect 4982 10694 5016 10730
rect 9466 10738 9508 10778
rect 9656 10755 9698 10768
rect 9656 10728 9659 10755
rect 9659 10728 9693 10755
rect 9693 10728 9698 10755
rect 9848 10698 9882 10734
rect 4515 10485 4549 10519
rect 4607 10485 4641 10519
rect 4699 10485 4733 10519
rect 4791 10485 4825 10519
rect 4883 10485 4917 10519
rect 4975 10485 5009 10519
rect 9381 10489 9415 10523
rect 9473 10489 9507 10523
rect 9565 10489 9599 10523
rect 9657 10489 9691 10523
rect 9749 10489 9783 10523
rect 9841 10489 9875 10523
rect 6141 6583 6175 6617
rect 6233 6583 6267 6617
rect 6325 6583 6359 6617
rect 6407 6583 6441 6617
rect 6178 6348 6212 6382
rect 6274 6351 6308 6384
rect 6274 6350 6308 6351
rect 6141 6039 6175 6073
rect 6233 6039 6267 6073
rect 6325 6039 6359 6073
rect 6407 6039 6441 6073
rect 9957 5951 9991 5985
rect 10047 5951 10081 5985
rect 10139 5951 10173 5985
rect 10231 5951 10265 5985
rect 10323 5951 10357 5985
rect 10415 5951 10449 5985
rect 10507 5951 10541 5985
rect 10599 5951 10633 5985
rect 10691 5951 10725 5985
rect 10783 5951 10817 5985
rect 10875 5951 10909 5985
rect 10967 5951 11001 5985
rect 11059 5951 11093 5985
rect 11151 5951 11185 5985
rect 11243 5951 11277 5985
rect 11335 5951 11369 5985
rect 11427 5951 11461 5985
rect 1775 5531 1809 5565
rect 1865 5531 1899 5565
rect 1957 5531 1991 5565
rect 2049 5531 2083 5565
rect 2141 5531 2175 5565
rect 2233 5531 2267 5565
rect 2325 5531 2359 5565
rect 2417 5531 2451 5565
rect 2509 5531 2543 5565
rect 2601 5531 2635 5565
rect 2693 5531 2727 5565
rect 2785 5531 2819 5565
rect 2877 5531 2911 5565
rect 2969 5531 3003 5565
rect 3061 5531 3095 5565
rect 3153 5531 3187 5565
rect 3245 5531 3279 5565
rect 2228 5361 2262 5395
rect 3909 5523 3943 5557
rect 3999 5523 4033 5557
rect 4091 5523 4125 5557
rect 4183 5523 4217 5557
rect 4275 5523 4309 5557
rect 4367 5523 4401 5557
rect 4459 5523 4493 5557
rect 4551 5523 4585 5557
rect 4643 5523 4677 5557
rect 4735 5523 4769 5557
rect 4827 5523 4861 5557
rect 4919 5523 4953 5557
rect 5011 5523 5045 5557
rect 5103 5523 5137 5557
rect 5195 5523 5229 5557
rect 5287 5523 5321 5557
rect 5379 5523 5413 5557
rect 5859 5523 5893 5557
rect 5951 5523 5985 5557
rect 6043 5523 6077 5557
rect 6135 5523 6169 5557
rect 6227 5523 6261 5557
rect 6319 5523 6353 5557
rect 6411 5523 6445 5557
rect 6503 5523 6537 5557
rect 6595 5523 6629 5557
rect 6687 5523 6721 5557
rect 6779 5523 6813 5557
rect 6871 5523 6905 5557
rect 6963 5523 6997 5557
rect 7055 5523 7089 5557
rect 7147 5523 7181 5557
rect 7239 5523 7273 5557
rect 7331 5523 7365 5557
rect 7861 5529 7895 5563
rect 7953 5529 7987 5563
rect 8045 5529 8079 5563
rect 8137 5529 8171 5563
rect 8229 5529 8263 5563
rect 8321 5529 8355 5563
rect 8413 5529 8447 5563
rect 8505 5529 8539 5563
rect 8597 5529 8631 5563
rect 8689 5529 8723 5563
rect 8781 5529 8815 5563
rect 8873 5529 8907 5563
rect 8965 5529 8999 5563
rect 9057 5529 9091 5563
rect 9149 5529 9183 5563
rect 9241 5529 9275 5563
rect 9333 5529 9367 5563
rect 2968 5361 3002 5395
rect 2044 5307 2059 5327
rect 2059 5307 2078 5327
rect 2412 5323 2433 5327
rect 2433 5323 2446 5327
rect 2044 5293 2078 5307
rect 2412 5293 2446 5323
rect 2136 5229 2170 5259
rect 2136 5225 2165 5229
rect 2165 5225 2170 5229
rect 2596 5245 2630 5259
rect 2596 5225 2601 5245
rect 2601 5225 2630 5245
rect 2784 5293 2818 5327
rect 3060 5299 3092 5327
rect 3092 5299 3094 5327
rect 3060 5293 3094 5299
rect 2968 5225 3002 5259
rect 2236 5160 2270 5194
rect 3244 5176 3273 5186
rect 3273 5176 3284 5186
rect 3244 5150 3284 5176
rect 1775 4987 1809 5021
rect 1865 4987 1899 5021
rect 1957 4987 1991 5021
rect 2049 4987 2083 5021
rect 2141 4987 2175 5021
rect 2233 4987 2267 5021
rect 2325 4987 2359 5021
rect 2417 4987 2451 5021
rect 2509 4987 2543 5021
rect 2601 4987 2635 5021
rect 2693 4987 2727 5021
rect 2785 4987 2819 5021
rect 2877 4987 2911 5021
rect 2969 4987 3003 5021
rect 3061 4987 3095 5021
rect 3153 4987 3187 5021
rect 3245 4987 3279 5021
rect 4362 5353 4396 5387
rect 5102 5353 5136 5387
rect 4178 5299 4193 5319
rect 4193 5299 4212 5319
rect 4546 5315 4567 5319
rect 4567 5315 4580 5319
rect 4178 5285 4212 5299
rect 4546 5285 4580 5315
rect 4270 5221 4304 5251
rect 4270 5217 4299 5221
rect 4299 5217 4304 5221
rect 4730 5237 4764 5251
rect 4730 5217 4735 5237
rect 4735 5217 4764 5237
rect 4918 5285 4952 5319
rect 5194 5291 5226 5319
rect 5226 5291 5228 5319
rect 5194 5285 5228 5291
rect 5102 5217 5136 5251
rect 4368 5150 4402 5184
rect 5384 5168 5407 5178
rect 5407 5168 5418 5178
rect 5384 5142 5418 5168
rect 6314 5353 6348 5387
rect 7054 5353 7088 5387
rect 6130 5299 6145 5319
rect 6145 5299 6164 5319
rect 6498 5315 6519 5319
rect 6519 5315 6532 5319
rect 6130 5285 6164 5299
rect 6498 5285 6532 5315
rect 6222 5221 6256 5251
rect 6222 5217 6251 5221
rect 6251 5217 6256 5221
rect 6682 5237 6716 5251
rect 6682 5217 6687 5237
rect 6687 5217 6716 5237
rect 6870 5285 6904 5319
rect 7146 5291 7178 5319
rect 7178 5291 7180 5319
rect 7146 5285 7180 5291
rect 7054 5217 7088 5251
rect 6320 5150 6354 5184
rect 7336 5168 7359 5178
rect 7359 5168 7370 5178
rect 7336 5142 7370 5168
rect 8316 5359 8350 5393
rect 9056 5359 9090 5393
rect 8132 5305 8147 5325
rect 8147 5305 8166 5325
rect 8500 5321 8521 5325
rect 8521 5321 8534 5325
rect 8132 5291 8166 5305
rect 8500 5291 8534 5321
rect 10410 5781 10444 5815
rect 12017 5939 12051 5973
rect 12109 5939 12143 5973
rect 12201 5939 12235 5973
rect 12293 5939 12327 5973
rect 12385 5939 12419 5973
rect 12477 5939 12511 5973
rect 12569 5939 12603 5973
rect 12661 5939 12695 5973
rect 12753 5939 12787 5973
rect 12845 5939 12879 5973
rect 12937 5939 12971 5973
rect 13029 5939 13063 5973
rect 13121 5939 13155 5973
rect 13213 5939 13247 5973
rect 13305 5939 13339 5973
rect 13397 5939 13431 5973
rect 13489 5939 13523 5973
rect 13975 5947 14009 5981
rect 14067 5947 14101 5981
rect 14159 5947 14193 5981
rect 14251 5947 14285 5981
rect 14343 5947 14377 5981
rect 14435 5947 14469 5981
rect 14527 5947 14561 5981
rect 14619 5947 14653 5981
rect 14711 5947 14745 5981
rect 14803 5947 14837 5981
rect 14895 5947 14929 5981
rect 14987 5947 15021 5981
rect 15079 5947 15113 5981
rect 15171 5947 15205 5981
rect 15263 5947 15297 5981
rect 15355 5947 15389 5981
rect 15447 5947 15481 5981
rect 15971 5953 16005 5987
rect 16061 5953 16095 5987
rect 16153 5953 16187 5987
rect 16245 5953 16279 5987
rect 16337 5953 16371 5987
rect 16429 5953 16463 5987
rect 16521 5953 16555 5987
rect 16613 5953 16647 5987
rect 16705 5953 16739 5987
rect 16797 5953 16831 5987
rect 16889 5953 16923 5987
rect 16981 5953 17015 5987
rect 17073 5953 17107 5987
rect 17165 5953 17199 5987
rect 17257 5953 17291 5987
rect 17349 5953 17383 5987
rect 17441 5953 17475 5987
rect 11150 5781 11184 5815
rect 10226 5727 10241 5747
rect 10241 5727 10260 5747
rect 10594 5743 10615 5747
rect 10615 5743 10628 5747
rect 10226 5713 10260 5727
rect 10594 5713 10628 5743
rect 10318 5649 10352 5679
rect 10318 5645 10347 5649
rect 10347 5645 10352 5649
rect 10778 5665 10812 5679
rect 10778 5645 10783 5665
rect 10783 5645 10812 5665
rect 10966 5713 11000 5747
rect 11242 5719 11274 5747
rect 11274 5719 11276 5747
rect 11242 5713 11276 5719
rect 11150 5645 11184 5679
rect 10418 5580 10452 5614
rect 11426 5596 11455 5606
rect 11455 5596 11466 5606
rect 11426 5570 11466 5596
rect 9957 5407 9991 5441
rect 10047 5407 10081 5441
rect 10139 5407 10173 5441
rect 10231 5407 10265 5441
rect 10323 5407 10357 5441
rect 10415 5407 10449 5441
rect 10507 5407 10541 5441
rect 10599 5407 10633 5441
rect 10691 5407 10725 5441
rect 10783 5407 10817 5441
rect 10875 5407 10909 5441
rect 10967 5407 11001 5441
rect 11059 5407 11093 5441
rect 11151 5407 11185 5441
rect 11243 5407 11277 5441
rect 11335 5407 11369 5441
rect 11427 5407 11461 5441
rect 12472 5769 12506 5803
rect 13212 5769 13246 5803
rect 12288 5715 12303 5735
rect 12303 5715 12322 5735
rect 12656 5731 12677 5735
rect 12677 5731 12690 5735
rect 12288 5701 12322 5715
rect 12656 5701 12690 5731
rect 12380 5637 12414 5667
rect 12380 5633 12409 5637
rect 12409 5633 12414 5637
rect 12840 5653 12874 5667
rect 12840 5633 12845 5653
rect 12845 5633 12874 5653
rect 13028 5701 13062 5735
rect 13304 5707 13336 5735
rect 13336 5707 13338 5735
rect 13304 5701 13338 5707
rect 13212 5633 13246 5667
rect 12478 5566 12512 5600
rect 13494 5584 13517 5594
rect 13517 5584 13528 5594
rect 13494 5558 13528 5584
rect 14430 5777 14464 5811
rect 15170 5777 15204 5811
rect 14246 5723 14261 5743
rect 14261 5723 14280 5743
rect 14614 5739 14635 5743
rect 14635 5739 14648 5743
rect 14246 5709 14280 5723
rect 14614 5709 14648 5739
rect 14338 5645 14372 5675
rect 14338 5641 14367 5645
rect 14367 5641 14372 5645
rect 14798 5661 14832 5675
rect 14798 5641 14803 5661
rect 14803 5641 14832 5661
rect 14986 5709 15020 5743
rect 15262 5715 15294 5743
rect 15294 5715 15296 5743
rect 15262 5709 15296 5715
rect 15170 5641 15204 5675
rect 14436 5574 14470 5608
rect 15452 5592 15475 5602
rect 15475 5592 15486 5602
rect 15452 5566 15486 5592
rect 16424 5783 16458 5817
rect 17164 5783 17198 5817
rect 16240 5729 16255 5749
rect 16255 5729 16274 5749
rect 16608 5745 16629 5749
rect 16629 5745 16642 5749
rect 16240 5715 16274 5729
rect 16608 5715 16642 5745
rect 16332 5651 16366 5681
rect 16332 5647 16361 5651
rect 16361 5647 16366 5651
rect 16792 5667 16826 5681
rect 16792 5647 16797 5667
rect 16797 5647 16826 5667
rect 16980 5715 17014 5749
rect 17256 5721 17288 5749
rect 17288 5721 17290 5749
rect 17256 5715 17290 5721
rect 17164 5647 17198 5681
rect 16430 5580 16464 5614
rect 17446 5598 17469 5608
rect 17469 5598 17480 5608
rect 17446 5572 17480 5598
rect 12017 5395 12051 5429
rect 12109 5395 12143 5429
rect 12201 5395 12235 5429
rect 12293 5395 12327 5429
rect 12385 5395 12419 5429
rect 12477 5395 12511 5429
rect 12569 5395 12603 5429
rect 12661 5395 12695 5429
rect 12753 5395 12787 5429
rect 12845 5395 12879 5429
rect 12937 5395 12971 5429
rect 13029 5395 13063 5429
rect 13121 5395 13155 5429
rect 13213 5395 13247 5429
rect 13305 5395 13339 5429
rect 13397 5395 13431 5429
rect 13489 5395 13523 5429
rect 13975 5403 14009 5437
rect 14067 5403 14101 5437
rect 14159 5403 14193 5437
rect 14251 5403 14285 5437
rect 14343 5403 14377 5437
rect 14435 5403 14469 5437
rect 14527 5403 14561 5437
rect 14619 5403 14653 5437
rect 14711 5403 14745 5437
rect 14803 5403 14837 5437
rect 14895 5403 14929 5437
rect 14987 5403 15021 5437
rect 15079 5403 15113 5437
rect 15171 5403 15205 5437
rect 15263 5403 15297 5437
rect 15355 5403 15389 5437
rect 15447 5403 15481 5437
rect 15971 5409 16005 5443
rect 16061 5409 16095 5443
rect 16153 5409 16187 5443
rect 16245 5409 16279 5443
rect 16337 5409 16371 5443
rect 16429 5409 16463 5443
rect 16521 5409 16555 5443
rect 16613 5409 16647 5443
rect 16705 5409 16739 5443
rect 16797 5409 16831 5443
rect 16889 5409 16923 5443
rect 16981 5409 17015 5443
rect 17073 5409 17107 5443
rect 17165 5409 17199 5443
rect 17257 5409 17291 5443
rect 17349 5409 17383 5443
rect 17441 5409 17475 5443
rect 8224 5227 8258 5257
rect 8224 5223 8253 5227
rect 8253 5223 8258 5227
rect 8684 5243 8718 5257
rect 8684 5223 8689 5243
rect 8689 5223 8718 5243
rect 8872 5291 8906 5325
rect 9148 5297 9180 5325
rect 9180 5297 9182 5325
rect 9148 5291 9182 5297
rect 9056 5223 9090 5257
rect 18331 5379 18365 5413
rect 18423 5379 18457 5413
rect 18515 5379 18549 5413
rect 18607 5379 18641 5413
rect 18699 5379 18733 5413
rect 18791 5379 18825 5413
rect 18883 5379 18917 5413
rect 18975 5379 19009 5413
rect 19067 5379 19101 5413
rect 19159 5379 19193 5413
rect 8322 5156 8356 5190
rect 9338 5174 9361 5184
rect 9361 5174 9372 5184
rect 9338 5148 9372 5174
rect 18608 5188 18642 5222
rect 10075 5077 10109 5111
rect 10167 5077 10201 5111
rect 10259 5077 10293 5111
rect 10351 5077 10385 5111
rect 10443 5077 10477 5111
rect 10535 5077 10569 5111
rect 10627 5077 10661 5111
rect 10719 5077 10753 5111
rect 10811 5077 10845 5111
rect 10903 5077 10937 5111
rect 10995 5077 11029 5111
rect 11087 5077 11121 5111
rect 11179 5077 11213 5111
rect 11271 5077 11305 5111
rect 11363 5077 11397 5111
rect 11455 5077 11489 5111
rect 11547 5077 11581 5111
rect 3909 4979 3943 5013
rect 3999 4979 4033 5013
rect 4091 4979 4125 5013
rect 4183 4979 4217 5013
rect 4275 4979 4309 5013
rect 4367 4979 4401 5013
rect 4459 4979 4493 5013
rect 4551 4979 4585 5013
rect 4643 4979 4677 5013
rect 4735 4979 4769 5013
rect 4827 4979 4861 5013
rect 4919 4979 4953 5013
rect 5011 4979 5045 5013
rect 5103 4979 5137 5013
rect 5195 4979 5229 5013
rect 5287 4979 5321 5013
rect 5379 4979 5413 5013
rect 5859 4979 5893 5013
rect 5951 4979 5985 5013
rect 6043 4979 6077 5013
rect 6135 4979 6169 5013
rect 6227 4979 6261 5013
rect 6319 4979 6353 5013
rect 6411 4979 6445 5013
rect 6503 4979 6537 5013
rect 6595 4979 6629 5013
rect 6687 4979 6721 5013
rect 6779 4979 6813 5013
rect 6871 4979 6905 5013
rect 6963 4979 6997 5013
rect 7055 4979 7089 5013
rect 7147 4979 7181 5013
rect 7239 4979 7273 5013
rect 7331 4979 7365 5013
rect 7861 4985 7895 5019
rect 7953 4985 7987 5019
rect 8045 4985 8079 5019
rect 8137 4985 8171 5019
rect 8229 4985 8263 5019
rect 8321 4985 8355 5019
rect 8413 4985 8447 5019
rect 8505 4985 8539 5019
rect 8597 4985 8631 5019
rect 8689 4985 8723 5019
rect 8781 4985 8815 5019
rect 8873 4985 8907 5019
rect 8965 4985 8999 5019
rect 9057 4985 9091 5019
rect 9149 4985 9183 5019
rect 9241 4985 9275 5019
rect 9333 4985 9367 5019
rect 10438 4907 10472 4941
rect 11178 4907 11212 4941
rect 10254 4853 10269 4873
rect 10269 4853 10288 4873
rect 10622 4869 10643 4873
rect 10643 4869 10656 4873
rect 10254 4839 10288 4853
rect 10622 4839 10656 4869
rect 12257 5033 12291 5067
rect 12345 5033 12379 5067
rect 12437 5033 12471 5067
rect 12529 5033 12563 5067
rect 12621 5033 12655 5067
rect 12713 5033 12747 5067
rect 12805 5033 12839 5067
rect 12897 5033 12931 5067
rect 12989 5033 13023 5067
rect 13081 5033 13115 5067
rect 13173 5033 13207 5067
rect 13265 5033 13299 5067
rect 13357 5033 13391 5067
rect 13449 5033 13483 5067
rect 13541 5033 13575 5067
rect 13633 5033 13667 5067
rect 13725 5033 13759 5067
rect 10346 4775 10380 4805
rect 10346 4771 10375 4775
rect 10375 4771 10380 4775
rect 10806 4791 10840 4805
rect 10806 4771 10811 4791
rect 10811 4771 10840 4791
rect 10994 4839 11028 4873
rect 11270 4845 11302 4873
rect 11302 4845 11304 4873
rect 11270 4839 11304 4845
rect 11178 4771 11212 4805
rect 10446 4706 10480 4740
rect 11454 4722 11483 4732
rect 11483 4722 11494 4732
rect 11454 4696 11494 4722
rect 10075 4533 10109 4567
rect 10167 4533 10201 4567
rect 10259 4533 10293 4567
rect 10351 4533 10385 4567
rect 10443 4533 10477 4567
rect 10535 4533 10569 4567
rect 10627 4533 10661 4567
rect 10719 4533 10753 4567
rect 10811 4533 10845 4567
rect 10903 4533 10937 4567
rect 10995 4533 11029 4567
rect 11087 4533 11121 4567
rect 11179 4533 11213 4567
rect 11271 4533 11305 4567
rect 11363 4533 11397 4567
rect 11455 4533 11489 4567
rect 11547 4533 11581 4567
rect 12708 4863 12742 4897
rect 14257 5027 14291 5061
rect 14347 5027 14381 5061
rect 14439 5027 14473 5061
rect 14531 5027 14565 5061
rect 14623 5027 14657 5061
rect 14715 5027 14749 5061
rect 14807 5027 14841 5061
rect 14899 5027 14933 5061
rect 14991 5027 15025 5061
rect 15083 5027 15117 5061
rect 15175 5027 15209 5061
rect 15267 5027 15301 5061
rect 15359 5027 15393 5061
rect 15451 5027 15485 5061
rect 15543 5027 15577 5061
rect 15635 5027 15669 5061
rect 15727 5027 15761 5061
rect 13448 4863 13482 4897
rect 12524 4809 12539 4829
rect 12539 4809 12558 4829
rect 12892 4825 12913 4829
rect 12913 4825 12926 4829
rect 12524 4795 12558 4809
rect 12892 4795 12926 4825
rect 12616 4731 12650 4761
rect 12616 4727 12645 4731
rect 12645 4727 12650 4731
rect 13076 4747 13110 4761
rect 13076 4727 13081 4747
rect 13081 4727 13110 4747
rect 13264 4795 13298 4829
rect 13540 4801 13572 4829
rect 13572 4801 13574 4829
rect 13540 4795 13574 4801
rect 13448 4727 13482 4761
rect 12714 4660 12748 4694
rect 13730 4678 13753 4688
rect 13753 4678 13764 4688
rect 13730 4652 13764 4678
rect 12257 4489 12291 4523
rect 12345 4489 12379 4523
rect 12437 4489 12471 4523
rect 12529 4489 12563 4523
rect 12621 4489 12655 4523
rect 12713 4489 12747 4523
rect 12805 4489 12839 4523
rect 12897 4489 12931 4523
rect 12989 4489 13023 4523
rect 13081 4489 13115 4523
rect 13173 4489 13207 4523
rect 13265 4489 13299 4523
rect 13357 4489 13391 4523
rect 13449 4489 13483 4523
rect 13541 4489 13575 4523
rect 13633 4489 13667 4523
rect 13725 4489 13759 4523
rect 14710 4857 14744 4891
rect 16281 5009 16315 5043
rect 16369 5009 16403 5043
rect 16461 5009 16495 5043
rect 16553 5009 16587 5043
rect 16645 5009 16679 5043
rect 16737 5009 16771 5043
rect 16829 5009 16863 5043
rect 16921 5009 16955 5043
rect 17013 5009 17047 5043
rect 17105 5009 17139 5043
rect 17197 5009 17231 5043
rect 17289 5009 17323 5043
rect 17381 5009 17415 5043
rect 17473 5009 17507 5043
rect 17565 5009 17599 5043
rect 17657 5009 17691 5043
rect 17749 5009 17783 5043
rect 18432 5104 18470 5108
rect 18432 5070 18437 5104
rect 18437 5070 18470 5104
rect 15450 4857 15484 4891
rect 14526 4803 14541 4823
rect 14541 4803 14560 4823
rect 14894 4819 14915 4823
rect 14915 4819 14928 4823
rect 14526 4789 14560 4803
rect 14894 4789 14928 4819
rect 14618 4725 14652 4755
rect 14618 4721 14647 4725
rect 14647 4721 14652 4725
rect 15078 4741 15112 4755
rect 15078 4721 15083 4741
rect 15083 4721 15112 4741
rect 15266 4789 15300 4823
rect 15542 4795 15574 4823
rect 15574 4795 15576 4823
rect 15542 4789 15576 4795
rect 15450 4721 15484 4755
rect 14716 4654 14750 4688
rect 15732 4672 15755 4682
rect 15755 4672 15766 4682
rect 15732 4646 15766 4672
rect 14257 4483 14291 4517
rect 14347 4483 14381 4517
rect 14439 4483 14473 4517
rect 14531 4483 14565 4517
rect 14623 4483 14657 4517
rect 14715 4483 14749 4517
rect 14807 4483 14841 4517
rect 14899 4483 14933 4517
rect 14991 4483 15025 4517
rect 15083 4483 15117 4517
rect 15175 4483 15209 4517
rect 15267 4483 15301 4517
rect 15359 4483 15393 4517
rect 15451 4483 15485 4517
rect 15543 4483 15577 4517
rect 15635 4483 15669 4517
rect 15727 4483 15761 4517
rect 16732 4839 16766 4873
rect 17472 4839 17506 4873
rect 16548 4785 16563 4805
rect 16563 4785 16582 4805
rect 16916 4801 16937 4805
rect 16937 4801 16950 4805
rect 16548 4771 16582 4785
rect 16916 4771 16950 4801
rect 18690 5183 18711 5194
rect 18711 5183 18724 5194
rect 18690 5160 18724 5183
rect 19064 5013 19102 5042
rect 19064 5004 19095 5013
rect 19095 5004 19102 5013
rect 16640 4707 16674 4737
rect 16640 4703 16669 4707
rect 16669 4703 16674 4707
rect 17100 4723 17134 4737
rect 17100 4703 17105 4723
rect 17105 4703 17134 4723
rect 17288 4771 17322 4805
rect 17564 4777 17596 4805
rect 17596 4777 17598 4805
rect 17564 4771 17598 4777
rect 17472 4703 17506 4737
rect 18331 4835 18365 4869
rect 18423 4835 18457 4869
rect 18515 4835 18549 4869
rect 18607 4835 18641 4869
rect 18699 4835 18733 4869
rect 18791 4835 18825 4869
rect 18883 4835 18917 4869
rect 18975 4835 19009 4869
rect 19067 4835 19101 4869
rect 19159 4835 19193 4869
rect 16738 4636 16772 4670
rect 17754 4654 17777 4664
rect 17777 4654 17788 4664
rect 17754 4628 17788 4654
rect 16281 4465 16315 4499
rect 16369 4465 16403 4499
rect 16461 4465 16495 4499
rect 16553 4465 16587 4499
rect 16645 4465 16679 4499
rect 16737 4465 16771 4499
rect 16829 4465 16863 4499
rect 16921 4465 16955 4499
rect 17013 4465 17047 4499
rect 17105 4465 17139 4499
rect 17197 4465 17231 4499
rect 17289 4465 17323 4499
rect 17381 4465 17415 4499
rect 17473 4465 17507 4499
rect 17565 4465 17599 4499
rect 17657 4465 17691 4499
rect 17749 4465 17783 4499
rect 6023 3323 6057 3357
rect 6111 3323 6145 3357
rect 6203 3323 6237 3357
rect 6295 3323 6329 3357
rect 6148 3088 6182 3122
rect 6244 3091 6278 3124
rect 6244 3090 6278 3091
rect 6023 2779 6057 2813
rect 6111 2779 6145 2813
rect 6203 2779 6237 2813
rect 6295 2779 6329 2813
rect 1745 2271 1779 2305
rect 1835 2271 1869 2305
rect 1927 2271 1961 2305
rect 2019 2271 2053 2305
rect 2111 2271 2145 2305
rect 2203 2271 2237 2305
rect 2295 2271 2329 2305
rect 2387 2271 2421 2305
rect 2479 2271 2513 2305
rect 2571 2271 2605 2305
rect 2663 2271 2697 2305
rect 2755 2271 2789 2305
rect 2847 2271 2881 2305
rect 2939 2271 2973 2305
rect 3031 2271 3065 2305
rect 3123 2271 3157 2305
rect 3215 2271 3249 2305
rect 2198 2101 2232 2135
rect 3815 2267 3849 2301
rect 3905 2267 3939 2301
rect 3997 2267 4031 2301
rect 4089 2267 4123 2301
rect 4181 2267 4215 2301
rect 4273 2267 4307 2301
rect 4365 2267 4399 2301
rect 4457 2267 4491 2301
rect 4549 2267 4583 2301
rect 4641 2267 4675 2301
rect 4733 2267 4767 2301
rect 4825 2267 4859 2301
rect 4917 2267 4951 2301
rect 5009 2267 5043 2301
rect 5101 2267 5135 2301
rect 5193 2267 5227 2301
rect 5285 2267 5319 2301
rect 5771 2267 5805 2301
rect 5857 2267 5891 2301
rect 5949 2267 5983 2301
rect 6041 2267 6075 2301
rect 6133 2267 6167 2301
rect 6225 2267 6259 2301
rect 6317 2267 6351 2301
rect 6409 2267 6443 2301
rect 6501 2267 6535 2301
rect 6593 2267 6627 2301
rect 6685 2267 6719 2301
rect 6777 2267 6811 2301
rect 6869 2267 6903 2301
rect 6961 2267 6995 2301
rect 7053 2267 7087 2301
rect 7145 2267 7179 2301
rect 7237 2267 7271 2301
rect 7769 2273 7803 2307
rect 7859 2273 7893 2307
rect 7951 2273 7985 2307
rect 8043 2273 8077 2307
rect 8135 2273 8169 2307
rect 8227 2273 8261 2307
rect 8319 2273 8353 2307
rect 8411 2273 8445 2307
rect 8503 2273 8537 2307
rect 8595 2273 8629 2307
rect 8687 2273 8721 2307
rect 8779 2273 8813 2307
rect 8871 2273 8905 2307
rect 8963 2273 8997 2307
rect 9055 2273 9089 2307
rect 9147 2273 9181 2307
rect 9239 2273 9273 2307
rect 9725 2273 9759 2307
rect 9811 2273 9845 2307
rect 9903 2273 9937 2307
rect 9995 2273 10029 2307
rect 10087 2273 10121 2307
rect 10179 2273 10213 2307
rect 10271 2273 10305 2307
rect 10363 2273 10397 2307
rect 10455 2273 10489 2307
rect 10547 2273 10581 2307
rect 10639 2273 10673 2307
rect 10731 2273 10765 2307
rect 10823 2273 10857 2307
rect 10915 2273 10949 2307
rect 11007 2273 11041 2307
rect 11099 2273 11133 2307
rect 11191 2273 11225 2307
rect 11713 2273 11747 2307
rect 11803 2273 11837 2307
rect 11895 2273 11929 2307
rect 11987 2273 12021 2307
rect 12079 2273 12113 2307
rect 12171 2273 12205 2307
rect 12263 2273 12297 2307
rect 12355 2273 12389 2307
rect 12447 2273 12481 2307
rect 12539 2273 12573 2307
rect 12631 2273 12665 2307
rect 12723 2273 12757 2307
rect 12815 2273 12849 2307
rect 12907 2273 12941 2307
rect 12999 2273 13033 2307
rect 13091 2273 13125 2307
rect 13183 2273 13217 2307
rect 13667 2273 13701 2307
rect 13755 2273 13789 2307
rect 13847 2273 13881 2307
rect 13939 2273 13973 2307
rect 14031 2273 14065 2307
rect 14123 2273 14157 2307
rect 14215 2273 14249 2307
rect 14307 2273 14341 2307
rect 14399 2273 14433 2307
rect 14491 2273 14525 2307
rect 14583 2273 14617 2307
rect 14675 2273 14709 2307
rect 14767 2273 14801 2307
rect 14859 2273 14893 2307
rect 14951 2273 14985 2307
rect 15043 2273 15077 2307
rect 15135 2273 15169 2307
rect 15729 2273 15763 2307
rect 15819 2273 15853 2307
rect 15911 2273 15945 2307
rect 16003 2273 16037 2307
rect 16095 2273 16129 2307
rect 16187 2273 16221 2307
rect 16279 2273 16313 2307
rect 16371 2273 16405 2307
rect 16463 2273 16497 2307
rect 16555 2273 16589 2307
rect 16647 2273 16681 2307
rect 16739 2273 16773 2307
rect 16831 2273 16865 2307
rect 16923 2273 16957 2307
rect 17015 2273 17049 2307
rect 17107 2273 17141 2307
rect 17199 2273 17233 2307
rect 2938 2101 2972 2135
rect 2014 2047 2029 2067
rect 2029 2047 2048 2067
rect 2382 2063 2403 2067
rect 2403 2063 2416 2067
rect 2014 2033 2048 2047
rect 2382 2033 2416 2063
rect 2106 1969 2140 1999
rect 2106 1965 2135 1969
rect 2135 1965 2140 1969
rect 2566 1985 2600 1999
rect 2566 1965 2571 1985
rect 2571 1965 2600 1985
rect 2754 2033 2788 2067
rect 3030 2039 3062 2067
rect 3062 2039 3064 2067
rect 3030 2033 3064 2039
rect 2938 1965 2972 1999
rect 2206 1900 2240 1934
rect 3214 1916 3243 1926
rect 3243 1916 3254 1926
rect 3214 1890 3254 1916
rect 1745 1727 1779 1761
rect 1835 1727 1869 1761
rect 1927 1727 1961 1761
rect 2019 1727 2053 1761
rect 2111 1727 2145 1761
rect 2203 1727 2237 1761
rect 2295 1727 2329 1761
rect 2387 1727 2421 1761
rect 2479 1727 2513 1761
rect 2571 1727 2605 1761
rect 2663 1727 2697 1761
rect 2755 1727 2789 1761
rect 2847 1727 2881 1761
rect 2939 1727 2973 1761
rect 3031 1727 3065 1761
rect 3123 1727 3157 1761
rect 3215 1727 3249 1761
rect 4268 2097 4302 2131
rect 5008 2097 5042 2131
rect 4084 2043 4099 2063
rect 4099 2043 4118 2063
rect 4452 2059 4473 2063
rect 4473 2059 4486 2063
rect 4084 2029 4118 2043
rect 4452 2029 4486 2059
rect 4176 1965 4210 1995
rect 4176 1961 4205 1965
rect 4205 1961 4210 1965
rect 4636 1981 4670 1995
rect 4636 1961 4641 1981
rect 4641 1961 4670 1981
rect 4824 2029 4858 2063
rect 5100 2035 5132 2063
rect 5132 2035 5134 2063
rect 5100 2029 5134 2035
rect 5008 1961 5042 1995
rect 4274 1894 4308 1928
rect 5290 1912 5313 1922
rect 5313 1912 5324 1922
rect 5290 1886 5324 1912
rect 6220 2097 6254 2131
rect 6960 2097 6994 2131
rect 6036 2043 6051 2063
rect 6051 2043 6070 2063
rect 6404 2059 6425 2063
rect 6425 2059 6438 2063
rect 6036 2029 6070 2043
rect 6404 2029 6438 2059
rect 6128 1965 6162 1995
rect 6128 1961 6157 1965
rect 6157 1961 6162 1965
rect 6588 1981 6622 1995
rect 6588 1961 6593 1981
rect 6593 1961 6622 1981
rect 6776 2029 6810 2063
rect 7052 2035 7084 2063
rect 7084 2035 7086 2063
rect 7052 2029 7086 2035
rect 6960 1961 6994 1995
rect 6226 1894 6260 1928
rect 7242 1912 7265 1922
rect 7265 1912 7276 1922
rect 7242 1886 7276 1912
rect 8222 2103 8256 2137
rect 8962 2103 8996 2137
rect 8038 2049 8053 2069
rect 8053 2049 8072 2069
rect 8406 2065 8427 2069
rect 8427 2065 8440 2069
rect 8038 2035 8072 2049
rect 8406 2035 8440 2065
rect 8130 1971 8164 2001
rect 8130 1967 8159 1971
rect 8159 1967 8164 1971
rect 8590 1987 8624 2001
rect 8590 1967 8595 1987
rect 8595 1967 8624 1987
rect 8778 2035 8812 2069
rect 9054 2041 9086 2069
rect 9086 2041 9088 2069
rect 9054 2035 9088 2041
rect 8962 1967 8996 2001
rect 8228 1900 8262 1934
rect 9244 1918 9267 1928
rect 9267 1918 9278 1928
rect 9244 1892 9278 1918
rect 10174 2103 10208 2137
rect 10914 2103 10948 2137
rect 9990 2049 10005 2069
rect 10005 2049 10024 2069
rect 10358 2065 10379 2069
rect 10379 2065 10392 2069
rect 9990 2035 10024 2049
rect 10358 2035 10392 2065
rect 10082 1971 10116 2001
rect 10082 1967 10111 1971
rect 10111 1967 10116 1971
rect 10542 1987 10576 2001
rect 10542 1967 10547 1987
rect 10547 1967 10576 1987
rect 10730 2035 10764 2069
rect 11006 2041 11038 2069
rect 11038 2041 11040 2069
rect 11006 2035 11040 2041
rect 10914 1967 10948 2001
rect 10180 1900 10214 1934
rect 11196 1918 11219 1928
rect 11219 1918 11230 1928
rect 11196 1892 11230 1918
rect 12166 2103 12200 2137
rect 12906 2103 12940 2137
rect 11982 2049 11997 2069
rect 11997 2049 12016 2069
rect 12350 2065 12371 2069
rect 12371 2065 12384 2069
rect 11982 2035 12016 2049
rect 12350 2035 12384 2065
rect 12074 1971 12108 2001
rect 12074 1967 12103 1971
rect 12103 1967 12108 1971
rect 12534 1987 12568 2001
rect 12534 1967 12539 1987
rect 12539 1967 12568 1987
rect 12722 2035 12756 2069
rect 12998 2041 13030 2069
rect 13030 2041 13032 2069
rect 12998 2035 13032 2041
rect 12906 1967 12940 2001
rect 12172 1900 12206 1934
rect 13188 1918 13211 1928
rect 13211 1918 13222 1928
rect 13188 1892 13222 1918
rect 14118 2103 14152 2137
rect 14858 2103 14892 2137
rect 13934 2049 13949 2069
rect 13949 2049 13968 2069
rect 14302 2065 14323 2069
rect 14323 2065 14336 2069
rect 13934 2035 13968 2049
rect 14302 2035 14336 2065
rect 14026 1971 14060 2001
rect 14026 1967 14055 1971
rect 14055 1967 14060 1971
rect 14486 1987 14520 2001
rect 14486 1967 14491 1987
rect 14491 1967 14520 1987
rect 14674 2035 14708 2069
rect 14950 2041 14982 2069
rect 14982 2041 14984 2069
rect 14950 2035 14984 2041
rect 14858 1967 14892 2001
rect 14124 1900 14158 1934
rect 15140 1918 15163 1928
rect 15163 1918 15174 1928
rect 15140 1892 15174 1918
rect 16182 2103 16216 2137
rect 16922 2103 16956 2137
rect 15998 2049 16013 2069
rect 16013 2049 16032 2069
rect 16366 2065 16387 2069
rect 16387 2065 16400 2069
rect 15998 2035 16032 2049
rect 16366 2035 16400 2065
rect 16090 1971 16124 2001
rect 16090 1967 16119 1971
rect 16119 1967 16124 1971
rect 16550 1987 16584 2001
rect 16550 1967 16555 1987
rect 16555 1967 16584 1987
rect 16738 2035 16772 2069
rect 17014 2041 17046 2069
rect 17046 2041 17048 2069
rect 17014 2035 17048 2041
rect 16922 1967 16956 2001
rect 16188 1900 16222 1934
rect 17204 1918 17227 1928
rect 17227 1918 17238 1928
rect 17204 1892 17238 1918
rect 3815 1723 3849 1757
rect 3905 1723 3939 1757
rect 3997 1723 4031 1757
rect 4089 1723 4123 1757
rect 4181 1723 4215 1757
rect 4273 1723 4307 1757
rect 4365 1723 4399 1757
rect 4457 1723 4491 1757
rect 4549 1723 4583 1757
rect 4641 1723 4675 1757
rect 4733 1723 4767 1757
rect 4825 1723 4859 1757
rect 4917 1723 4951 1757
rect 5009 1723 5043 1757
rect 5101 1723 5135 1757
rect 5193 1723 5227 1757
rect 5285 1723 5319 1757
rect 5771 1723 5805 1757
rect 5857 1723 5891 1757
rect 5949 1723 5983 1757
rect 6041 1723 6075 1757
rect 6133 1723 6167 1757
rect 6225 1723 6259 1757
rect 6317 1723 6351 1757
rect 6409 1723 6443 1757
rect 6501 1723 6535 1757
rect 6593 1723 6627 1757
rect 6685 1723 6719 1757
rect 6777 1723 6811 1757
rect 6869 1723 6903 1757
rect 6961 1723 6995 1757
rect 7053 1723 7087 1757
rect 7145 1723 7179 1757
rect 7237 1723 7271 1757
rect 7769 1729 7803 1763
rect 7859 1729 7893 1763
rect 7951 1729 7985 1763
rect 8043 1729 8077 1763
rect 8135 1729 8169 1763
rect 8227 1729 8261 1763
rect 8319 1729 8353 1763
rect 8411 1729 8445 1763
rect 8503 1729 8537 1763
rect 8595 1729 8629 1763
rect 8687 1729 8721 1763
rect 8779 1729 8813 1763
rect 8871 1729 8905 1763
rect 8963 1729 8997 1763
rect 9055 1729 9089 1763
rect 9147 1729 9181 1763
rect 9239 1729 9273 1763
rect 9725 1729 9759 1763
rect 9811 1729 9845 1763
rect 9903 1729 9937 1763
rect 9995 1729 10029 1763
rect 10087 1729 10121 1763
rect 10179 1729 10213 1763
rect 10271 1729 10305 1763
rect 10363 1729 10397 1763
rect 10455 1729 10489 1763
rect 10547 1729 10581 1763
rect 10639 1729 10673 1763
rect 10731 1729 10765 1763
rect 10823 1729 10857 1763
rect 10915 1729 10949 1763
rect 11007 1729 11041 1763
rect 11099 1729 11133 1763
rect 11191 1729 11225 1763
rect 11713 1729 11747 1763
rect 11803 1729 11837 1763
rect 11895 1729 11929 1763
rect 11987 1729 12021 1763
rect 12079 1729 12113 1763
rect 12171 1729 12205 1763
rect 12263 1729 12297 1763
rect 12355 1729 12389 1763
rect 12447 1729 12481 1763
rect 12539 1729 12573 1763
rect 12631 1729 12665 1763
rect 12723 1729 12757 1763
rect 12815 1729 12849 1763
rect 12907 1729 12941 1763
rect 12999 1729 13033 1763
rect 13091 1729 13125 1763
rect 13183 1729 13217 1763
rect 13667 1729 13701 1763
rect 13755 1729 13789 1763
rect 13847 1729 13881 1763
rect 13939 1729 13973 1763
rect 14031 1729 14065 1763
rect 14123 1729 14157 1763
rect 14215 1729 14249 1763
rect 14307 1729 14341 1763
rect 14399 1729 14433 1763
rect 14491 1729 14525 1763
rect 14583 1729 14617 1763
rect 14675 1729 14709 1763
rect 14767 1729 14801 1763
rect 14859 1729 14893 1763
rect 14951 1729 14985 1763
rect 15043 1729 15077 1763
rect 15135 1729 15169 1763
rect 15729 1729 15763 1763
rect 15819 1729 15853 1763
rect 15911 1729 15945 1763
rect 16003 1729 16037 1763
rect 16095 1729 16129 1763
rect 16187 1729 16221 1763
rect 16279 1729 16313 1763
rect 16371 1729 16405 1763
rect 16463 1729 16497 1763
rect 16555 1729 16589 1763
rect 16647 1729 16681 1763
rect 16739 1729 16773 1763
rect 16831 1729 16865 1763
rect 16923 1729 16957 1763
rect 17015 1729 17049 1763
rect 17107 1729 17141 1763
rect 17199 1729 17233 1763
<< metal1 >>
rect 18590 44096 19128 44168
rect 18590 43898 18768 44096
rect 18962 43898 19128 44096
rect 18590 43828 19128 43898
rect 18548 43481 18644 43510
rect 18548 43447 18579 43481
rect 18613 43447 18644 43481
rect 18548 43391 18644 43447
rect 18548 43357 18579 43391
rect 18613 43357 18644 43391
rect 18548 43299 18644 43357
rect 18548 43265 18579 43299
rect 18613 43265 18644 43299
rect 18548 43207 18644 43265
rect 18866 43294 18936 43828
rect 18866 43258 18882 43294
rect 18916 43258 18936 43294
rect 18866 43244 18936 43258
rect 19092 43481 19188 43510
rect 19092 43447 19123 43481
rect 19157 43447 19188 43481
rect 19092 43391 19188 43447
rect 19092 43357 19123 43391
rect 19157 43357 19188 43391
rect 19092 43299 19188 43357
rect 19092 43265 19123 43299
rect 19157 43265 19188 43299
rect 18548 43173 18579 43207
rect 18613 43173 18644 43207
rect 18548 43115 18644 43173
rect 18548 43081 18579 43115
rect 18613 43081 18644 43115
rect 18548 43023 18644 43081
rect 18548 42989 18579 43023
rect 18613 42989 18644 43023
rect 18548 42931 18644 42989
rect 18548 42897 18579 42931
rect 18613 42897 18644 42931
rect 18548 42839 18644 42897
rect 18548 42820 18579 42839
rect 18613 42820 18644 42839
rect 18548 42762 18562 42820
rect 18624 42762 18644 42820
rect 18548 42747 18644 42762
rect 18548 42713 18579 42747
rect 18613 42713 18644 42747
rect 18548 42655 18644 42713
rect 18548 42621 18579 42655
rect 18613 42621 18644 42655
rect 18548 42563 18644 42621
rect 18548 42529 18579 42563
rect 18613 42529 18644 42563
rect 18548 42471 18644 42529
rect 18548 42437 18579 42471
rect 18613 42437 18644 42471
rect 18548 42379 18644 42437
rect 18548 42345 18579 42379
rect 18613 42345 18644 42379
rect 18548 42287 18644 42345
rect 18548 42253 18579 42287
rect 18613 42253 18644 42287
rect 18548 42195 18644 42253
rect 18548 42161 18579 42195
rect 18613 42161 18644 42195
rect 18548 42103 18644 42161
rect 18548 42069 18579 42103
rect 18613 42069 18644 42103
rect 18548 42011 18644 42069
rect 19092 43207 19188 43265
rect 19092 43173 19123 43207
rect 19157 43173 19188 43207
rect 19092 43115 19188 43173
rect 19092 43081 19123 43115
rect 19157 43081 19188 43115
rect 19092 43023 19188 43081
rect 19092 42989 19123 43023
rect 19157 42989 19188 43023
rect 19092 42931 19188 42989
rect 19092 42897 19123 42931
rect 19157 42897 19188 42931
rect 19092 42839 19188 42897
rect 19092 42805 19123 42839
rect 19157 42805 19188 42839
rect 19092 42782 19188 42805
rect 19092 42747 19124 42782
rect 19092 42713 19123 42747
rect 19186 42724 19188 42782
rect 19157 42713 19188 42724
rect 19092 42655 19188 42713
rect 19092 42621 19123 42655
rect 19157 42621 19188 42655
rect 19092 42563 19188 42621
rect 19092 42529 19123 42563
rect 19157 42529 19188 42563
rect 19092 42471 19188 42529
rect 19092 42437 19123 42471
rect 19157 42437 19188 42471
rect 19092 42379 19188 42437
rect 19092 42345 19123 42379
rect 19157 42345 19188 42379
rect 19092 42287 19188 42345
rect 19092 42253 19123 42287
rect 19157 42253 19188 42287
rect 19092 42195 19188 42253
rect 19092 42161 19123 42195
rect 19157 42161 19188 42195
rect 19092 42103 19188 42161
rect 19092 42069 19123 42103
rect 19157 42069 19188 42103
rect 18548 41977 18579 42011
rect 18613 41977 18644 42011
rect 18548 41948 18644 41977
rect 18856 42024 18938 42050
rect 18856 41990 18886 42024
rect 18920 41990 18938 42024
rect 18532 41495 18628 41524
rect 18532 41461 18563 41495
rect 18597 41461 18628 41495
rect 18532 41403 18628 41461
rect 18532 41369 18563 41403
rect 18597 41369 18628 41403
rect 18532 41311 18628 41369
rect 18856 41398 18938 41990
rect 19092 42011 19188 42069
rect 19092 41977 19123 42011
rect 19157 41977 19188 42011
rect 19092 41948 19188 41977
rect 18856 41364 18868 41398
rect 18902 41364 18938 41398
rect 18856 41346 18938 41364
rect 19076 41495 19172 41524
rect 19076 41461 19107 41495
rect 19141 41461 19172 41495
rect 19076 41403 19172 41461
rect 19076 41369 19107 41403
rect 19141 41369 19172 41403
rect 18532 41277 18563 41311
rect 18597 41277 18628 41311
rect 18532 41219 18628 41277
rect 18532 41185 18563 41219
rect 18597 41185 18628 41219
rect 18532 41127 18628 41185
rect 18532 41093 18563 41127
rect 18597 41093 18628 41127
rect 18532 41035 18628 41093
rect 18532 41001 18563 41035
rect 18597 41001 18628 41035
rect 18532 40948 18628 41001
rect 18532 40890 18540 40948
rect 18602 40890 18628 40948
rect 18532 40851 18628 40890
rect 18532 40817 18563 40851
rect 18597 40817 18628 40851
rect 18532 40759 18628 40817
rect 18532 40725 18563 40759
rect 18597 40725 18628 40759
rect 18532 40667 18628 40725
rect 18532 40633 18563 40667
rect 18597 40633 18628 40667
rect 18532 40575 18628 40633
rect 18532 40541 18563 40575
rect 18597 40541 18628 40575
rect 18532 40483 18628 40541
rect 19076 41311 19172 41369
rect 19076 41277 19107 41311
rect 19141 41277 19172 41311
rect 19076 41219 19172 41277
rect 19076 41185 19107 41219
rect 19141 41185 19172 41219
rect 19076 41127 19172 41185
rect 19076 41093 19107 41127
rect 19141 41093 19172 41127
rect 19076 41035 19172 41093
rect 19076 41001 19107 41035
rect 19141 41001 19172 41035
rect 19076 40943 19172 41001
rect 19076 40940 19107 40943
rect 19141 40940 19172 40943
rect 19076 40882 19106 40940
rect 19168 40882 19172 40940
rect 19076 40851 19172 40882
rect 19076 40817 19107 40851
rect 19141 40817 19172 40851
rect 19076 40759 19172 40817
rect 19076 40725 19107 40759
rect 19141 40725 19172 40759
rect 19076 40667 19172 40725
rect 19076 40633 19107 40667
rect 19141 40633 19172 40667
rect 19076 40575 19172 40633
rect 19076 40541 19107 40575
rect 19141 40541 19172 40575
rect 18532 40449 18563 40483
rect 18597 40449 18628 40483
rect 18532 40391 18628 40449
rect 18532 40357 18563 40391
rect 18597 40357 18628 40391
rect 18532 40299 18628 40357
rect 18532 40265 18563 40299
rect 18597 40265 18628 40299
rect 18532 40236 18628 40265
rect 18846 40468 18914 40510
rect 18846 40434 18870 40468
rect 18904 40434 18914 40468
rect 18540 39699 18636 39728
rect 18540 39665 18571 39699
rect 18605 39665 18636 39699
rect 18540 39607 18636 39665
rect 18540 39573 18571 39607
rect 18605 39573 18636 39607
rect 18540 39515 18636 39573
rect 18846 39606 18914 40434
rect 19076 40483 19172 40541
rect 19076 40449 19107 40483
rect 19141 40449 19172 40483
rect 19076 40391 19172 40449
rect 19076 40357 19107 40391
rect 19141 40357 19172 40391
rect 19076 40299 19172 40357
rect 19076 40265 19107 40299
rect 19141 40265 19172 40299
rect 19076 40236 19172 40265
rect 18846 39570 18862 39606
rect 18896 39570 18914 39606
rect 18846 39554 18914 39570
rect 19084 39699 19180 39728
rect 19084 39665 19115 39699
rect 19149 39665 19180 39699
rect 19084 39607 19180 39665
rect 19084 39573 19115 39607
rect 19149 39573 19180 39607
rect 18540 39481 18571 39515
rect 18605 39481 18636 39515
rect 18540 39423 18636 39481
rect 18540 39389 18571 39423
rect 18605 39389 18636 39423
rect 18540 39331 18636 39389
rect 18540 39320 18571 39331
rect 18605 39320 18636 39331
rect 18540 39262 18564 39320
rect 18626 39262 18636 39320
rect 18540 39239 18636 39262
rect 18540 39205 18571 39239
rect 18605 39205 18636 39239
rect 18540 39147 18636 39205
rect 18540 39113 18571 39147
rect 18605 39113 18636 39147
rect 19084 39515 19180 39573
rect 19084 39481 19115 39515
rect 19149 39481 19180 39515
rect 19084 39423 19180 39481
rect 19084 39389 19115 39423
rect 19149 39389 19180 39423
rect 19084 39331 19180 39389
rect 19084 39316 19115 39331
rect 19149 39316 19180 39331
rect 19084 39258 19106 39316
rect 19168 39258 19180 39316
rect 19084 39239 19180 39258
rect 19084 39205 19115 39239
rect 19149 39205 19180 39239
rect 19084 39147 19180 39205
rect 18540 39055 18636 39113
rect 18540 39021 18571 39055
rect 18605 39021 18636 39055
rect 18540 38963 18636 39021
rect 18540 38929 18571 38963
rect 18605 38929 18636 38963
rect 18540 38871 18636 38929
rect 18540 38837 18571 38871
rect 18605 38837 18636 38871
rect 18540 38808 18636 38837
rect 18864 39090 18946 39114
rect 18864 39056 18876 39090
rect 18910 39056 18946 39090
rect 18554 38437 18650 38466
rect 18554 38403 18585 38437
rect 18619 38403 18650 38437
rect 18554 38345 18650 38403
rect 18554 38311 18585 38345
rect 18619 38311 18650 38345
rect 18554 38253 18650 38311
rect 18864 38340 18946 39056
rect 19084 39113 19115 39147
rect 19149 39113 19180 39147
rect 19084 39055 19180 39113
rect 19084 39021 19115 39055
rect 19149 39021 19180 39055
rect 19084 38963 19180 39021
rect 19084 38929 19115 38963
rect 19149 38929 19180 38963
rect 19084 38871 19180 38929
rect 19084 38837 19115 38871
rect 19149 38837 19180 38871
rect 19084 38808 19180 38837
rect 18864 38306 18886 38340
rect 18920 38306 18946 38340
rect 18864 38284 18946 38306
rect 19098 38437 19194 38466
rect 19098 38403 19129 38437
rect 19163 38403 19194 38437
rect 19098 38345 19194 38403
rect 19098 38311 19129 38345
rect 19163 38311 19194 38345
rect 18554 38219 18585 38253
rect 18619 38219 18650 38253
rect 18554 38161 18650 38219
rect 18554 38127 18585 38161
rect 18619 38127 18650 38161
rect 18554 38124 18650 38127
rect 18554 38066 18572 38124
rect 18634 38066 18650 38124
rect 18554 38035 18585 38066
rect 18619 38035 18650 38066
rect 18554 37977 18650 38035
rect 18554 37943 18585 37977
rect 18619 37943 18650 37977
rect 19098 38253 19194 38311
rect 19098 38219 19129 38253
rect 19163 38219 19194 38253
rect 19098 38161 19194 38219
rect 19098 38140 19129 38161
rect 19163 38140 19194 38161
rect 19098 38082 19122 38140
rect 19184 38082 19194 38140
rect 19098 38069 19194 38082
rect 19098 38035 19129 38069
rect 19163 38035 19194 38069
rect 19098 37977 19194 38035
rect 18554 37885 18650 37943
rect 18554 37851 18585 37885
rect 18619 37851 18650 37885
rect 18554 37793 18650 37851
rect 18554 37759 18585 37793
rect 18619 37759 18650 37793
rect 18554 37730 18650 37759
rect 18872 37794 18934 37954
rect 18872 37760 18888 37794
rect 18922 37760 18934 37794
rect 18566 37283 18662 37312
rect 18566 37249 18597 37283
rect 18631 37249 18662 37283
rect 18566 37195 18662 37249
rect 18872 37198 18934 37760
rect 19098 37943 19129 37977
rect 19163 37943 19194 37977
rect 19098 37885 19194 37943
rect 19098 37851 19129 37885
rect 19163 37851 19194 37885
rect 19098 37793 19194 37851
rect 19098 37759 19129 37793
rect 19163 37759 19194 37793
rect 19098 37730 19194 37759
rect 19110 37283 19206 37312
rect 19110 37249 19141 37283
rect 19175 37249 19206 37283
rect 18566 37161 18597 37195
rect 18631 37161 18662 37195
rect 18566 37103 18662 37161
rect 18870 37192 18952 37198
rect 18870 37158 18892 37192
rect 18926 37158 18952 37192
rect 18870 37144 18952 37158
rect 19110 37195 19206 37249
rect 19110 37161 19141 37195
rect 19175 37161 19206 37195
rect 18566 37069 18597 37103
rect 18631 37069 18662 37103
rect 18566 37054 18662 37069
rect 18566 36996 18580 37054
rect 18642 36996 18662 37054
rect 18566 36977 18597 36996
rect 18631 36977 18662 36996
rect 18566 36919 18662 36977
rect 19110 37103 19206 37161
rect 19110 37069 19141 37103
rect 19175 37069 19206 37103
rect 19110 37044 19206 37069
rect 19110 36986 19128 37044
rect 19190 36986 19206 37044
rect 19110 36977 19141 36986
rect 19175 36977 19206 36986
rect 18566 36885 18597 36919
rect 18631 36885 18662 36919
rect 18566 36827 18662 36885
rect 18886 36920 18950 36928
rect 18886 36884 18900 36920
rect 18934 36884 18950 36920
rect 18886 36868 18950 36884
rect 19110 36919 19206 36977
rect 19110 36885 19141 36919
rect 19175 36885 19206 36919
rect 18566 36793 18597 36827
rect 18631 36793 18662 36827
rect 18566 36764 18662 36793
rect 18574 36399 18670 36428
rect 18574 36365 18605 36399
rect 18639 36365 18670 36399
rect 18574 36307 18670 36365
rect 18574 36273 18605 36307
rect 18639 36273 18670 36307
rect 18574 36256 18670 36273
rect 18574 36200 18598 36256
rect 18652 36200 18670 36256
rect 18898 36236 18944 36868
rect 19110 36827 19206 36885
rect 19110 36793 19141 36827
rect 19175 36793 19206 36827
rect 19110 36764 19206 36793
rect 19118 36399 19214 36428
rect 19118 36365 19149 36399
rect 19183 36365 19214 36399
rect 19118 36307 19214 36365
rect 19118 36284 19149 36307
rect 19183 36284 19214 36307
rect 18574 36181 18605 36200
rect 18639 36181 18670 36200
rect 18574 36123 18670 36181
rect 18890 36226 18954 36236
rect 18890 36190 18904 36226
rect 18940 36190 18954 36226
rect 18890 36176 18954 36190
rect 19118 36228 19142 36284
rect 19200 36228 19214 36284
rect 19118 36215 19214 36228
rect 19118 36181 19149 36215
rect 19183 36181 19214 36215
rect 18574 36089 18605 36123
rect 18639 36089 18670 36123
rect 18574 36060 18670 36089
rect 18896 36130 18958 36146
rect 18896 36094 18904 36130
rect 18948 36094 18958 36130
rect 18896 36080 18958 36094
rect 19118 36123 19214 36181
rect 19118 36089 19149 36123
rect 19183 36089 19214 36123
rect 18911 35879 18953 36080
rect 19118 36060 19214 36089
rect 18870 35837 18953 35879
rect 18870 35518 18912 35837
rect 18870 35476 19094 35518
rect 18598 35011 18694 35040
rect 18598 34977 18629 35011
rect 18663 34977 18694 35011
rect 18598 34919 18694 34977
rect 18598 34885 18629 34919
rect 18663 34885 18694 34919
rect 18598 34827 18694 34885
rect 18598 34793 18629 34827
rect 18663 34793 18694 34827
rect 18598 34735 18694 34793
rect 18598 34701 18629 34735
rect 18663 34701 18694 34735
rect 18598 34643 18694 34701
rect 18598 34609 18629 34643
rect 18663 34609 18694 34643
rect 18598 34551 18694 34609
rect 18598 34517 18629 34551
rect 18663 34517 18694 34551
rect 18598 34459 18694 34517
rect 18598 34425 18629 34459
rect 18663 34425 18694 34459
rect 18598 34367 18694 34425
rect 18598 34333 18629 34367
rect 18663 34333 18694 34367
rect 18598 34275 18694 34333
rect 18823 34914 18885 34929
rect 18823 34880 18836 34914
rect 18870 34880 18885 34914
rect 18823 34347 18885 34880
rect 19054 34674 19094 35476
rect 19142 35011 19238 35040
rect 19142 34977 19173 35011
rect 19207 34977 19238 35011
rect 19142 34919 19238 34977
rect 19142 34885 19173 34919
rect 19207 34885 19238 34919
rect 19142 34827 19238 34885
rect 19142 34793 19173 34827
rect 19207 34793 19238 34827
rect 19142 34735 19238 34793
rect 19142 34701 19173 34735
rect 19207 34701 19238 34735
rect 19050 34634 19106 34674
rect 19050 34600 19058 34634
rect 19092 34600 19106 34634
rect 19050 34578 19106 34600
rect 19142 34643 19238 34701
rect 19142 34609 19173 34643
rect 19207 34609 19238 34643
rect 19142 34551 19238 34609
rect 19142 34517 19173 34551
rect 19207 34517 19238 34551
rect 19142 34459 19238 34517
rect 19142 34425 19173 34459
rect 19207 34425 19238 34459
rect 19142 34367 19238 34425
rect 18823 34285 19032 34347
rect 18598 34241 18629 34275
rect 18663 34241 18694 34275
rect 18598 34183 18694 34241
rect 18598 34149 18629 34183
rect 18663 34149 18694 34183
rect 18598 34132 18694 34149
rect 18861 34181 18907 34193
rect 18861 34147 18867 34181
rect 18901 34147 18907 34181
rect 18861 34135 18907 34147
rect 18598 34066 18618 34132
rect 18684 34066 18694 34132
rect 18598 34057 18629 34066
rect 18663 34057 18694 34066
rect 18598 33999 18694 34057
rect 18793 34094 18839 34106
rect 18793 34060 18799 34094
rect 18833 34060 18839 34094
rect 18793 34048 18839 34060
rect 18598 33965 18629 33999
rect 18663 33965 18694 33999
rect 18598 33907 18694 33965
rect 18598 33873 18629 33907
rect 18663 33873 18694 33907
rect 18598 33815 18694 33873
rect 18598 33781 18629 33815
rect 18663 33781 18694 33815
rect 18802 33792 18830 34048
rect 18598 33723 18694 33781
rect 18793 33780 18839 33792
rect 18793 33746 18799 33780
rect 18833 33746 18839 33780
rect 18793 33734 18839 33746
rect 18598 33689 18629 33723
rect 18663 33689 18694 33723
rect 18598 33631 18694 33689
rect 18598 33597 18629 33631
rect 18663 33597 18694 33631
rect 18598 33539 18694 33597
rect 18598 33505 18629 33539
rect 18663 33505 18694 33539
rect 18598 33447 18694 33505
rect 18598 33413 18629 33447
rect 18663 33413 18694 33447
rect 18598 33355 18694 33413
rect 18802 33372 18830 33734
rect 18870 33689 18898 34135
rect 18861 33677 18907 33689
rect 18861 33643 18867 33677
rect 18901 33643 18907 33677
rect 18861 33631 18907 33643
rect 18870 33451 18898 33631
rect 18970 33586 19032 34285
rect 19142 34333 19173 34367
rect 19207 34333 19238 34367
rect 19142 34275 19238 34333
rect 19142 34241 19173 34275
rect 19207 34241 19238 34275
rect 19142 34183 19238 34241
rect 19142 34149 19173 34183
rect 19207 34149 19238 34183
rect 19142 34142 19238 34149
rect 19142 34076 19160 34142
rect 19226 34076 19238 34142
rect 19142 34057 19173 34076
rect 19207 34057 19238 34076
rect 19142 33999 19238 34057
rect 19142 33965 19173 33999
rect 19207 33965 19238 33999
rect 19142 33907 19238 33965
rect 19142 33873 19173 33907
rect 19207 33873 19238 33907
rect 19142 33815 19238 33873
rect 19142 33781 19173 33815
rect 19207 33781 19238 33815
rect 19142 33723 19238 33781
rect 19142 33689 19173 33723
rect 19207 33689 19238 33723
rect 19142 33631 19238 33689
rect 19142 33597 19173 33631
rect 19207 33597 19238 33631
rect 18970 33524 19046 33586
rect 18970 33484 18988 33524
rect 19028 33484 19046 33524
rect 18970 33466 19046 33484
rect 19142 33539 19238 33597
rect 19142 33505 19173 33539
rect 19207 33505 19238 33539
rect 18861 33439 18907 33451
rect 18861 33405 18867 33439
rect 18901 33405 18907 33439
rect 18861 33393 18907 33405
rect 19142 33447 19238 33505
rect 19142 33413 19173 33447
rect 19207 33413 19238 33447
rect 18598 33321 18629 33355
rect 18663 33321 18694 33355
rect 18598 33263 18694 33321
rect 18793 33360 18839 33372
rect 18793 33326 18799 33360
rect 18833 33326 18839 33360
rect 18793 33314 18839 33326
rect 19142 33355 19238 33413
rect 19142 33321 19173 33355
rect 19207 33321 19238 33355
rect 18598 33229 18629 33263
rect 18663 33229 18694 33263
rect 18598 33200 18694 33229
rect 18879 33266 19025 33293
rect 18879 33232 18940 33266
rect 18976 33232 19025 33266
rect 18879 33070 19025 33232
rect 19142 33263 19238 33321
rect 19142 33229 19173 33263
rect 19207 33229 19238 33263
rect 19142 33200 19238 33229
rect 18879 33042 19102 33070
rect 18994 33032 19102 33042
rect 18598 32729 18694 32758
rect 18598 32695 18629 32729
rect 18663 32695 18694 32729
rect 18598 32637 18694 32695
rect 18598 32603 18629 32637
rect 18663 32603 18694 32637
rect 18598 32545 18694 32603
rect 18598 32511 18629 32545
rect 18663 32511 18694 32545
rect 18598 32453 18694 32511
rect 18598 32419 18629 32453
rect 18663 32419 18694 32453
rect 18598 32361 18694 32419
rect 18598 32327 18629 32361
rect 18663 32327 18694 32361
rect 18598 32269 18694 32327
rect 18598 32235 18629 32269
rect 18663 32235 18694 32269
rect 18598 32177 18694 32235
rect 18598 32143 18629 32177
rect 18663 32143 18694 32177
rect 18598 32085 18694 32143
rect 18598 32051 18629 32085
rect 18663 32051 18694 32085
rect 18598 31993 18694 32051
rect 18823 32632 18885 32647
rect 18823 32598 18836 32632
rect 18870 32598 18885 32632
rect 18823 32065 18885 32598
rect 19054 32392 19094 33032
rect 19142 32729 19238 32758
rect 19142 32695 19173 32729
rect 19207 32695 19238 32729
rect 19142 32637 19238 32695
rect 19142 32603 19173 32637
rect 19207 32603 19238 32637
rect 19142 32545 19238 32603
rect 19142 32511 19173 32545
rect 19207 32511 19238 32545
rect 19142 32453 19238 32511
rect 19142 32419 19173 32453
rect 19207 32419 19238 32453
rect 19050 32352 19106 32392
rect 19050 32318 19058 32352
rect 19092 32318 19106 32352
rect 19050 32296 19106 32318
rect 19142 32361 19238 32419
rect 19142 32327 19173 32361
rect 19207 32327 19238 32361
rect 19142 32269 19238 32327
rect 19142 32235 19173 32269
rect 19207 32235 19238 32269
rect 19142 32177 19238 32235
rect 19142 32143 19173 32177
rect 19207 32143 19238 32177
rect 19142 32085 19238 32143
rect 18823 32003 19032 32065
rect 18598 31959 18629 31993
rect 18663 31959 18694 31993
rect 18598 31901 18694 31959
rect 18598 31867 18629 31901
rect 18663 31867 18694 31901
rect 18598 31850 18694 31867
rect 18861 31899 18907 31911
rect 18861 31865 18867 31899
rect 18901 31865 18907 31899
rect 18861 31853 18907 31865
rect 18598 31784 18618 31850
rect 18684 31784 18694 31850
rect 18598 31775 18629 31784
rect 18663 31775 18694 31784
rect 18598 31717 18694 31775
rect 18793 31812 18839 31824
rect 18793 31778 18799 31812
rect 18833 31778 18839 31812
rect 18793 31766 18839 31778
rect 18598 31683 18629 31717
rect 18663 31683 18694 31717
rect 18598 31625 18694 31683
rect 18598 31591 18629 31625
rect 18663 31591 18694 31625
rect 18598 31533 18694 31591
rect 18598 31499 18629 31533
rect 18663 31499 18694 31533
rect 18802 31510 18830 31766
rect 18598 31441 18694 31499
rect 18793 31498 18839 31510
rect 18793 31464 18799 31498
rect 18833 31464 18839 31498
rect 18793 31452 18839 31464
rect 18598 31407 18629 31441
rect 18663 31407 18694 31441
rect 18598 31349 18694 31407
rect 18598 31315 18629 31349
rect 18663 31315 18694 31349
rect 18598 31257 18694 31315
rect 18598 31223 18629 31257
rect 18663 31223 18694 31257
rect 18598 31165 18694 31223
rect 18598 31131 18629 31165
rect 18663 31131 18694 31165
rect 18598 31073 18694 31131
rect 18802 31090 18830 31452
rect 18870 31407 18898 31853
rect 18861 31395 18907 31407
rect 18861 31361 18867 31395
rect 18901 31361 18907 31395
rect 18861 31349 18907 31361
rect 18870 31169 18898 31349
rect 18970 31304 19032 32003
rect 19142 32051 19173 32085
rect 19207 32051 19238 32085
rect 19142 31993 19238 32051
rect 19142 31959 19173 31993
rect 19207 31959 19238 31993
rect 19142 31901 19238 31959
rect 19142 31867 19173 31901
rect 19207 31867 19238 31901
rect 19142 31860 19238 31867
rect 19142 31794 19160 31860
rect 19226 31794 19238 31860
rect 19142 31775 19173 31794
rect 19207 31775 19238 31794
rect 19142 31717 19238 31775
rect 19142 31683 19173 31717
rect 19207 31683 19238 31717
rect 19142 31625 19238 31683
rect 19142 31591 19173 31625
rect 19207 31591 19238 31625
rect 19142 31533 19238 31591
rect 19142 31499 19173 31533
rect 19207 31499 19238 31533
rect 19142 31441 19238 31499
rect 19142 31407 19173 31441
rect 19207 31407 19238 31441
rect 19142 31349 19238 31407
rect 19142 31315 19173 31349
rect 19207 31315 19238 31349
rect 18970 31242 19046 31304
rect 18970 31202 18988 31242
rect 19028 31202 19046 31242
rect 18970 31184 19046 31202
rect 19142 31257 19238 31315
rect 19142 31223 19173 31257
rect 19207 31223 19238 31257
rect 18861 31157 18907 31169
rect 18861 31123 18867 31157
rect 18901 31123 18907 31157
rect 18861 31111 18907 31123
rect 19142 31165 19238 31223
rect 19142 31131 19173 31165
rect 19207 31131 19238 31165
rect 18598 31039 18629 31073
rect 18663 31039 18694 31073
rect 18598 30981 18694 31039
rect 18793 31078 18839 31090
rect 18793 31044 18799 31078
rect 18833 31044 18839 31078
rect 18793 31032 18839 31044
rect 19142 31073 19238 31131
rect 19142 31039 19173 31073
rect 19207 31039 19238 31073
rect 18598 30947 18629 30981
rect 18663 30947 18694 30981
rect 18598 30918 18694 30947
rect 18879 30984 19025 31011
rect 18879 30950 18940 30984
rect 18976 30950 19025 30984
rect 18879 30780 19025 30950
rect 19142 30981 19238 31039
rect 19142 30947 19173 30981
rect 19207 30947 19238 30981
rect 19142 30918 19238 30947
rect 18879 30740 19098 30780
rect 18602 30483 18698 30512
rect 18602 30449 18633 30483
rect 18667 30449 18698 30483
rect 18602 30391 18698 30449
rect 18602 30357 18633 30391
rect 18667 30357 18698 30391
rect 18602 30299 18698 30357
rect 18602 30265 18633 30299
rect 18667 30265 18698 30299
rect 18602 30207 18698 30265
rect 18602 30173 18633 30207
rect 18667 30173 18698 30207
rect 18602 30115 18698 30173
rect 18602 30081 18633 30115
rect 18667 30081 18698 30115
rect 18602 30023 18698 30081
rect 18602 29989 18633 30023
rect 18667 29989 18698 30023
rect 18602 29931 18698 29989
rect 18602 29897 18633 29931
rect 18667 29897 18698 29931
rect 18602 29839 18698 29897
rect 18602 29805 18633 29839
rect 18667 29805 18698 29839
rect 18602 29747 18698 29805
rect 18827 30386 18889 30401
rect 18827 30352 18840 30386
rect 18874 30352 18889 30386
rect 18827 29819 18889 30352
rect 19058 30146 19098 30740
rect 19146 30483 19242 30512
rect 19146 30449 19177 30483
rect 19211 30449 19242 30483
rect 19146 30391 19242 30449
rect 19146 30357 19177 30391
rect 19211 30357 19242 30391
rect 19146 30299 19242 30357
rect 19146 30265 19177 30299
rect 19211 30265 19242 30299
rect 19146 30207 19242 30265
rect 19146 30173 19177 30207
rect 19211 30173 19242 30207
rect 19054 30106 19110 30146
rect 19054 30072 19062 30106
rect 19096 30072 19110 30106
rect 19054 30050 19110 30072
rect 19146 30115 19242 30173
rect 19146 30081 19177 30115
rect 19211 30081 19242 30115
rect 19146 30023 19242 30081
rect 19146 29989 19177 30023
rect 19211 29989 19242 30023
rect 19146 29931 19242 29989
rect 19146 29897 19177 29931
rect 19211 29897 19242 29931
rect 19146 29839 19242 29897
rect 18827 29757 19036 29819
rect 18602 29713 18633 29747
rect 18667 29713 18698 29747
rect 18602 29655 18698 29713
rect 18602 29621 18633 29655
rect 18667 29621 18698 29655
rect 18602 29604 18698 29621
rect 18865 29653 18911 29665
rect 18865 29619 18871 29653
rect 18905 29619 18911 29653
rect 18865 29607 18911 29619
rect 18602 29538 18622 29604
rect 18688 29538 18698 29604
rect 18602 29529 18633 29538
rect 18667 29529 18698 29538
rect 18602 29471 18698 29529
rect 18797 29566 18843 29578
rect 18797 29532 18803 29566
rect 18837 29532 18843 29566
rect 18797 29520 18843 29532
rect 18602 29437 18633 29471
rect 18667 29437 18698 29471
rect 18602 29379 18698 29437
rect 18602 29345 18633 29379
rect 18667 29345 18698 29379
rect 18602 29287 18698 29345
rect 18602 29253 18633 29287
rect 18667 29253 18698 29287
rect 18806 29264 18834 29520
rect 18602 29195 18698 29253
rect 18797 29252 18843 29264
rect 18797 29218 18803 29252
rect 18837 29218 18843 29252
rect 18797 29206 18843 29218
rect 18602 29161 18633 29195
rect 18667 29161 18698 29195
rect 18602 29103 18698 29161
rect 18602 29069 18633 29103
rect 18667 29069 18698 29103
rect 18602 29011 18698 29069
rect 18602 28977 18633 29011
rect 18667 28977 18698 29011
rect 18602 28919 18698 28977
rect 18602 28885 18633 28919
rect 18667 28885 18698 28919
rect 18602 28827 18698 28885
rect 18806 28844 18834 29206
rect 18874 29161 18902 29607
rect 18865 29149 18911 29161
rect 18865 29115 18871 29149
rect 18905 29115 18911 29149
rect 18865 29103 18911 29115
rect 18874 28923 18902 29103
rect 18974 29058 19036 29757
rect 19146 29805 19177 29839
rect 19211 29805 19242 29839
rect 19146 29747 19242 29805
rect 19146 29713 19177 29747
rect 19211 29713 19242 29747
rect 19146 29655 19242 29713
rect 19146 29621 19177 29655
rect 19211 29621 19242 29655
rect 19146 29614 19242 29621
rect 19146 29548 19164 29614
rect 19230 29548 19242 29614
rect 19146 29529 19177 29548
rect 19211 29529 19242 29548
rect 19146 29471 19242 29529
rect 19146 29437 19177 29471
rect 19211 29437 19242 29471
rect 19146 29379 19242 29437
rect 19146 29345 19177 29379
rect 19211 29345 19242 29379
rect 19146 29287 19242 29345
rect 19146 29253 19177 29287
rect 19211 29253 19242 29287
rect 19146 29195 19242 29253
rect 19146 29161 19177 29195
rect 19211 29161 19242 29195
rect 19146 29103 19242 29161
rect 19146 29069 19177 29103
rect 19211 29069 19242 29103
rect 18974 28996 19050 29058
rect 18974 28956 18992 28996
rect 19032 28956 19050 28996
rect 18974 28938 19050 28956
rect 19146 29011 19242 29069
rect 19146 28977 19177 29011
rect 19211 28977 19242 29011
rect 18865 28911 18911 28923
rect 18865 28877 18871 28911
rect 18905 28877 18911 28911
rect 18865 28865 18911 28877
rect 19146 28919 19242 28977
rect 19146 28885 19177 28919
rect 19211 28885 19242 28919
rect 18602 28793 18633 28827
rect 18667 28793 18698 28827
rect 18602 28735 18698 28793
rect 18797 28832 18843 28844
rect 18797 28798 18803 28832
rect 18837 28798 18843 28832
rect 18797 28786 18843 28798
rect 19146 28827 19242 28885
rect 19146 28793 19177 28827
rect 19211 28793 19242 28827
rect 18602 28701 18633 28735
rect 18667 28701 18698 28735
rect 18602 28672 18698 28701
rect 18883 28738 19029 28765
rect 18883 28704 18944 28738
rect 18980 28704 19029 28738
rect 18883 28558 19029 28704
rect 19146 28735 19242 28793
rect 19146 28701 19177 28735
rect 19211 28701 19242 28735
rect 19146 28672 19242 28701
rect 18883 28514 19090 28558
rect 18594 28297 18690 28326
rect 18594 28263 18625 28297
rect 18659 28263 18690 28297
rect 18594 28205 18690 28263
rect 18594 28171 18625 28205
rect 18659 28171 18690 28205
rect 18594 28113 18690 28171
rect 18594 28079 18625 28113
rect 18659 28079 18690 28113
rect 18594 28021 18690 28079
rect 18594 27987 18625 28021
rect 18659 27987 18690 28021
rect 18594 27929 18690 27987
rect 18594 27895 18625 27929
rect 18659 27895 18690 27929
rect 18594 27837 18690 27895
rect 18594 27803 18625 27837
rect 18659 27803 18690 27837
rect 18594 27745 18690 27803
rect 18594 27711 18625 27745
rect 18659 27711 18690 27745
rect 18594 27653 18690 27711
rect 18594 27619 18625 27653
rect 18659 27619 18690 27653
rect 18594 27561 18690 27619
rect 18819 28200 18881 28215
rect 18819 28166 18832 28200
rect 18866 28166 18881 28200
rect 18819 27633 18881 28166
rect 19050 27960 19090 28514
rect 19138 28297 19234 28326
rect 19138 28263 19169 28297
rect 19203 28263 19234 28297
rect 19138 28205 19234 28263
rect 19138 28171 19169 28205
rect 19203 28171 19234 28205
rect 19138 28113 19234 28171
rect 19138 28079 19169 28113
rect 19203 28079 19234 28113
rect 19138 28021 19234 28079
rect 19138 27987 19169 28021
rect 19203 27987 19234 28021
rect 19046 27920 19102 27960
rect 19046 27886 19054 27920
rect 19088 27886 19102 27920
rect 19046 27864 19102 27886
rect 19138 27929 19234 27987
rect 19138 27895 19169 27929
rect 19203 27895 19234 27929
rect 19138 27837 19234 27895
rect 19138 27803 19169 27837
rect 19203 27803 19234 27837
rect 19138 27745 19234 27803
rect 19138 27711 19169 27745
rect 19203 27711 19234 27745
rect 19138 27653 19234 27711
rect 18819 27571 19028 27633
rect 18594 27527 18625 27561
rect 18659 27527 18690 27561
rect 18594 27469 18690 27527
rect 18594 27435 18625 27469
rect 18659 27435 18690 27469
rect 18594 27418 18690 27435
rect 18857 27467 18903 27479
rect 18857 27433 18863 27467
rect 18897 27433 18903 27467
rect 18857 27421 18903 27433
rect 18594 27352 18614 27418
rect 18680 27352 18690 27418
rect 18594 27343 18625 27352
rect 18659 27343 18690 27352
rect 18594 27285 18690 27343
rect 18789 27380 18835 27392
rect 18789 27346 18795 27380
rect 18829 27346 18835 27380
rect 18789 27334 18835 27346
rect 18594 27251 18625 27285
rect 18659 27251 18690 27285
rect 18594 27193 18690 27251
rect 18594 27159 18625 27193
rect 18659 27159 18690 27193
rect 18594 27101 18690 27159
rect 18594 27067 18625 27101
rect 18659 27067 18690 27101
rect 18798 27078 18826 27334
rect 18594 27009 18690 27067
rect 18789 27066 18835 27078
rect 18789 27032 18795 27066
rect 18829 27032 18835 27066
rect 18789 27020 18835 27032
rect 18594 26975 18625 27009
rect 18659 26975 18690 27009
rect 18594 26917 18690 26975
rect 18594 26883 18625 26917
rect 18659 26883 18690 26917
rect 18594 26825 18690 26883
rect 18594 26791 18625 26825
rect 18659 26791 18690 26825
rect 18594 26733 18690 26791
rect 18594 26699 18625 26733
rect 18659 26699 18690 26733
rect 18594 26641 18690 26699
rect 18798 26658 18826 27020
rect 18866 26975 18894 27421
rect 18857 26963 18903 26975
rect 18857 26929 18863 26963
rect 18897 26929 18903 26963
rect 18857 26917 18903 26929
rect 18866 26737 18894 26917
rect 18966 26872 19028 27571
rect 19138 27619 19169 27653
rect 19203 27619 19234 27653
rect 19138 27561 19234 27619
rect 19138 27527 19169 27561
rect 19203 27527 19234 27561
rect 19138 27469 19234 27527
rect 19138 27435 19169 27469
rect 19203 27435 19234 27469
rect 19138 27428 19234 27435
rect 19138 27362 19156 27428
rect 19222 27362 19234 27428
rect 19138 27343 19169 27362
rect 19203 27343 19234 27362
rect 19138 27285 19234 27343
rect 19138 27251 19169 27285
rect 19203 27251 19234 27285
rect 19138 27193 19234 27251
rect 19138 27159 19169 27193
rect 19203 27159 19234 27193
rect 19138 27101 19234 27159
rect 19138 27067 19169 27101
rect 19203 27067 19234 27101
rect 19138 27009 19234 27067
rect 19138 26975 19169 27009
rect 19203 26975 19234 27009
rect 19138 26917 19234 26975
rect 19138 26883 19169 26917
rect 19203 26883 19234 26917
rect 18966 26810 19042 26872
rect 18966 26770 18984 26810
rect 19024 26770 19042 26810
rect 18966 26752 19042 26770
rect 19138 26825 19234 26883
rect 19138 26791 19169 26825
rect 19203 26791 19234 26825
rect 18857 26725 18903 26737
rect 18857 26691 18863 26725
rect 18897 26691 18903 26725
rect 18857 26679 18903 26691
rect 19138 26733 19234 26791
rect 19138 26699 19169 26733
rect 19203 26699 19234 26733
rect 18594 26607 18625 26641
rect 18659 26607 18690 26641
rect 18594 26549 18690 26607
rect 18789 26646 18835 26658
rect 18789 26612 18795 26646
rect 18829 26612 18835 26646
rect 18789 26600 18835 26612
rect 19138 26641 19234 26699
rect 19138 26607 19169 26641
rect 19203 26607 19234 26641
rect 18594 26515 18625 26549
rect 18659 26515 18690 26549
rect 18594 26486 18690 26515
rect 18875 26552 19021 26579
rect 18875 26518 18936 26552
rect 18972 26518 19021 26552
rect 18875 26348 19021 26518
rect 19138 26549 19234 26607
rect 19138 26515 19169 26549
rect 19203 26515 19234 26549
rect 19138 26486 19234 26515
rect 18875 26308 19094 26348
rect 18598 26051 18694 26080
rect 18598 26017 18629 26051
rect 18663 26017 18694 26051
rect 18598 25959 18694 26017
rect 18598 25925 18629 25959
rect 18663 25925 18694 25959
rect 18598 25867 18694 25925
rect 18598 25833 18629 25867
rect 18663 25833 18694 25867
rect 18598 25775 18694 25833
rect 18598 25741 18629 25775
rect 18663 25741 18694 25775
rect 18598 25683 18694 25741
rect 18598 25649 18629 25683
rect 18663 25649 18694 25683
rect 18598 25591 18694 25649
rect 18598 25557 18629 25591
rect 18663 25557 18694 25591
rect 18598 25499 18694 25557
rect 18598 25465 18629 25499
rect 18663 25465 18694 25499
rect 18598 25407 18694 25465
rect 18598 25373 18629 25407
rect 18663 25373 18694 25407
rect 18598 25315 18694 25373
rect 18823 25954 18885 25969
rect 18823 25920 18836 25954
rect 18870 25920 18885 25954
rect 18823 25387 18885 25920
rect 19054 25714 19094 26308
rect 19142 26051 19238 26080
rect 19142 26017 19173 26051
rect 19207 26017 19238 26051
rect 19142 25959 19238 26017
rect 19142 25925 19173 25959
rect 19207 25925 19238 25959
rect 19142 25867 19238 25925
rect 19142 25833 19173 25867
rect 19207 25833 19238 25867
rect 19142 25775 19238 25833
rect 19142 25741 19173 25775
rect 19207 25741 19238 25775
rect 19050 25674 19106 25714
rect 19050 25640 19058 25674
rect 19092 25640 19106 25674
rect 19050 25618 19106 25640
rect 19142 25683 19238 25741
rect 19142 25649 19173 25683
rect 19207 25649 19238 25683
rect 19142 25591 19238 25649
rect 19142 25557 19173 25591
rect 19207 25557 19238 25591
rect 19142 25499 19238 25557
rect 19142 25465 19173 25499
rect 19207 25465 19238 25499
rect 19142 25407 19238 25465
rect 18823 25325 19032 25387
rect 18598 25281 18629 25315
rect 18663 25281 18694 25315
rect 18598 25223 18694 25281
rect 18598 25189 18629 25223
rect 18663 25189 18694 25223
rect 18598 25172 18694 25189
rect 18861 25221 18907 25233
rect 18861 25187 18867 25221
rect 18901 25187 18907 25221
rect 18861 25175 18907 25187
rect 18598 25106 18618 25172
rect 18684 25106 18694 25172
rect 18598 25097 18629 25106
rect 18663 25097 18694 25106
rect 18598 25039 18694 25097
rect 18793 25134 18839 25146
rect 18793 25100 18799 25134
rect 18833 25100 18839 25134
rect 18793 25088 18839 25100
rect 18598 25005 18629 25039
rect 18663 25005 18694 25039
rect 18598 24947 18694 25005
rect 18598 24913 18629 24947
rect 18663 24913 18694 24947
rect 18598 24855 18694 24913
rect 18598 24821 18629 24855
rect 18663 24821 18694 24855
rect 18802 24832 18830 25088
rect 18598 24763 18694 24821
rect 18793 24820 18839 24832
rect 18793 24786 18799 24820
rect 18833 24786 18839 24820
rect 18793 24774 18839 24786
rect 18598 24729 18629 24763
rect 18663 24729 18694 24763
rect 18598 24671 18694 24729
rect 18598 24637 18629 24671
rect 18663 24637 18694 24671
rect 18598 24579 18694 24637
rect 18598 24545 18629 24579
rect 18663 24545 18694 24579
rect 18598 24487 18694 24545
rect 18598 24453 18629 24487
rect 18663 24453 18694 24487
rect 18598 24395 18694 24453
rect 18802 24412 18830 24774
rect 18870 24729 18898 25175
rect 18861 24717 18907 24729
rect 18861 24683 18867 24717
rect 18901 24683 18907 24717
rect 18861 24671 18907 24683
rect 18870 24491 18898 24671
rect 18970 24626 19032 25325
rect 19142 25373 19173 25407
rect 19207 25373 19238 25407
rect 19142 25315 19238 25373
rect 19142 25281 19173 25315
rect 19207 25281 19238 25315
rect 19142 25223 19238 25281
rect 19142 25189 19173 25223
rect 19207 25189 19238 25223
rect 19142 25182 19238 25189
rect 19142 25116 19160 25182
rect 19226 25116 19238 25182
rect 19142 25097 19173 25116
rect 19207 25097 19238 25116
rect 19142 25039 19238 25097
rect 19142 25005 19173 25039
rect 19207 25005 19238 25039
rect 19142 24947 19238 25005
rect 19142 24913 19173 24947
rect 19207 24913 19238 24947
rect 19142 24855 19238 24913
rect 19142 24821 19173 24855
rect 19207 24821 19238 24855
rect 19142 24763 19238 24821
rect 19142 24729 19173 24763
rect 19207 24729 19238 24763
rect 19142 24671 19238 24729
rect 19142 24637 19173 24671
rect 19207 24637 19238 24671
rect 18970 24564 19046 24626
rect 18970 24524 18988 24564
rect 19028 24524 19046 24564
rect 18970 24506 19046 24524
rect 19142 24579 19238 24637
rect 19142 24545 19173 24579
rect 19207 24545 19238 24579
rect 18861 24479 18907 24491
rect 18861 24445 18867 24479
rect 18901 24445 18907 24479
rect 18861 24433 18907 24445
rect 19142 24487 19238 24545
rect 19142 24453 19173 24487
rect 19207 24453 19238 24487
rect 18598 24361 18629 24395
rect 18663 24361 18694 24395
rect 18598 24303 18694 24361
rect 18793 24400 18839 24412
rect 18793 24366 18799 24400
rect 18833 24366 18839 24400
rect 18793 24354 18839 24366
rect 19142 24395 19238 24453
rect 19142 24361 19173 24395
rect 19207 24361 19238 24395
rect 18598 24269 18629 24303
rect 18663 24269 18694 24303
rect 18598 24240 18694 24269
rect 18879 24306 19025 24333
rect 18879 24272 18940 24306
rect 18976 24272 19025 24306
rect 18879 23936 19025 24272
rect 19142 24303 19238 24361
rect 19142 24269 19173 24303
rect 19207 24269 19238 24303
rect 19142 24240 19238 24269
rect 7670 23400 9510 23420
rect 7670 23389 8536 23400
rect 8602 23389 9510 23400
rect 7670 23355 7699 23389
rect 7733 23355 7791 23389
rect 7825 23355 7883 23389
rect 7917 23355 7975 23389
rect 8009 23355 8067 23389
rect 8101 23355 8159 23389
rect 8193 23355 8251 23389
rect 8285 23355 8343 23389
rect 8377 23355 8435 23389
rect 8469 23355 8527 23389
rect 8602 23355 8619 23389
rect 8653 23355 8711 23389
rect 8745 23355 8803 23389
rect 8837 23355 8895 23389
rect 8929 23355 8987 23389
rect 9021 23355 9079 23389
rect 9113 23355 9171 23389
rect 9205 23355 9263 23389
rect 9297 23355 9355 23389
rect 9389 23355 9447 23389
rect 9481 23355 9510 23389
rect 7670 23334 8536 23355
rect 8602 23334 9510 23355
rect 7670 23324 9510 23334
rect 9916 23404 11756 23424
rect 9916 23393 10782 23404
rect 10848 23393 11756 23404
rect 9916 23359 9945 23393
rect 9979 23359 10037 23393
rect 10071 23359 10129 23393
rect 10163 23359 10221 23393
rect 10255 23359 10313 23393
rect 10347 23359 10405 23393
rect 10439 23359 10497 23393
rect 10531 23359 10589 23393
rect 10623 23359 10681 23393
rect 10715 23359 10773 23393
rect 10848 23359 10865 23393
rect 10899 23359 10957 23393
rect 10991 23359 11049 23393
rect 11083 23359 11141 23393
rect 11175 23359 11233 23393
rect 11267 23359 11325 23393
rect 11359 23359 11417 23393
rect 11451 23359 11509 23393
rect 11543 23359 11601 23393
rect 11635 23359 11693 23393
rect 11727 23359 11756 23393
rect 9916 23338 10782 23359
rect 10848 23338 11756 23359
rect 9916 23328 11756 23338
rect 12102 23396 13942 23416
rect 12102 23385 12968 23396
rect 13034 23385 13942 23396
rect 12102 23351 12131 23385
rect 12165 23351 12223 23385
rect 12257 23351 12315 23385
rect 12349 23351 12407 23385
rect 12441 23351 12499 23385
rect 12533 23351 12591 23385
rect 12625 23351 12683 23385
rect 12717 23351 12775 23385
rect 12809 23351 12867 23385
rect 12901 23351 12959 23385
rect 13034 23351 13051 23385
rect 13085 23351 13143 23385
rect 13177 23351 13235 23385
rect 13269 23351 13327 23385
rect 13361 23351 13419 23385
rect 13453 23351 13511 23385
rect 13545 23351 13603 23385
rect 13637 23351 13695 23385
rect 13729 23351 13787 23385
rect 13821 23351 13879 23385
rect 13913 23351 13942 23385
rect 12102 23330 12968 23351
rect 13034 23330 13942 23351
rect 12102 23320 13942 23330
rect 14348 23400 16188 23420
rect 14348 23389 15214 23400
rect 15280 23389 16188 23400
rect 14348 23355 14377 23389
rect 14411 23355 14469 23389
rect 14503 23355 14561 23389
rect 14595 23355 14653 23389
rect 14687 23355 14745 23389
rect 14779 23355 14837 23389
rect 14871 23355 14929 23389
rect 14963 23355 15021 23389
rect 15055 23355 15113 23389
rect 15147 23355 15205 23389
rect 15280 23355 15297 23389
rect 15331 23355 15389 23389
rect 15423 23355 15481 23389
rect 15515 23355 15573 23389
rect 15607 23355 15665 23389
rect 15699 23355 15757 23389
rect 15791 23355 15849 23389
rect 15883 23355 15941 23389
rect 15975 23355 16033 23389
rect 16067 23355 16125 23389
rect 16159 23355 16188 23389
rect 14348 23334 15214 23355
rect 15280 23334 16188 23355
rect 14348 23324 16188 23334
rect 16630 23400 18470 23420
rect 16630 23389 17496 23400
rect 17562 23389 18470 23400
rect 16630 23355 16659 23389
rect 16693 23355 16751 23389
rect 16785 23355 16843 23389
rect 16877 23355 16935 23389
rect 16969 23355 17027 23389
rect 17061 23355 17119 23389
rect 17153 23355 17211 23389
rect 17245 23355 17303 23389
rect 17337 23355 17395 23389
rect 17429 23355 17487 23389
rect 17562 23355 17579 23389
rect 17613 23355 17671 23389
rect 17705 23355 17763 23389
rect 17797 23355 17855 23389
rect 17889 23355 17947 23389
rect 17981 23355 18039 23389
rect 18073 23355 18131 23389
rect 18165 23355 18223 23389
rect 18257 23355 18315 23389
rect 18349 23355 18407 23389
rect 18441 23355 18470 23389
rect 16630 23334 17496 23355
rect 17562 23334 18470 23355
rect 16630 23324 18470 23334
rect 7784 23219 7842 23225
rect 7784 23185 7796 23219
rect 7830 23216 7842 23219
rect 8204 23219 8262 23225
rect 8204 23216 8216 23219
rect 7830 23188 8216 23216
rect 7830 23185 7842 23188
rect 7784 23179 7842 23185
rect 8204 23185 8216 23188
rect 8250 23216 8262 23219
rect 8518 23219 8576 23225
rect 8518 23216 8530 23219
rect 8250 23188 8530 23216
rect 8250 23185 8262 23188
rect 8204 23179 8262 23185
rect 8518 23185 8530 23188
rect 8564 23185 8576 23219
rect 10030 23223 10088 23229
rect 8518 23179 8576 23185
rect 8755 23182 9399 23195
rect 10030 23189 10042 23223
rect 10076 23220 10088 23223
rect 10450 23223 10508 23229
rect 10450 23220 10462 23223
rect 10076 23192 10462 23220
rect 10076 23189 10088 23192
rect 10030 23183 10088 23189
rect 10450 23189 10462 23192
rect 10496 23220 10508 23223
rect 10764 23223 10822 23229
rect 10764 23220 10776 23223
rect 10496 23192 10776 23220
rect 10496 23189 10508 23192
rect 10450 23183 10508 23189
rect 10764 23189 10776 23192
rect 10810 23189 10822 23223
rect 12216 23215 12274 23221
rect 10764 23183 10822 23189
rect 11001 23186 11645 23199
rect 7863 23151 7921 23157
rect 6269 23078 7763 23139
rect 7863 23117 7875 23151
rect 7909 23148 7921 23151
rect 8101 23151 8159 23157
rect 8101 23148 8113 23151
rect 7909 23120 8113 23148
rect 7909 23117 7921 23120
rect 7863 23111 7921 23117
rect 8101 23117 8113 23120
rect 8147 23148 8159 23151
rect 8605 23151 8663 23157
rect 8605 23148 8617 23151
rect 8147 23120 8617 23148
rect 8147 23117 8159 23120
rect 8101 23111 8159 23117
rect 8605 23117 8617 23120
rect 8651 23117 8663 23151
rect 8605 23111 8663 23117
rect 8755 23148 9350 23182
rect 9384 23148 9399 23182
rect 8755 23133 9399 23148
rect 10109 23155 10167 23161
rect 6269 23042 7702 23078
rect 7736 23042 7763 23078
rect 8755 23048 8817 23133
rect 6269 22993 7763 23042
rect 7936 23030 8817 23048
rect 6269 18485 6415 22993
rect 7936 22990 7954 23030
rect 7994 22990 8817 23030
rect 7936 22986 8817 22990
rect 9738 23082 10009 23143
rect 10109 23121 10121 23155
rect 10155 23152 10167 23155
rect 10347 23155 10405 23161
rect 10347 23152 10359 23155
rect 10155 23124 10359 23152
rect 10155 23121 10167 23124
rect 10109 23115 10167 23121
rect 10347 23121 10359 23124
rect 10393 23152 10405 23155
rect 10851 23155 10909 23161
rect 10851 23152 10863 23155
rect 10393 23124 10863 23152
rect 10393 23121 10405 23124
rect 10347 23115 10405 23121
rect 10851 23121 10863 23124
rect 10897 23121 10909 23155
rect 10851 23115 10909 23121
rect 11001 23152 11596 23186
rect 11630 23152 11645 23186
rect 12216 23181 12228 23215
rect 12262 23212 12274 23215
rect 12636 23215 12694 23221
rect 12636 23212 12648 23215
rect 12262 23184 12648 23212
rect 12262 23181 12274 23184
rect 12216 23175 12274 23181
rect 12636 23181 12648 23184
rect 12682 23212 12694 23215
rect 12950 23215 13008 23221
rect 12950 23212 12962 23215
rect 12682 23184 12962 23212
rect 12682 23181 12694 23184
rect 12636 23175 12694 23181
rect 12950 23181 12962 23184
rect 12996 23181 13008 23215
rect 14462 23219 14520 23225
rect 12950 23175 13008 23181
rect 13187 23178 13831 23191
rect 14462 23185 14474 23219
rect 14508 23216 14520 23219
rect 14882 23219 14940 23225
rect 14882 23216 14894 23219
rect 14508 23188 14894 23216
rect 14508 23185 14520 23188
rect 14462 23179 14520 23185
rect 14882 23185 14894 23188
rect 14928 23216 14940 23219
rect 15196 23219 15254 23225
rect 15196 23216 15208 23219
rect 14928 23188 15208 23216
rect 14928 23185 14940 23188
rect 14882 23179 14940 23185
rect 15196 23185 15208 23188
rect 15242 23185 15254 23219
rect 16744 23219 16802 23225
rect 15196 23179 15254 23185
rect 15433 23182 16077 23195
rect 11001 23137 11645 23152
rect 12295 23147 12353 23153
rect 9738 23046 9948 23082
rect 9982 23046 10009 23082
rect 11001 23052 11063 23137
rect 9738 22997 10009 23046
rect 10182 23034 11063 23052
rect 7936 22972 8056 22986
rect 9048 22964 9144 22968
rect 9738 22964 9778 22997
rect 10182 22994 10200 23034
rect 10240 22994 11063 23034
rect 10182 22990 11063 22994
rect 11944 23074 12195 23135
rect 12295 23113 12307 23147
rect 12341 23144 12353 23147
rect 12533 23147 12591 23153
rect 12533 23144 12545 23147
rect 12341 23116 12545 23144
rect 12341 23113 12353 23116
rect 12295 23107 12353 23113
rect 12533 23113 12545 23116
rect 12579 23144 12591 23147
rect 13037 23147 13095 23153
rect 13037 23144 13049 23147
rect 12579 23116 13049 23144
rect 12579 23113 12591 23116
rect 12533 23107 12591 23113
rect 13037 23113 13049 23116
rect 13083 23113 13095 23147
rect 13037 23107 13095 23113
rect 13187 23144 13782 23178
rect 13816 23144 13831 23178
rect 13187 23129 13831 23144
rect 14541 23151 14599 23157
rect 11944 23038 12134 23074
rect 12168 23038 12195 23074
rect 13187 23044 13249 23129
rect 10182 22976 10302 22990
rect 11944 22989 12195 23038
rect 12368 23026 13249 23044
rect 9048 22960 9778 22964
rect 9048 22926 9070 22960
rect 9104 22926 9778 22960
rect 9048 22924 9778 22926
rect 11294 22968 11390 22972
rect 11944 22968 11988 22989
rect 12368 22986 12386 23026
rect 12426 22986 13249 23026
rect 12368 22982 13249 22986
rect 14170 23078 14441 23139
rect 14541 23117 14553 23151
rect 14587 23148 14599 23151
rect 14779 23151 14837 23157
rect 14779 23148 14791 23151
rect 14587 23120 14791 23148
rect 14587 23117 14599 23120
rect 14541 23111 14599 23117
rect 14779 23117 14791 23120
rect 14825 23148 14837 23151
rect 15283 23151 15341 23157
rect 15283 23148 15295 23151
rect 14825 23120 15295 23148
rect 14825 23117 14837 23120
rect 14779 23111 14837 23117
rect 15283 23117 15295 23120
rect 15329 23117 15341 23151
rect 15283 23111 15341 23117
rect 15433 23148 16028 23182
rect 16062 23148 16077 23182
rect 16744 23185 16756 23219
rect 16790 23216 16802 23219
rect 17164 23219 17222 23225
rect 17164 23216 17176 23219
rect 16790 23188 17176 23216
rect 16790 23185 16802 23188
rect 16744 23179 16802 23185
rect 17164 23185 17176 23188
rect 17210 23216 17222 23219
rect 17478 23219 17536 23225
rect 17478 23216 17490 23219
rect 17210 23188 17490 23216
rect 17210 23185 17222 23188
rect 17164 23179 17222 23185
rect 17478 23185 17490 23188
rect 17524 23185 17536 23219
rect 17478 23179 17536 23185
rect 17715 23182 18359 23195
rect 15433 23133 16077 23148
rect 16823 23151 16881 23157
rect 14170 23042 14380 23078
rect 14414 23042 14441 23078
rect 15433 23048 15495 23133
rect 14170 22993 14441 23042
rect 14614 23030 15495 23048
rect 12368 22968 12488 22982
rect 11294 22964 11988 22968
rect 11294 22930 11316 22964
rect 11350 22930 11988 22964
rect 11294 22928 11988 22930
rect 13480 22960 13576 22964
rect 14170 22960 14210 22993
rect 14614 22990 14632 23030
rect 14672 22990 15495 23030
rect 16472 23078 16723 23139
rect 16823 23117 16835 23151
rect 16869 23148 16881 23151
rect 17061 23151 17119 23157
rect 17061 23148 17073 23151
rect 16869 23120 17073 23148
rect 16869 23117 16881 23120
rect 16823 23111 16881 23117
rect 17061 23117 17073 23120
rect 17107 23148 17119 23151
rect 17565 23151 17623 23157
rect 17565 23148 17577 23151
rect 17107 23120 17577 23148
rect 17107 23117 17119 23120
rect 17061 23111 17119 23117
rect 17565 23117 17577 23120
rect 17611 23117 17623 23151
rect 17565 23111 17623 23117
rect 17715 23148 18310 23182
rect 18344 23148 18359 23182
rect 17715 23133 18359 23148
rect 16472 23042 16662 23078
rect 16696 23042 16723 23078
rect 17715 23048 17777 23133
rect 16472 23024 16723 23042
rect 14614 22986 15495 22990
rect 16462 22993 16723 23024
rect 16896 23030 17777 23048
rect 14614 22972 14734 22986
rect 13480 22956 14210 22960
rect 9048 22912 9144 22924
rect 11294 22916 11390 22928
rect 13480 22922 13502 22956
rect 13536 22922 14210 22956
rect 13480 22920 14210 22922
rect 15726 22964 15822 22968
rect 16462 22964 16500 22993
rect 16896 22990 16914 23030
rect 16954 22990 17777 23030
rect 16896 22986 17777 22990
rect 16896 22972 17016 22986
rect 15726 22960 16500 22964
rect 15726 22926 15748 22960
rect 15782 22926 16500 22960
rect 15726 22924 16500 22926
rect 13480 22908 13576 22920
rect 15726 22912 15822 22924
rect 16462 22916 16500 22924
rect 18008 22964 18104 22968
rect 18922 22964 18962 23936
rect 18008 22960 18962 22964
rect 18008 22926 18030 22960
rect 18064 22926 18962 22960
rect 18008 22924 18962 22926
rect 18008 22912 18104 22924
rect 7670 22858 9510 22876
rect 7670 22845 8546 22858
rect 8612 22845 9510 22858
rect 7670 22811 7699 22845
rect 7733 22811 7791 22845
rect 7825 22811 7883 22845
rect 7917 22811 7975 22845
rect 8009 22811 8067 22845
rect 8101 22811 8159 22845
rect 8193 22811 8251 22845
rect 8285 22811 8343 22845
rect 8377 22811 8435 22845
rect 8469 22811 8527 22845
rect 8612 22811 8619 22845
rect 8653 22811 8711 22845
rect 8745 22811 8803 22845
rect 8837 22811 8895 22845
rect 8929 22811 8987 22845
rect 9021 22811 9079 22845
rect 9113 22811 9171 22845
rect 9205 22811 9263 22845
rect 9297 22811 9355 22845
rect 9389 22811 9447 22845
rect 9481 22811 9510 22845
rect 7670 22792 8546 22811
rect 8612 22792 9510 22811
rect 7670 22780 9510 22792
rect 9916 22862 11756 22880
rect 9916 22849 10792 22862
rect 10858 22849 11756 22862
rect 9916 22815 9945 22849
rect 9979 22815 10037 22849
rect 10071 22815 10129 22849
rect 10163 22815 10221 22849
rect 10255 22815 10313 22849
rect 10347 22815 10405 22849
rect 10439 22815 10497 22849
rect 10531 22815 10589 22849
rect 10623 22815 10681 22849
rect 10715 22815 10773 22849
rect 10858 22815 10865 22849
rect 10899 22815 10957 22849
rect 10991 22815 11049 22849
rect 11083 22815 11141 22849
rect 11175 22815 11233 22849
rect 11267 22815 11325 22849
rect 11359 22815 11417 22849
rect 11451 22815 11509 22849
rect 11543 22815 11601 22849
rect 11635 22815 11693 22849
rect 11727 22815 11756 22849
rect 9916 22796 10792 22815
rect 10858 22796 11756 22815
rect 9916 22784 11756 22796
rect 12102 22854 13942 22872
rect 12102 22841 12978 22854
rect 13044 22841 13942 22854
rect 12102 22807 12131 22841
rect 12165 22807 12223 22841
rect 12257 22807 12315 22841
rect 12349 22807 12407 22841
rect 12441 22807 12499 22841
rect 12533 22807 12591 22841
rect 12625 22807 12683 22841
rect 12717 22807 12775 22841
rect 12809 22807 12867 22841
rect 12901 22807 12959 22841
rect 13044 22807 13051 22841
rect 13085 22807 13143 22841
rect 13177 22807 13235 22841
rect 13269 22807 13327 22841
rect 13361 22807 13419 22841
rect 13453 22807 13511 22841
rect 13545 22807 13603 22841
rect 13637 22807 13695 22841
rect 13729 22807 13787 22841
rect 13821 22807 13879 22841
rect 13913 22807 13942 22841
rect 12102 22788 12978 22807
rect 13044 22788 13942 22807
rect 12102 22776 13942 22788
rect 14348 22858 16188 22876
rect 14348 22845 15224 22858
rect 15290 22845 16188 22858
rect 14348 22811 14377 22845
rect 14411 22811 14469 22845
rect 14503 22811 14561 22845
rect 14595 22811 14653 22845
rect 14687 22811 14745 22845
rect 14779 22811 14837 22845
rect 14871 22811 14929 22845
rect 14963 22811 15021 22845
rect 15055 22811 15113 22845
rect 15147 22811 15205 22845
rect 15290 22811 15297 22845
rect 15331 22811 15389 22845
rect 15423 22811 15481 22845
rect 15515 22811 15573 22845
rect 15607 22811 15665 22845
rect 15699 22811 15757 22845
rect 15791 22811 15849 22845
rect 15883 22811 15941 22845
rect 15975 22811 16033 22845
rect 16067 22811 16125 22845
rect 16159 22811 16188 22845
rect 14348 22792 15224 22811
rect 15290 22792 16188 22811
rect 14348 22780 16188 22792
rect 16630 22858 18470 22876
rect 16630 22845 17506 22858
rect 17572 22845 18470 22858
rect 16630 22811 16659 22845
rect 16693 22811 16751 22845
rect 16785 22811 16843 22845
rect 16877 22811 16935 22845
rect 16969 22811 17027 22845
rect 17061 22811 17119 22845
rect 17153 22811 17211 22845
rect 17245 22811 17303 22845
rect 17337 22811 17395 22845
rect 17429 22811 17487 22845
rect 17572 22811 17579 22845
rect 17613 22811 17671 22845
rect 17705 22811 17763 22845
rect 17797 22811 17855 22845
rect 17889 22811 17947 22845
rect 17981 22811 18039 22845
rect 18073 22811 18131 22845
rect 18165 22811 18223 22845
rect 18257 22811 18315 22845
rect 18349 22811 18407 22845
rect 18441 22811 18470 22845
rect 16630 22792 17506 22811
rect 17572 22792 18470 22811
rect 16630 22780 18470 22792
rect 6269 18339 26063 18485
rect 9430 17822 9782 17842
rect 9430 17811 9540 17822
rect 9600 17811 9782 17822
rect 9430 17777 9459 17811
rect 9493 17777 9540 17811
rect 9600 17777 9643 17811
rect 9677 17777 9719 17811
rect 9753 17777 9782 17811
rect 9430 17762 9540 17777
rect 9600 17762 9782 17777
rect 9430 17746 9782 17762
rect 16267 17714 16621 17732
rect 16267 17701 16455 17714
rect 16523 17701 16621 17714
rect 15481 17674 15843 17694
rect 15481 17663 15683 17674
rect 15751 17663 15843 17674
rect 15481 17629 15510 17663
rect 15544 17629 15596 17663
rect 15630 17629 15683 17663
rect 15751 17629 15780 17663
rect 15814 17629 15843 17663
rect 16267 17667 16296 17701
rect 16330 17667 16374 17701
rect 16408 17667 16455 17701
rect 16523 17667 16558 17701
rect 16592 17667 16621 17701
rect 16267 17652 16455 17667
rect 16523 17652 16621 17667
rect 16267 17636 16621 17652
rect 17133 17714 17495 17734
rect 17133 17703 17335 17714
rect 17403 17703 17495 17714
rect 17133 17669 17162 17703
rect 17196 17669 17248 17703
rect 17282 17669 17335 17703
rect 17403 17669 17432 17703
rect 17466 17669 17495 17703
rect 17911 17704 18263 17724
rect 19027 17708 19385 17726
rect 19027 17706 19219 17708
rect 17911 17698 18121 17704
rect 17133 17652 17335 17669
rect 17403 17652 17495 17669
rect 17133 17638 17495 17652
rect 17909 17693 18121 17698
rect 18189 17693 18263 17704
rect 17909 17659 17940 17693
rect 17974 17659 18016 17693
rect 18050 17659 18108 17693
rect 18189 17659 18200 17693
rect 18234 17659 18263 17693
rect 17909 17642 18121 17659
rect 18189 17642 18263 17659
rect 17909 17632 18263 17642
rect 19025 17695 19219 17706
rect 19287 17695 19385 17708
rect 19025 17661 19056 17695
rect 19090 17661 19138 17695
rect 19172 17661 19219 17695
rect 19287 17661 19322 17695
rect 19356 17661 19385 17695
rect 19025 17646 19219 17661
rect 19287 17646 19385 17661
rect 19025 17640 19385 17646
rect 15481 17612 15683 17629
rect 15751 17612 15843 17629
rect 17911 17628 18263 17632
rect 19027 17630 19385 17640
rect 19893 17708 20259 17728
rect 19893 17697 20099 17708
rect 20167 17697 20259 17708
rect 19893 17663 19922 17697
rect 19956 17663 20012 17697
rect 20046 17663 20099 17697
rect 20167 17663 20196 17697
rect 20230 17663 20259 17697
rect 19893 17646 20099 17663
rect 20167 17646 20259 17663
rect 19893 17632 20259 17646
rect 20663 17698 21027 17718
rect 20663 17687 20885 17698
rect 20953 17687 21027 17698
rect 20663 17653 20692 17687
rect 20726 17653 20780 17687
rect 20814 17653 20872 17687
rect 20953 17653 20964 17687
rect 20998 17653 21027 17687
rect 20663 17636 20885 17653
rect 20953 17636 21027 17653
rect 20663 17622 21027 17636
rect 21365 17698 21733 17716
rect 21365 17685 21475 17698
rect 21543 17685 21733 17698
rect 21365 17651 21394 17685
rect 21428 17651 21475 17685
rect 21543 17651 21578 17685
rect 21612 17651 21670 17685
rect 21704 17651 21733 17685
rect 21365 17636 21475 17651
rect 21543 17636 21733 17651
rect 21365 17620 21733 17636
rect 22149 17698 22515 17718
rect 22149 17687 22355 17698
rect 22423 17687 22515 17698
rect 22149 17653 22178 17687
rect 22212 17653 22268 17687
rect 22302 17653 22355 17687
rect 22423 17653 22452 17687
rect 22486 17653 22515 17687
rect 22149 17636 22355 17653
rect 22423 17636 22515 17653
rect 22149 17622 22515 17636
rect 23007 17688 23373 17708
rect 23007 17677 23141 17688
rect 23209 17677 23373 17688
rect 23007 17643 23036 17677
rect 23070 17643 23128 17677
rect 23209 17643 23220 17677
rect 23254 17643 23310 17677
rect 23344 17643 23373 17677
rect 23007 17626 23141 17643
rect 23209 17626 23373 17643
rect 23007 17612 23373 17626
rect 15481 17598 15843 17612
rect 6603 17576 9539 17587
rect 6603 17504 6646 17576
rect 6722 17568 9539 17576
rect 6722 17532 9496 17568
rect 9532 17532 9539 17568
rect 6722 17504 9539 17532
rect 6603 17497 9539 17504
rect 9573 17572 13733 17587
rect 9573 17536 9596 17572
rect 9632 17536 13733 17572
rect 9573 17497 13733 17536
rect 9430 17286 9782 17298
rect 9430 17278 9796 17286
rect 9430 17267 9536 17278
rect 9594 17267 9796 17278
rect 9430 17233 9459 17267
rect 9493 17233 9536 17267
rect 9594 17233 9643 17267
rect 9677 17233 9719 17267
rect 9753 17233 9796 17267
rect 9430 17218 9536 17233
rect 9594 17220 9796 17233
rect 9594 17218 9782 17220
rect 9430 17202 9782 17218
rect 9045 17054 11482 17055
rect 9036 17042 11482 17054
rect 9036 17041 11414 17042
rect 8787 16986 11414 17041
rect 11474 16986 11482 17042
rect 8787 16977 11482 16986
rect 8787 16964 9497 16977
rect 8787 16963 9000 16964
rect 9160 16963 9497 16964
rect 4376 16624 5112 16634
rect 4376 16616 4590 16624
rect 4364 16603 4590 16616
rect 4642 16603 5112 16624
rect 4364 16569 4405 16603
rect 4439 16569 4497 16603
rect 4531 16569 4589 16603
rect 4642 16570 4681 16603
rect 4623 16569 4681 16570
rect 4715 16569 4773 16603
rect 4807 16569 4865 16603
rect 4899 16569 4957 16603
rect 4991 16569 5049 16603
rect 5083 16569 5112 16603
rect 4364 16550 5112 16569
rect 4376 16538 5112 16550
rect 4546 16292 4606 16538
rect 5946 16406 6148 16438
rect 5946 16404 6006 16406
rect 5032 16390 6006 16404
rect 5032 16352 5044 16390
rect 5078 16352 6006 16390
rect 5032 16340 6006 16352
rect 6076 16404 6148 16406
rect 6076 16340 6259 16404
rect 5032 16338 6259 16340
rect 5946 16312 6148 16338
rect 4546 16258 4554 16292
rect 4588 16258 4606 16292
rect 4546 16238 4606 16258
rect 4636 16294 4746 16308
rect 4636 16260 4674 16294
rect 4708 16260 4746 16294
rect 4636 16252 4746 16260
rect 4670 16090 4701 16252
rect 4376 16076 5112 16090
rect 4360 16074 5112 16076
rect 4360 16059 4976 16074
rect 5034 16059 5112 16074
rect 4360 16025 4405 16059
rect 4439 16025 4497 16059
rect 4531 16025 4589 16059
rect 4623 16025 4681 16059
rect 4715 16025 4773 16059
rect 4807 16025 4865 16059
rect 4899 16025 4957 16059
rect 5034 16025 5049 16059
rect 5083 16025 5112 16059
rect 4360 16020 4976 16025
rect 5034 16020 5112 16025
rect 4360 16010 5112 16020
rect 4376 15994 5112 16010
rect 4476 15874 5026 15890
rect 4476 15859 4746 15874
rect 4808 15859 5026 15874
rect 4476 15825 4505 15859
rect 4539 15825 4595 15859
rect 4629 15825 4687 15859
rect 4721 15825 4746 15859
rect 4813 15825 4871 15859
rect 4905 15825 4963 15859
rect 4997 15825 5026 15859
rect 4476 15814 4746 15825
rect 4808 15814 5026 15825
rect 4476 15794 5026 15814
rect 4574 15570 4650 15586
rect 4776 15570 4830 15794
rect 6193 15633 6259 16338
rect 6608 15768 7344 15780
rect 6608 15756 6712 15768
rect 6548 15749 6712 15756
rect 6780 15749 7344 15768
rect 6548 15715 6637 15749
rect 6671 15715 6712 15749
rect 6780 15715 6821 15749
rect 6855 15715 6913 15749
rect 6947 15715 7005 15749
rect 7039 15715 7097 15749
rect 7131 15715 7189 15749
rect 7223 15715 7281 15749
rect 7315 15715 7344 15749
rect 6548 15706 6712 15715
rect 6780 15706 7344 15715
rect 6548 15690 7344 15706
rect 6608 15684 7344 15690
rect 4574 15530 4588 15570
rect 4630 15530 4650 15570
rect 4574 15514 4650 15530
rect 4766 15560 4834 15570
rect 6193 15567 7047 15633
rect 6791 15564 6857 15567
rect 4766 15520 4778 15560
rect 4820 15520 4834 15560
rect 4584 15346 4638 15514
rect 4766 15508 4834 15520
rect 4958 15502 5044 15510
rect 4958 15490 4976 15502
rect 4958 15456 4970 15490
rect 4958 15448 4976 15456
rect 5030 15448 5044 15502
rect 4958 15436 5044 15448
rect 5194 15458 6856 15516
rect 5194 15452 6857 15458
rect 4766 15346 4834 15348
rect 4476 15332 5026 15346
rect 4476 15315 4898 15332
rect 4966 15315 5026 15332
rect 4476 15281 4505 15315
rect 4539 15281 4595 15315
rect 4629 15281 4687 15315
rect 4721 15281 4779 15315
rect 4813 15281 4871 15315
rect 4997 15281 5026 15315
rect 4476 15270 4898 15281
rect 4966 15270 5026 15281
rect 4476 15250 5026 15270
rect 4386 15052 5122 15070
rect 4386 15039 4582 15052
rect 4648 15039 5122 15052
rect 4386 15005 4415 15039
rect 4449 15005 4507 15039
rect 4541 15005 4582 15039
rect 4648 15005 4691 15039
rect 4725 15005 4783 15039
rect 4817 15005 4875 15039
rect 4909 15005 4967 15039
rect 5001 15005 5059 15039
rect 5093 15005 5122 15039
rect 4386 14986 4582 15005
rect 4648 14986 5122 15005
rect 4386 14974 5122 14986
rect 4556 14728 4616 14974
rect 5194 14942 5258 15452
rect 6791 15434 6857 15452
rect 6578 15408 6682 15424
rect 6578 15356 6608 15408
rect 6660 15400 6682 15408
rect 6668 15364 6682 15400
rect 6791 15398 6804 15434
rect 6838 15398 6857 15434
rect 6791 15390 6857 15398
rect 6660 15356 6682 15364
rect 6578 15342 6682 15356
rect 6981 15380 7047 15567
rect 7178 15440 7234 15444
rect 7178 15432 7619 15440
rect 7178 15398 7190 15432
rect 7224 15398 7619 15432
rect 7178 15390 7619 15398
rect 7178 15386 7234 15390
rect 7347 15388 7397 15390
rect 6981 15344 6998 15380
rect 7032 15344 7047 15380
rect 6890 15314 6948 15330
rect 6348 15310 6948 15314
rect 5750 15274 6302 15280
rect 5748 15264 6302 15274
rect 6348 15276 6902 15310
rect 6936 15276 6948 15310
rect 6348 15270 6948 15276
rect 5748 15249 6130 15264
rect 6198 15249 6302 15264
rect 5748 15215 5779 15249
rect 5813 15215 5871 15249
rect 5905 15215 5963 15249
rect 5997 15215 6055 15249
rect 6089 15215 6130 15249
rect 6198 15215 6239 15249
rect 6273 15215 6302 15249
rect 5748 15208 6130 15215
rect 5750 15202 6130 15208
rect 6198 15202 6302 15215
rect 5750 15184 6302 15202
rect 6350 15156 6430 15270
rect 6890 15264 6948 15270
rect 6981 15266 7047 15344
rect 6608 15222 7344 15236
rect 6546 15218 7344 15222
rect 6546 15205 7114 15218
rect 7182 15205 7344 15218
rect 6546 15171 6637 15205
rect 6671 15171 6729 15205
rect 6763 15171 6821 15205
rect 6855 15171 6913 15205
rect 6947 15171 7005 15205
rect 7039 15171 7097 15205
rect 7182 15171 7189 15205
rect 7223 15171 7281 15205
rect 7315 15171 7344 15205
rect 6546 15156 7114 15171
rect 7182 15156 7344 15171
rect 6104 15148 6430 15156
rect 5040 14930 5258 14942
rect 5040 14896 5056 14930
rect 5090 14896 5258 14930
rect 5040 14878 5258 14896
rect 5290 15080 6020 15132
rect 6104 15112 6144 15148
rect 6184 15112 6430 15148
rect 6608 15140 7344 15156
rect 6104 15098 6430 15112
rect 4556 14694 4564 14728
rect 4598 14694 4616 14728
rect 4556 14674 4616 14694
rect 4646 14730 4756 14744
rect 4646 14696 4684 14730
rect 4718 14696 4756 14730
rect 4646 14688 4756 14696
rect 4680 14526 4711 14688
rect 4386 14508 5122 14526
rect 4386 14495 5012 14508
rect 5078 14495 5122 14508
rect 4386 14461 4415 14495
rect 4449 14461 4507 14495
rect 4541 14461 4599 14495
rect 4633 14461 4691 14495
rect 4725 14461 4783 14495
rect 4817 14461 4875 14495
rect 4909 14461 4967 14495
rect 5001 14461 5012 14495
rect 5093 14461 5122 14495
rect 4386 14442 5012 14461
rect 5078 14442 5122 14461
rect 4386 14430 5122 14442
rect 4486 14314 5036 14326
rect 4486 14295 4682 14314
rect 4754 14295 5036 14314
rect 4486 14261 4515 14295
rect 4549 14261 4605 14295
rect 4639 14261 4682 14295
rect 4754 14261 4789 14295
rect 4823 14261 4881 14295
rect 4915 14261 4973 14295
rect 5007 14261 5036 14295
rect 4486 14244 4682 14261
rect 4754 14244 5036 14261
rect 4486 14230 5036 14244
rect 4584 14006 4660 14024
rect 4788 14006 4834 14230
rect 4584 13966 4598 14006
rect 4640 13966 4660 14006
rect 4584 13950 4660 13966
rect 4776 13996 4844 14006
rect 4776 13956 4788 13996
rect 4830 13956 4844 13996
rect 4592 13782 4646 13950
rect 4776 13944 4844 13956
rect 4966 13900 5138 13914
rect 4966 13884 5030 13900
rect 4966 13850 4978 13884
rect 5014 13850 5030 13884
rect 4966 13838 5030 13850
rect 5090 13838 5138 13900
rect 4966 13820 5138 13838
rect 4486 13770 5036 13782
rect 4486 13751 4884 13770
rect 4956 13751 5036 13770
rect 4486 13717 4515 13751
rect 4549 13717 4605 13751
rect 4639 13717 4697 13751
rect 4731 13717 4789 13751
rect 4823 13717 4881 13751
rect 4956 13717 4973 13751
rect 5007 13717 5036 13751
rect 4486 13700 4884 13717
rect 4956 13700 5036 13717
rect 4486 13686 5036 13700
rect 4378 13384 5114 13402
rect 4378 13371 4576 13384
rect 4648 13371 5114 13384
rect 4378 13337 4407 13371
rect 4441 13337 4499 13371
rect 4533 13337 4576 13371
rect 4648 13337 4683 13371
rect 4717 13337 4775 13371
rect 4809 13337 4867 13371
rect 4901 13337 4959 13371
rect 4993 13337 5051 13371
rect 5085 13337 5114 13371
rect 4378 13318 4576 13337
rect 4648 13318 5114 13337
rect 4378 13306 5114 13318
rect 5290 13366 5342 15080
rect 5968 14956 6020 15080
rect 5770 14951 5906 14952
rect 5562 14938 5906 14951
rect 5562 14904 5824 14938
rect 5858 14904 5906 14938
rect 5562 14878 5906 14904
rect 5940 14938 6020 14956
rect 5940 14904 5964 14938
rect 6000 14904 6020 14938
rect 5940 14890 6020 14904
rect 5562 14873 5845 14878
rect 5562 13971 5640 14873
rect 5750 14716 6302 14736
rect 5748 14705 5794 14716
rect 5862 14705 6302 14716
rect 5748 14671 5779 14705
rect 5862 14671 5871 14705
rect 5905 14671 5963 14705
rect 5997 14671 6055 14705
rect 6089 14671 6147 14705
rect 6181 14671 6239 14705
rect 6273 14671 6302 14705
rect 5748 14654 5794 14671
rect 5862 14654 6302 14671
rect 5748 14650 6302 14654
rect 5750 14640 6302 14650
rect 7347 14673 7397 14674
rect 7569 14673 7619 15390
rect 7347 14623 7619 14673
rect 5732 14294 6468 14314
rect 5732 14283 6350 14294
rect 6418 14283 6468 14294
rect 5732 14249 5761 14283
rect 5795 14249 5853 14283
rect 5887 14249 5945 14283
rect 5979 14249 6037 14283
rect 6071 14249 6129 14283
rect 6163 14249 6221 14283
rect 6255 14249 6313 14283
rect 6347 14249 6350 14283
rect 6439 14249 6468 14283
rect 5732 14232 6350 14249
rect 6418 14232 6468 14249
rect 5732 14218 6468 14232
rect 7347 14177 7397 14623
rect 7722 14284 8366 14298
rect 7722 14267 7916 14284
rect 7984 14267 8366 14284
rect 7722 14233 7751 14267
rect 7785 14233 7843 14267
rect 7877 14233 7916 14267
rect 7984 14233 8027 14267
rect 8061 14233 8119 14267
rect 8153 14233 8211 14267
rect 8245 14233 8303 14267
rect 8337 14233 8366 14267
rect 7722 14222 7916 14233
rect 7984 14222 8366 14233
rect 7722 14202 8366 14222
rect 7347 14172 7398 14177
rect 7347 14166 8074 14172
rect 7347 14132 7896 14166
rect 7932 14132 8074 14166
rect 7347 14125 8074 14132
rect 7390 14124 8074 14125
rect 8787 14096 8865 16963
rect 9242 16628 9978 16638
rect 9242 16607 9456 16628
rect 9508 16607 9978 16628
rect 9242 16573 9271 16607
rect 9305 16573 9363 16607
rect 9397 16573 9455 16607
rect 9508 16574 9547 16607
rect 9489 16573 9547 16574
rect 9581 16573 9639 16607
rect 9673 16573 9731 16607
rect 9765 16573 9823 16607
rect 9857 16573 9915 16607
rect 9949 16573 9978 16607
rect 9242 16542 9978 16573
rect 9412 16296 9472 16542
rect 10812 16410 11014 16442
rect 10812 16408 10872 16410
rect 9898 16394 10872 16408
rect 9898 16356 9910 16394
rect 9944 16356 10872 16394
rect 9898 16344 10872 16356
rect 10942 16408 11014 16410
rect 10942 16344 11125 16408
rect 9898 16342 11125 16344
rect 10812 16316 11014 16342
rect 9412 16262 9420 16296
rect 9454 16262 9472 16296
rect 9412 16242 9472 16262
rect 9502 16298 9612 16312
rect 9502 16264 9540 16298
rect 9574 16264 9612 16298
rect 9502 16256 9612 16264
rect 9536 16094 9567 16256
rect 9242 16088 9978 16094
rect 9232 16078 9978 16088
rect 9232 16063 9842 16078
rect 9900 16063 9978 16078
rect 9232 16029 9271 16063
rect 9305 16029 9363 16063
rect 9397 16029 9455 16063
rect 9489 16029 9547 16063
rect 9581 16029 9639 16063
rect 9673 16029 9731 16063
rect 9765 16029 9823 16063
rect 9900 16029 9915 16063
rect 9949 16029 9978 16063
rect 9232 16024 9842 16029
rect 9900 16024 9978 16029
rect 9232 16022 9978 16024
rect 9242 15998 9978 16022
rect 9342 15878 9892 15894
rect 9342 15863 9612 15878
rect 9674 15863 9892 15878
rect 9342 15829 9371 15863
rect 9405 15829 9461 15863
rect 9495 15829 9553 15863
rect 9587 15829 9612 15863
rect 9679 15829 9737 15863
rect 9771 15829 9829 15863
rect 9863 15829 9892 15863
rect 9342 15818 9612 15829
rect 9674 15818 9892 15829
rect 9342 15798 9892 15818
rect 9440 15574 9516 15590
rect 9642 15574 9696 15798
rect 11059 15637 11125 16342
rect 11474 15772 12210 15784
rect 11410 15753 11578 15772
rect 11646 15753 12210 15772
rect 11410 15719 11503 15753
rect 11537 15719 11578 15753
rect 11646 15719 11687 15753
rect 11721 15719 11779 15753
rect 11813 15719 11871 15753
rect 11905 15719 11963 15753
rect 11997 15719 12055 15753
rect 12089 15719 12147 15753
rect 12181 15719 12210 15753
rect 11410 15710 11578 15719
rect 11646 15710 12210 15719
rect 11410 15706 12210 15710
rect 11474 15688 12210 15706
rect 9440 15534 9454 15574
rect 9496 15534 9516 15574
rect 9440 15518 9516 15534
rect 9632 15564 9700 15574
rect 11059 15571 11913 15637
rect 11657 15568 11723 15571
rect 9632 15524 9644 15564
rect 9686 15524 9700 15564
rect 9450 15350 9504 15518
rect 9632 15512 9700 15524
rect 9824 15506 9910 15514
rect 9824 15494 9842 15506
rect 9824 15460 9836 15494
rect 9824 15452 9842 15460
rect 9896 15452 9910 15506
rect 9824 15440 9910 15452
rect 10060 15462 11722 15520
rect 10060 15456 11723 15462
rect 9632 15350 9700 15352
rect 9342 15336 9892 15350
rect 9342 15319 9764 15336
rect 9832 15319 9892 15336
rect 9342 15285 9371 15319
rect 9405 15285 9461 15319
rect 9495 15285 9553 15319
rect 9587 15285 9645 15319
rect 9679 15285 9737 15319
rect 9863 15285 9892 15319
rect 9342 15274 9764 15285
rect 9832 15274 9892 15285
rect 9342 15254 9892 15274
rect 9252 15056 9988 15074
rect 9252 15043 9448 15056
rect 9514 15043 9988 15056
rect 9252 15009 9281 15043
rect 9315 15009 9373 15043
rect 9407 15009 9448 15043
rect 9514 15009 9557 15043
rect 9591 15009 9649 15043
rect 9683 15009 9741 15043
rect 9775 15009 9833 15043
rect 9867 15009 9925 15043
rect 9959 15009 9988 15043
rect 9252 14990 9448 15009
rect 9514 14990 9988 15009
rect 9252 14978 9988 14990
rect 9422 14732 9482 14978
rect 10060 14946 10124 15456
rect 11657 15438 11723 15456
rect 11444 15412 11548 15428
rect 11444 15360 11474 15412
rect 11526 15404 11548 15412
rect 11534 15368 11548 15404
rect 11657 15402 11670 15438
rect 11704 15402 11723 15438
rect 11657 15394 11723 15402
rect 11526 15360 11548 15368
rect 11444 15346 11548 15360
rect 11847 15384 11913 15571
rect 12044 15444 12100 15448
rect 12044 15436 12485 15444
rect 12044 15402 12056 15436
rect 12090 15402 12485 15436
rect 12044 15394 12485 15402
rect 12044 15390 12100 15394
rect 12213 15390 12263 15394
rect 11847 15348 11864 15384
rect 11898 15348 11913 15384
rect 11756 15318 11814 15334
rect 11214 15314 11814 15318
rect 10616 15268 11168 15284
rect 11214 15280 11768 15314
rect 11802 15280 11814 15314
rect 11214 15274 11814 15280
rect 10616 15253 10996 15268
rect 11064 15253 11168 15268
rect 10616 15219 10645 15253
rect 10679 15219 10737 15253
rect 10771 15219 10829 15253
rect 10863 15219 10921 15253
rect 10955 15219 10996 15253
rect 11064 15219 11105 15253
rect 11139 15219 11168 15253
rect 10616 15206 10996 15219
rect 11064 15206 11168 15219
rect 10616 15188 11168 15206
rect 11216 15160 11296 15274
rect 11756 15268 11814 15274
rect 11847 15270 11913 15348
rect 11474 15230 12210 15240
rect 11404 15222 12210 15230
rect 11404 15209 11980 15222
rect 12048 15209 12210 15222
rect 11404 15175 11503 15209
rect 11537 15175 11595 15209
rect 11629 15175 11687 15209
rect 11721 15175 11779 15209
rect 11813 15175 11871 15209
rect 11905 15175 11963 15209
rect 12048 15175 12055 15209
rect 12089 15175 12147 15209
rect 12181 15175 12210 15209
rect 11404 15164 11980 15175
rect 10970 15152 11296 15160
rect 9906 14934 10124 14946
rect 9906 14900 9922 14934
rect 9956 14900 10124 14934
rect 9906 14882 10124 14900
rect 10156 15084 10886 15136
rect 10970 15116 11010 15152
rect 11050 15116 11296 15152
rect 11474 15160 11980 15164
rect 12048 15160 12210 15175
rect 11474 15144 12210 15160
rect 10970 15102 11296 15116
rect 9422 14698 9430 14732
rect 9464 14698 9482 14732
rect 9422 14678 9482 14698
rect 9512 14734 9622 14748
rect 9512 14700 9550 14734
rect 9584 14700 9622 14734
rect 9512 14692 9622 14700
rect 9546 14530 9577 14692
rect 9252 14512 9988 14530
rect 9252 14499 9878 14512
rect 9944 14499 9988 14512
rect 9252 14465 9281 14499
rect 9315 14465 9373 14499
rect 9407 14465 9465 14499
rect 9499 14465 9557 14499
rect 9591 14465 9649 14499
rect 9683 14465 9741 14499
rect 9775 14465 9833 14499
rect 9867 14465 9878 14499
rect 9959 14465 9988 14499
rect 9252 14446 9878 14465
rect 9944 14446 9988 14465
rect 9252 14434 9988 14446
rect 9350 14318 9902 14330
rect 9350 14299 9548 14318
rect 9620 14299 9902 14318
rect 9350 14265 9379 14299
rect 9413 14265 9471 14299
rect 9505 14265 9548 14299
rect 9620 14265 9655 14299
rect 9689 14265 9747 14299
rect 9781 14265 9839 14299
rect 9873 14265 9902 14299
rect 9350 14248 9548 14265
rect 9620 14248 9902 14265
rect 9350 14234 9902 14248
rect 7446 14030 8114 14090
rect 5823 13976 5901 14029
rect 7446 14018 7520 14030
rect 5823 13971 5850 13976
rect 5562 13942 5850 13971
rect 5884 13942 5901 13976
rect 5562 13893 5901 13942
rect 5290 13356 5376 13366
rect 4548 13060 4608 13306
rect 5290 13304 5298 13356
rect 5360 13304 5376 13356
rect 5290 13296 5376 13304
rect 5290 13228 5342 13296
rect 5036 13220 5342 13228
rect 5036 13186 5048 13220
rect 5082 13186 5342 13220
rect 5036 13176 5342 13186
rect 5562 13085 5640 13893
rect 6002 13890 6072 13936
rect 6002 13838 6012 13890
rect 6064 13838 6072 13890
rect 6002 13798 6072 13838
rect 6100 13930 6168 13986
rect 6100 13878 6110 13930
rect 6162 13878 6168 13930
rect 6100 13800 6168 13878
rect 6202 13970 6274 13988
rect 6202 13932 6212 13970
rect 6248 13932 6274 13970
rect 6202 13886 6274 13932
rect 6202 13830 6208 13886
rect 6260 13830 6274 13886
rect 6794 13918 7342 13940
rect 6794 13909 6828 13918
rect 6896 13909 7342 13918
rect 6794 13875 6823 13909
rect 6896 13875 6915 13909
rect 6949 13875 7007 13909
rect 7041 13875 7099 13909
rect 7133 13875 7191 13909
rect 7225 13875 7279 13909
rect 7313 13875 7342 13909
rect 6202 13804 6274 13830
rect 6380 13852 6666 13872
rect 6380 13814 6394 13852
rect 6432 13814 6666 13852
rect 6794 13856 6828 13875
rect 6896 13856 7342 13875
rect 6794 13844 7342 13856
rect 7446 13930 7518 14018
rect 7836 13980 7976 13992
rect 7636 13974 7742 13976
rect 7636 13938 7806 13974
rect 7636 13936 7752 13938
rect 6380 13798 6666 13814
rect 6585 13785 6666 13798
rect 7446 13786 7516 13930
rect 7636 13882 7652 13936
rect 7704 13904 7752 13936
rect 7792 13904 7806 13938
rect 7704 13882 7806 13904
rect 7836 13904 7866 13980
rect 7946 13958 7976 13980
rect 8042 13972 8114 14030
rect 8182 14076 8865 14096
rect 8182 14036 8212 14076
rect 8254 14036 8865 14076
rect 8182 14018 8865 14036
rect 8602 13990 8638 14018
rect 9450 14010 9526 14028
rect 9654 14010 9700 14234
rect 7946 13904 7974 13958
rect 8020 13956 8114 13972
rect 8020 13920 8052 13956
rect 8090 13920 8114 13956
rect 9450 13970 9464 14010
rect 9506 13970 9526 14010
rect 9450 13954 9526 13970
rect 9642 14000 9710 14010
rect 9642 13960 9654 14000
rect 9696 13960 9710 14000
rect 8020 13904 8114 13920
rect 7836 13890 7974 13904
rect 7636 13856 7806 13882
rect 9458 13786 9512 13954
rect 9642 13948 9710 13960
rect 9832 13904 10004 13918
rect 9832 13888 9896 13904
rect 9832 13854 9844 13888
rect 9880 13854 9896 13888
rect 9832 13842 9896 13854
rect 9956 13842 10004 13904
rect 9832 13824 10004 13842
rect 5732 13754 6468 13770
rect 5732 13739 5862 13754
rect 5930 13739 6468 13754
rect 5732 13705 5761 13739
rect 5795 13705 5853 13739
rect 5930 13705 5945 13739
rect 5979 13705 6037 13739
rect 6071 13705 6129 13739
rect 6163 13705 6221 13739
rect 6255 13705 6313 13739
rect 6347 13705 6405 13739
rect 6439 13705 6468 13739
rect 6585 13711 7063 13785
rect 7120 13764 7516 13786
rect 7120 13730 7162 13764
rect 7196 13730 7516 13764
rect 9350 13774 9902 13786
rect 9350 13755 9750 13774
rect 9822 13755 9902 13774
rect 7120 13714 7516 13730
rect 7640 13738 8366 13754
rect 5732 13692 5862 13705
rect 5930 13692 6468 13705
rect 5732 13674 6468 13692
rect 6989 13604 7063 13711
rect 7640 13676 7656 13738
rect 7724 13723 8366 13738
rect 7724 13689 7751 13723
rect 7785 13689 7843 13723
rect 7877 13689 7935 13723
rect 7969 13689 8027 13723
rect 8061 13689 8119 13723
rect 8153 13689 8211 13723
rect 8245 13689 8303 13723
rect 8337 13689 8366 13723
rect 9350 13721 9379 13755
rect 9413 13721 9471 13755
rect 9505 13721 9563 13755
rect 9597 13721 9655 13755
rect 9689 13721 9747 13755
rect 9822 13721 9839 13755
rect 9873 13721 9902 13755
rect 9350 13704 9750 13721
rect 9822 13704 9902 13721
rect 9350 13690 9902 13704
rect 7724 13676 8366 13689
rect 7640 13658 8366 13676
rect 7640 13656 7734 13658
rect 6544 13554 6893 13577
rect 6544 13520 6834 13554
rect 6868 13520 6893 13554
rect 6544 13503 6893 13520
rect 6989 13570 7012 13604
rect 7046 13570 7063 13604
rect 5856 13450 6408 13472
rect 5856 13441 5984 13450
rect 6052 13441 6408 13450
rect 5856 13407 5885 13441
rect 5919 13407 5977 13441
rect 6052 13407 6069 13441
rect 6103 13407 6161 13441
rect 6195 13407 6253 13441
rect 6287 13407 6345 13441
rect 6379 13407 6408 13441
rect 5856 13390 5984 13407
rect 6052 13390 6408 13407
rect 5856 13376 6408 13390
rect 6120 13338 6218 13344
rect 6120 13286 6140 13338
rect 6194 13286 6218 13338
rect 6544 13298 6618 13503
rect 6989 13489 7063 13570
rect 6794 13378 7342 13396
rect 6794 13365 7136 13378
rect 7204 13365 7342 13378
rect 6794 13331 6823 13365
rect 6857 13331 6915 13365
rect 6949 13331 7007 13365
rect 7041 13331 7099 13365
rect 7133 13331 7136 13365
rect 7225 13331 7279 13365
rect 7313 13331 7342 13365
rect 6794 13316 7136 13331
rect 7204 13316 7342 13331
rect 6794 13300 7342 13316
rect 9244 13388 9980 13406
rect 9244 13375 9442 13388
rect 9514 13375 9980 13388
rect 9244 13341 9273 13375
rect 9307 13341 9365 13375
rect 9399 13341 9442 13375
rect 9514 13341 9549 13375
rect 9583 13341 9641 13375
rect 9675 13341 9733 13375
rect 9767 13341 9825 13375
rect 9859 13341 9917 13375
rect 9951 13341 9980 13375
rect 9244 13322 9442 13341
rect 9514 13322 9980 13341
rect 9244 13310 9980 13322
rect 10156 13370 10208 15084
rect 10834 14960 10886 15084
rect 10636 14955 10772 14956
rect 10428 14942 10772 14955
rect 10428 14908 10690 14942
rect 10724 14908 10772 14942
rect 10428 14882 10772 14908
rect 10806 14942 10886 14960
rect 10806 14908 10830 14942
rect 10866 14908 10886 14942
rect 10806 14894 10886 14908
rect 10428 14877 10711 14882
rect 10428 13975 10506 14877
rect 12435 14741 12485 15394
rect 12341 14740 12485 14741
rect 10616 14720 11168 14740
rect 10616 14709 10660 14720
rect 10728 14709 11168 14720
rect 10616 14675 10645 14709
rect 10728 14675 10737 14709
rect 10771 14675 10829 14709
rect 10863 14675 10921 14709
rect 10955 14675 11013 14709
rect 11047 14675 11105 14709
rect 11139 14675 11168 14709
rect 12209 14691 12485 14740
rect 13643 14697 13733 17497
rect 16399 17468 16461 17478
rect 16399 17466 16413 17468
rect 15360 17436 15683 17458
rect 14960 17407 15635 17436
rect 14960 16366 14989 17407
rect 15360 17402 15635 17407
rect 15669 17402 15683 17436
rect 15360 17368 15683 17402
rect 15713 17428 15902 17448
rect 15713 17394 15725 17428
rect 15763 17411 15902 17428
rect 15943 17436 16413 17466
rect 15943 17411 15973 17436
rect 16187 17434 16217 17436
rect 16399 17434 16413 17436
rect 16449 17434 16461 17468
rect 15763 17394 15973 17411
rect 16399 17410 16461 17434
rect 16493 17476 17335 17498
rect 16493 17464 17287 17476
rect 16493 17430 16517 17464
rect 16551 17442 17287 17464
rect 17321 17442 17335 17476
rect 16551 17430 17335 17442
rect 16493 17408 17335 17430
rect 17365 17472 18103 17488
rect 17365 17468 18059 17472
rect 17365 17434 17377 17468
rect 17415 17438 18059 17468
rect 18097 17438 18103 17472
rect 17415 17434 18103 17438
rect 17365 17414 18103 17434
rect 18133 17474 18201 17490
rect 18133 17472 19179 17474
rect 18133 17462 19225 17472
rect 18133 17460 19177 17462
rect 18133 17426 18147 17460
rect 18183 17428 19177 17460
rect 19213 17428 19225 17462
rect 18183 17426 19225 17428
rect 18133 17418 19225 17426
rect 18133 17406 18201 17418
rect 19163 17404 19225 17418
rect 19257 17470 20099 17492
rect 20897 17483 20963 17484
rect 19257 17458 20051 17470
rect 19257 17424 19281 17458
rect 19315 17436 20051 17458
rect 20085 17436 20099 17470
rect 19315 17424 20099 17436
rect 19257 17402 20099 17424
rect 20129 17466 20867 17482
rect 20129 17462 20823 17466
rect 20129 17428 20141 17462
rect 20179 17432 20823 17462
rect 20861 17432 20867 17466
rect 20179 17428 20867 17432
rect 20129 17408 20867 17428
rect 20897 17468 21107 17483
rect 20897 17462 21425 17468
rect 20897 17454 21481 17462
rect 20897 17420 20911 17454
rect 20947 17452 21481 17454
rect 20947 17422 21433 17452
rect 20947 17420 20963 17422
rect 21305 17420 21433 17422
rect 20897 17400 20963 17420
rect 21419 17418 21433 17420
rect 21469 17418 21481 17452
rect 21419 17394 21481 17418
rect 21513 17460 22355 17482
rect 23153 17473 23219 17474
rect 21513 17448 22307 17460
rect 21513 17414 21537 17448
rect 21571 17426 22307 17448
rect 22341 17426 22355 17460
rect 21571 17414 22355 17426
rect 15713 17381 15973 17394
rect 21513 17392 22355 17414
rect 22385 17456 23123 17472
rect 22385 17452 23079 17456
rect 22385 17418 22397 17452
rect 22435 17422 23079 17452
rect 23117 17422 23123 17456
rect 22435 17418 23123 17422
rect 22385 17398 23123 17418
rect 23153 17444 23432 17473
rect 23153 17410 23167 17444
rect 23203 17443 23432 17444
rect 23203 17410 23219 17443
rect 23153 17390 23219 17410
rect 15713 17374 15902 17381
rect 16267 17172 16621 17188
rect 16267 17157 16453 17172
rect 16521 17157 16621 17172
rect 15481 17134 15843 17150
rect 15481 17119 15691 17134
rect 15759 17119 15843 17134
rect 15481 17085 15510 17119
rect 15544 17085 15596 17119
rect 15630 17085 15688 17119
rect 15759 17085 15780 17119
rect 15814 17085 15843 17119
rect 16267 17123 16296 17157
rect 16330 17123 16374 17157
rect 16408 17123 16453 17157
rect 16521 17123 16558 17157
rect 16592 17123 16621 17157
rect 16267 17110 16453 17123
rect 16521 17110 16621 17123
rect 16267 17092 16621 17110
rect 17133 17174 17495 17190
rect 17133 17159 17343 17174
rect 17411 17159 17495 17174
rect 17911 17166 18263 17180
rect 17911 17160 18101 17166
rect 17133 17125 17162 17159
rect 17196 17125 17248 17159
rect 17282 17125 17340 17159
rect 17411 17125 17432 17159
rect 17466 17125 17495 17159
rect 17133 17112 17343 17125
rect 17411 17112 17495 17125
rect 17133 17094 17495 17112
rect 17905 17149 18101 17160
rect 18169 17149 18263 17166
rect 17905 17115 17940 17149
rect 17974 17115 18016 17149
rect 18050 17115 18101 17149
rect 18169 17115 18200 17149
rect 18234 17115 18263 17149
rect 17905 17104 18101 17115
rect 18169 17104 18263 17115
rect 17905 17094 18263 17104
rect 15481 17072 15691 17085
rect 15759 17072 15843 17085
rect 17911 17084 18263 17094
rect 19027 17166 19385 17182
rect 19027 17151 19217 17166
rect 19285 17151 19385 17166
rect 19027 17117 19056 17151
rect 19090 17117 19138 17151
rect 19172 17117 19217 17151
rect 19285 17117 19322 17151
rect 19356 17117 19385 17151
rect 19027 17104 19217 17117
rect 19285 17104 19385 17117
rect 19027 17086 19385 17104
rect 19893 17168 20259 17184
rect 19893 17153 20107 17168
rect 20175 17153 20259 17168
rect 19893 17119 19922 17153
rect 19956 17119 20012 17153
rect 20046 17119 20104 17153
rect 20175 17119 20196 17153
rect 20230 17119 20259 17153
rect 19893 17106 20107 17119
rect 20175 17106 20259 17119
rect 19893 17088 20259 17106
rect 20663 17160 21027 17174
rect 20663 17143 20865 17160
rect 20933 17143 21027 17160
rect 20663 17109 20692 17143
rect 20726 17109 20780 17143
rect 20814 17109 20865 17143
rect 20933 17109 20964 17143
rect 20998 17109 21027 17143
rect 20663 17098 20865 17109
rect 20933 17098 21027 17109
rect 20663 17078 21027 17098
rect 21365 17156 21733 17172
rect 21365 17141 21473 17156
rect 21541 17141 21733 17156
rect 21365 17107 21394 17141
rect 21428 17107 21473 17141
rect 21541 17107 21578 17141
rect 21612 17107 21670 17141
rect 21704 17107 21733 17141
rect 21365 17094 21473 17107
rect 21541 17094 21733 17107
rect 21365 17076 21733 17094
rect 22149 17158 22515 17174
rect 22149 17143 22363 17158
rect 22431 17143 22515 17158
rect 22149 17109 22178 17143
rect 22212 17109 22268 17143
rect 22302 17109 22360 17143
rect 22431 17109 22452 17143
rect 22486 17109 22515 17143
rect 22149 17096 22363 17109
rect 22431 17096 22515 17109
rect 22149 17078 22515 17096
rect 23007 17150 23373 17164
rect 23007 17133 23121 17150
rect 23189 17133 23373 17150
rect 23007 17099 23036 17133
rect 23070 17099 23121 17133
rect 23189 17099 23220 17133
rect 23254 17099 23310 17133
rect 23344 17099 23373 17133
rect 23007 17088 23121 17099
rect 23189 17088 23373 17099
rect 15481 17054 15843 17072
rect 23007 17068 23373 17088
rect 23402 16937 23432 17443
rect 23402 16906 23479 16937
rect 23403 16877 23479 16906
rect 16246 16722 16612 16742
rect 16246 16711 16430 16722
rect 16498 16711 16612 16722
rect 16246 16677 16275 16711
rect 16309 16677 16365 16711
rect 16399 16677 16430 16711
rect 16498 16677 16549 16711
rect 16583 16677 16612 16711
rect 16246 16660 16430 16677
rect 16498 16660 16612 16677
rect 16246 16646 16612 16660
rect 17104 16714 17470 16732
rect 17104 16701 17188 16714
rect 17256 16701 17470 16714
rect 17104 16667 17133 16701
rect 17167 16667 17188 16701
rect 17259 16667 17317 16701
rect 17351 16667 17407 16701
rect 17441 16667 17470 16701
rect 17104 16652 17188 16667
rect 17256 16652 17470 16667
rect 17104 16636 17470 16652
rect 17886 16716 18254 16734
rect 17886 16703 18078 16716
rect 18146 16703 18254 16716
rect 17886 16669 17915 16703
rect 17949 16669 18007 16703
rect 18041 16669 18078 16703
rect 18146 16669 18191 16703
rect 18225 16669 18254 16703
rect 17886 16654 18078 16669
rect 18146 16654 18254 16669
rect 17886 16638 18254 16654
rect 18592 16712 18956 16732
rect 18592 16701 18686 16712
rect 18754 16701 18956 16712
rect 18592 16667 18621 16701
rect 18655 16667 18686 16701
rect 18754 16667 18805 16701
rect 18839 16667 18893 16701
rect 18927 16667 18956 16701
rect 18592 16650 18686 16667
rect 18754 16650 18956 16667
rect 18592 16636 18956 16650
rect 19360 16704 19726 16722
rect 19360 16691 19444 16704
rect 19512 16691 19726 16704
rect 19360 16657 19389 16691
rect 19423 16657 19444 16691
rect 19515 16657 19573 16691
rect 19607 16657 19663 16691
rect 19697 16657 19726 16691
rect 19360 16642 19444 16657
rect 19512 16642 19726 16657
rect 19360 16626 19726 16642
rect 20234 16706 20592 16724
rect 20234 16693 20334 16706
rect 20402 16693 20592 16706
rect 20234 16659 20263 16693
rect 20297 16659 20334 16693
rect 20402 16659 20447 16693
rect 20481 16659 20529 16693
rect 20563 16659 20592 16693
rect 20234 16644 20334 16659
rect 20402 16644 20592 16659
rect 20234 16628 20592 16644
rect 21356 16716 21708 16726
rect 21356 16706 21714 16716
rect 21356 16695 21450 16706
rect 21518 16695 21714 16706
rect 21356 16661 21385 16695
rect 21419 16661 21450 16695
rect 21518 16661 21569 16695
rect 21603 16661 21645 16695
rect 21679 16661 21714 16695
rect 21356 16644 21450 16661
rect 21518 16650 21714 16661
rect 22124 16698 22486 16716
rect 22124 16685 22208 16698
rect 22276 16685 22486 16698
rect 22124 16651 22153 16685
rect 22187 16651 22208 16685
rect 22279 16651 22337 16685
rect 22371 16651 22423 16685
rect 22457 16651 22486 16685
rect 21518 16644 21708 16650
rect 21356 16630 21708 16644
rect 22124 16636 22208 16651
rect 22276 16636 22486 16651
rect 22124 16620 22486 16636
rect 22998 16700 23352 16718
rect 22998 16687 23098 16700
rect 23166 16687 23352 16700
rect 22998 16653 23027 16687
rect 23061 16653 23098 16687
rect 23166 16653 23211 16687
rect 23245 16653 23289 16687
rect 23323 16653 23352 16687
rect 22998 16638 23098 16653
rect 23166 16638 23352 16653
rect 22998 16622 23352 16638
rect 16400 16400 16466 16420
rect 16400 16367 16416 16400
rect 16224 16366 16416 16367
rect 16452 16366 16466 16400
rect 14960 16337 16466 16366
rect 16496 16392 17234 16412
rect 16496 16388 17184 16392
rect 16496 16354 16502 16388
rect 16540 16358 17184 16388
rect 17222 16358 17234 16392
rect 16540 16354 17234 16358
rect 16496 16338 17234 16354
rect 17264 16396 18106 16418
rect 17264 16384 18048 16396
rect 17264 16350 17278 16384
rect 17312 16362 18048 16384
rect 18082 16362 18106 16396
rect 17312 16350 18106 16362
rect 16400 16336 16466 16337
rect 17264 16328 18106 16350
rect 18138 16392 18200 16416
rect 18138 16358 18150 16392
rect 18186 16390 18200 16392
rect 18656 16390 18722 16410
rect 18186 16388 18314 16390
rect 18656 16388 18672 16390
rect 18186 16358 18672 16388
rect 18138 16356 18672 16358
rect 18708 16356 18722 16390
rect 18138 16348 18722 16356
rect 18194 16342 18722 16348
rect 18512 16327 18722 16342
rect 18752 16382 19490 16402
rect 18752 16378 19440 16382
rect 18752 16344 18758 16378
rect 18796 16348 19440 16378
rect 19478 16348 19490 16382
rect 18796 16344 19490 16348
rect 18752 16328 19490 16344
rect 19520 16386 20362 16408
rect 19520 16374 20304 16386
rect 19520 16340 19534 16374
rect 19568 16352 20304 16374
rect 20338 16352 20362 16386
rect 19568 16340 20362 16352
rect 18656 16326 18722 16327
rect 19520 16318 20362 16340
rect 20394 16392 20456 16406
rect 21418 16392 21486 16404
rect 20394 16384 21486 16392
rect 20394 16382 21436 16384
rect 20394 16348 20406 16382
rect 20442 16350 21436 16382
rect 21472 16350 21486 16384
rect 20442 16348 21486 16350
rect 20394 16338 21486 16348
rect 20440 16336 21486 16338
rect 21418 16320 21486 16336
rect 21516 16376 22254 16396
rect 21516 16372 22204 16376
rect 21516 16338 21522 16372
rect 21560 16342 22204 16372
rect 22242 16342 22254 16376
rect 21560 16338 22254 16342
rect 21516 16322 22254 16338
rect 22284 16380 23126 16402
rect 22284 16368 23068 16380
rect 22284 16334 22298 16368
rect 22332 16346 23068 16368
rect 23102 16346 23126 16380
rect 22332 16334 23126 16346
rect 22284 16312 23126 16334
rect 23158 16376 23220 16400
rect 23158 16342 23170 16376
rect 23206 16374 23220 16376
rect 23449 16374 23479 16877
rect 23206 16344 23479 16374
rect 23206 16342 23220 16344
rect 23158 16332 23220 16342
rect 16246 16184 16612 16198
rect 16246 16167 16410 16184
rect 16478 16167 16612 16184
rect 16246 16133 16275 16167
rect 16309 16133 16365 16167
rect 16399 16133 16410 16167
rect 16491 16133 16549 16167
rect 16583 16133 16612 16167
rect 16246 16122 16410 16133
rect 16478 16122 16612 16133
rect 16246 16102 16612 16122
rect 17104 16174 17470 16188
rect 17104 16157 17196 16174
rect 17264 16157 17470 16174
rect 17104 16123 17133 16157
rect 17167 16123 17196 16157
rect 17264 16123 17317 16157
rect 17351 16123 17407 16157
rect 17441 16123 17470 16157
rect 17104 16112 17196 16123
rect 17264 16112 17470 16123
rect 17104 16092 17470 16112
rect 17886 16174 18254 16190
rect 17886 16159 18076 16174
rect 18144 16159 18254 16174
rect 17886 16125 17915 16159
rect 17949 16125 18007 16159
rect 18041 16125 18076 16159
rect 18144 16125 18191 16159
rect 18225 16125 18254 16159
rect 17886 16112 18076 16125
rect 18144 16112 18254 16125
rect 17886 16094 18254 16112
rect 18592 16174 18956 16188
rect 18592 16157 18666 16174
rect 18734 16157 18956 16174
rect 18592 16123 18621 16157
rect 18655 16123 18666 16157
rect 18747 16123 18805 16157
rect 18839 16123 18893 16157
rect 18927 16123 18956 16157
rect 18592 16112 18666 16123
rect 18734 16112 18956 16123
rect 18592 16092 18956 16112
rect 19360 16164 19726 16178
rect 19360 16147 19452 16164
rect 19520 16147 19726 16164
rect 19360 16113 19389 16147
rect 19423 16113 19452 16147
rect 19520 16113 19573 16147
rect 19607 16113 19663 16147
rect 19697 16113 19726 16147
rect 19360 16102 19452 16113
rect 19520 16102 19726 16113
rect 19360 16082 19726 16102
rect 20234 16170 20592 16180
rect 21356 16178 21708 16182
rect 20234 16164 20594 16170
rect 20234 16149 20332 16164
rect 20400 16149 20594 16164
rect 20234 16115 20263 16149
rect 20297 16115 20332 16149
rect 20400 16115 20447 16149
rect 20481 16115 20529 16149
rect 20563 16115 20594 16149
rect 20234 16102 20332 16115
rect 20400 16104 20594 16115
rect 21356 16168 21710 16178
rect 21356 16151 21430 16168
rect 21498 16151 21710 16168
rect 21356 16117 21385 16151
rect 21419 16117 21430 16151
rect 21511 16117 21569 16151
rect 21603 16117 21645 16151
rect 21679 16117 21710 16151
rect 21356 16106 21430 16117
rect 21498 16112 21710 16117
rect 22124 16158 22486 16172
rect 22124 16141 22216 16158
rect 22284 16141 22486 16158
rect 21498 16106 21708 16112
rect 20400 16102 20592 16104
rect 20234 16084 20592 16102
rect 21356 16086 21708 16106
rect 22124 16107 22153 16141
rect 22187 16107 22216 16141
rect 22284 16107 22337 16141
rect 22371 16107 22423 16141
rect 22457 16107 22486 16141
rect 22124 16096 22216 16107
rect 22284 16096 22486 16107
rect 22124 16076 22486 16096
rect 22998 16158 23352 16174
rect 22998 16143 23096 16158
rect 23164 16143 23352 16158
rect 22998 16109 23027 16143
rect 23061 16109 23096 16143
rect 23164 16109 23211 16143
rect 23245 16109 23289 16143
rect 23323 16109 23352 16143
rect 22998 16096 23096 16109
rect 23164 16096 23352 16109
rect 22998 16078 23352 16096
rect 23373 15915 23403 15918
rect 23449 15915 23479 16344
rect 23373 15885 23479 15915
rect 23373 15607 23403 15885
rect 23372 15606 23403 15607
rect 22975 15577 23403 15606
rect 22975 14749 23005 15577
rect 23484 14870 25508 14880
rect 23484 14849 24400 14870
rect 24462 14849 25508 14870
rect 23484 14815 23513 14849
rect 23547 14815 23605 14849
rect 23639 14815 23697 14849
rect 23731 14815 23789 14849
rect 23823 14815 23881 14849
rect 23915 14815 23973 14849
rect 24007 14815 24065 14849
rect 24099 14815 24157 14849
rect 24191 14815 24249 14849
rect 24283 14815 24341 14849
rect 24375 14815 24400 14849
rect 24467 14815 24525 14849
rect 24559 14815 24617 14849
rect 24651 14815 24709 14849
rect 24743 14815 24801 14849
rect 24835 14815 24893 14849
rect 24927 14815 24985 14849
rect 25019 14815 25077 14849
rect 25111 14815 25169 14849
rect 25203 14815 25261 14849
rect 25295 14815 25353 14849
rect 25387 14815 25445 14849
rect 25479 14815 25508 14849
rect 23484 14810 24400 14815
rect 24462 14810 25508 14815
rect 23484 14784 25508 14810
rect 22975 14719 23418 14749
rect 10616 14658 10660 14675
rect 10728 14658 11168 14675
rect 10616 14644 11168 14658
rect 10598 14298 11334 14318
rect 10598 14287 11216 14298
rect 11284 14287 11334 14298
rect 10598 14253 10627 14287
rect 10661 14253 10719 14287
rect 10753 14253 10811 14287
rect 10845 14253 10903 14287
rect 10937 14253 10995 14287
rect 11029 14253 11087 14287
rect 11121 14253 11179 14287
rect 11213 14253 11216 14287
rect 11305 14253 11334 14287
rect 10598 14236 11216 14253
rect 11284 14236 11334 14253
rect 10598 14222 11334 14236
rect 12213 14181 12263 14691
rect 13643 14607 22797 14697
rect 23388 14675 23418 14719
rect 24138 14714 24198 14726
rect 23388 14674 23700 14675
rect 23388 14645 23731 14674
rect 23701 14614 23731 14645
rect 24138 14662 24144 14714
rect 24196 14662 24198 14714
rect 24138 14650 24198 14662
rect 24138 14616 24150 14650
rect 24186 14616 24198 14650
rect 24337 14679 24395 14685
rect 24337 14645 24349 14679
rect 24383 14676 24395 14679
rect 24983 14679 25041 14685
rect 24983 14676 24995 14679
rect 24383 14648 24995 14676
rect 24383 14645 24395 14648
rect 24337 14639 24395 14645
rect 24983 14645 24995 14648
rect 25029 14645 25041 14679
rect 25917 14658 26063 18339
rect 24983 14639 25041 14645
rect 12588 14288 13232 14302
rect 12588 14271 12782 14288
rect 12850 14271 13232 14288
rect 12588 14237 12617 14271
rect 12651 14237 12709 14271
rect 12743 14237 12782 14271
rect 12850 14237 12893 14271
rect 12927 14237 12985 14271
rect 13019 14237 13077 14271
rect 13111 14237 13169 14271
rect 13203 14237 13232 14271
rect 12588 14226 12782 14237
rect 12850 14226 13232 14237
rect 12588 14206 13232 14226
rect 13643 14182 13733 14607
rect 22618 14599 22797 14607
rect 22618 14580 23581 14599
rect 22618 14546 23530 14580
rect 23568 14546 23581 14580
rect 22618 14509 23581 14546
rect 23644 14562 23732 14614
rect 24138 14578 24198 14616
rect 23644 14528 23672 14562
rect 23708 14528 23732 14562
rect 24444 14564 24510 14620
rect 22618 14508 22736 14509
rect 23644 14490 23732 14528
rect 23962 14543 24020 14549
rect 23962 14509 23974 14543
rect 24008 14540 24020 14543
rect 24330 14543 24388 14549
rect 24330 14540 24342 14543
rect 24008 14512 24342 14540
rect 24008 14509 24020 14512
rect 23962 14503 24020 14509
rect 24330 14509 24342 14512
rect 24376 14509 24388 14543
rect 24330 14503 24388 14509
rect 24444 14512 24452 14564
rect 24504 14512 24510 14564
rect 24444 14502 24510 14512
rect 24550 14588 24604 14620
rect 24550 14578 24556 14588
rect 24592 14578 24604 14588
rect 24550 14526 24552 14578
rect 24550 14502 24604 14526
rect 24684 14602 24770 14618
rect 24684 14550 24698 14602
rect 24750 14550 24770 14602
rect 24684 14528 24712 14550
rect 24746 14528 24770 14550
rect 25348 14594 26063 14658
rect 25348 14560 25356 14594
rect 25390 14560 26063 14594
rect 24684 14518 24770 14528
rect 24799 14543 24857 14549
rect 24799 14509 24811 14543
rect 24845 14540 24857 14543
rect 25167 14543 25225 14549
rect 25167 14540 25179 14543
rect 24845 14512 25179 14540
rect 24845 14509 24857 14512
rect 24799 14503 24857 14509
rect 25167 14509 25179 14512
rect 25213 14509 25225 14543
rect 25348 14516 26063 14560
rect 25917 14514 26063 14516
rect 25167 14503 25225 14509
rect 23778 14475 23836 14481
rect 23778 14441 23790 14475
rect 23824 14472 23836 14475
rect 24882 14475 24940 14481
rect 24882 14472 24894 14475
rect 23824 14444 24894 14472
rect 23824 14441 23836 14444
rect 23778 14435 23836 14441
rect 24882 14441 24894 14444
rect 24928 14472 24940 14475
rect 25066 14475 25124 14481
rect 25066 14472 25078 14475
rect 24928 14444 25078 14472
rect 24928 14441 24940 14444
rect 24882 14435 24940 14441
rect 25066 14441 25078 14444
rect 25112 14441 25124 14475
rect 25066 14435 25124 14441
rect 23484 14318 25508 14336
rect 23484 14305 23992 14318
rect 24054 14305 25508 14318
rect 23484 14271 23513 14305
rect 23547 14271 23605 14305
rect 23639 14271 23697 14305
rect 23731 14271 23789 14305
rect 23823 14271 23881 14305
rect 23915 14271 23973 14305
rect 24054 14271 24065 14305
rect 24099 14271 24157 14305
rect 24191 14271 24249 14305
rect 24283 14271 24341 14305
rect 24375 14271 24433 14305
rect 24467 14271 24525 14305
rect 24559 14271 24617 14305
rect 24651 14271 24709 14305
rect 24743 14271 24801 14305
rect 24835 14271 24893 14305
rect 24927 14271 24985 14305
rect 25019 14271 25077 14305
rect 25111 14271 25169 14305
rect 25203 14271 25261 14305
rect 25295 14271 25353 14305
rect 25387 14271 25445 14305
rect 25479 14271 25508 14305
rect 23484 14258 23992 14271
rect 24054 14258 25508 14271
rect 23484 14240 25508 14258
rect 12213 14176 12264 14181
rect 12213 14170 12940 14176
rect 12213 14136 12762 14170
rect 12798 14136 12940 14170
rect 12213 14129 12940 14136
rect 12256 14128 12940 14129
rect 13470 14132 13733 14182
rect 13470 14100 13732 14132
rect 12312 14034 12980 14094
rect 10689 13980 10767 14033
rect 12312 14022 12386 14034
rect 10689 13975 10716 13980
rect 10428 13946 10716 13975
rect 10750 13946 10767 13980
rect 10428 13897 10767 13946
rect 10156 13360 10242 13370
rect 6120 13268 6218 13286
rect 6332 13278 6618 13298
rect 6332 13240 6342 13278
rect 6380 13240 6618 13278
rect 6332 13224 6618 13240
rect 4548 13026 4556 13060
rect 4590 13026 4608 13060
rect 4548 13006 4608 13026
rect 4638 13062 4748 13076
rect 4638 13028 4676 13062
rect 4710 13028 4748 13062
rect 4638 13020 4748 13028
rect 5562 13060 6081 13085
rect 5562 13026 5994 13060
rect 6028 13026 6081 13060
rect 4672 12858 4703 13020
rect 5562 13007 6081 13026
rect 6176 13082 6258 13154
rect 6176 13028 6196 13082
rect 6248 13028 6258 13082
rect 4378 12844 5114 12858
rect 4378 12827 4990 12844
rect 5062 12827 5114 12844
rect 4378 12793 4407 12827
rect 4441 12793 4499 12827
rect 4533 12793 4591 12827
rect 4625 12793 4683 12827
rect 4717 12793 4775 12827
rect 4809 12793 4867 12827
rect 4901 12793 4959 12827
rect 5085 12793 5114 12827
rect 4378 12778 4990 12793
rect 5062 12778 5114 12793
rect 4378 12762 5114 12778
rect 4478 12642 5028 12658
rect 4478 12627 4634 12642
rect 4708 12627 5028 12642
rect 4478 12593 4507 12627
rect 4541 12593 4597 12627
rect 4631 12593 4634 12627
rect 4723 12593 4781 12627
rect 4815 12593 4873 12627
rect 4907 12593 4965 12627
rect 4999 12593 5028 12627
rect 4478 12576 4634 12593
rect 4708 12576 5028 12593
rect 4478 12562 5028 12576
rect 4576 12338 4652 12364
rect 4776 12338 4826 12562
rect 4960 12390 5110 12404
rect 4960 12370 5006 12390
rect 4576 12298 4590 12338
rect 4632 12298 4652 12338
rect 4576 12282 4652 12298
rect 4768 12328 4836 12338
rect 4768 12288 4780 12328
rect 4822 12288 4836 12328
rect 4960 12336 4970 12370
rect 4960 12322 5006 12336
rect 5068 12322 5110 12390
rect 4960 12306 5110 12322
rect 4590 12114 4642 12282
rect 4768 12276 4836 12288
rect 5562 12121 5640 13007
rect 6176 12970 6258 13028
rect 9414 13064 9474 13310
rect 10156 13308 10164 13360
rect 10226 13308 10242 13360
rect 10156 13300 10242 13308
rect 10156 13232 10208 13300
rect 9902 13224 10208 13232
rect 9902 13190 9914 13224
rect 9948 13190 10208 13224
rect 9902 13180 10208 13190
rect 10428 13089 10506 13897
rect 10868 13894 10938 13940
rect 10868 13842 10878 13894
rect 10930 13842 10938 13894
rect 10868 13802 10938 13842
rect 10966 13934 11034 13990
rect 10966 13882 10976 13934
rect 11028 13882 11034 13934
rect 10966 13804 11034 13882
rect 11068 13974 11140 13992
rect 11068 13936 11078 13974
rect 11114 13936 11140 13974
rect 11068 13890 11140 13936
rect 11068 13834 11074 13890
rect 11126 13834 11140 13890
rect 11660 13922 12210 13944
rect 11660 13913 11694 13922
rect 11762 13913 12210 13922
rect 11660 13879 11689 13913
rect 11762 13879 11781 13913
rect 11815 13879 11873 13913
rect 11907 13879 11965 13913
rect 11999 13879 12057 13913
rect 12091 13879 12147 13913
rect 12181 13879 12210 13913
rect 11068 13808 11140 13834
rect 11246 13856 11532 13876
rect 11246 13818 11260 13856
rect 11298 13818 11532 13856
rect 11660 13860 11694 13879
rect 11762 13860 12210 13879
rect 11660 13848 12210 13860
rect 12312 13934 12384 14022
rect 12702 13984 12842 13996
rect 12502 13978 12608 13980
rect 12502 13942 12672 13978
rect 12502 13940 12618 13942
rect 11246 13802 11532 13818
rect 11451 13789 11532 13802
rect 12312 13790 12382 13934
rect 12502 13886 12518 13940
rect 12570 13908 12618 13940
rect 12658 13908 12672 13942
rect 12570 13886 12672 13908
rect 12702 13908 12732 13984
rect 12812 13962 12842 13984
rect 12908 13976 12980 14034
rect 13048 14080 13732 14100
rect 13048 14040 13078 14080
rect 13120 14040 13732 14080
rect 13048 14022 13732 14040
rect 13468 13996 13732 14022
rect 13468 13994 13504 13996
rect 12812 13908 12840 13962
rect 12886 13960 12980 13976
rect 12886 13924 12918 13960
rect 12956 13924 12980 13960
rect 12886 13908 12980 13924
rect 12702 13894 12840 13908
rect 12502 13860 12672 13886
rect 10598 13758 11334 13774
rect 10598 13743 10728 13758
rect 10796 13743 11334 13758
rect 10598 13709 10627 13743
rect 10661 13709 10719 13743
rect 10796 13709 10811 13743
rect 10845 13709 10903 13743
rect 10937 13709 10995 13743
rect 11029 13709 11087 13743
rect 11121 13709 11179 13743
rect 11213 13709 11271 13743
rect 11305 13709 11334 13743
rect 11451 13715 11929 13789
rect 11986 13768 12382 13790
rect 11986 13734 12028 13768
rect 12062 13734 12382 13768
rect 11986 13718 12382 13734
rect 12506 13742 13232 13758
rect 10598 13696 10728 13709
rect 10796 13696 11334 13709
rect 10598 13678 11334 13696
rect 11855 13608 11929 13715
rect 12506 13680 12522 13742
rect 12590 13727 13232 13742
rect 12590 13693 12617 13727
rect 12651 13693 12709 13727
rect 12743 13693 12801 13727
rect 12835 13693 12893 13727
rect 12927 13693 12985 13727
rect 13019 13693 13077 13727
rect 13111 13693 13169 13727
rect 13203 13693 13232 13727
rect 12590 13680 13232 13693
rect 12506 13662 13232 13680
rect 12506 13660 12600 13662
rect 11410 13558 11759 13581
rect 11410 13524 11700 13558
rect 11734 13524 11759 13558
rect 11410 13507 11759 13524
rect 11855 13574 11878 13608
rect 11912 13574 11929 13608
rect 10722 13454 11274 13476
rect 10722 13445 10850 13454
rect 10918 13445 11274 13454
rect 10722 13411 10751 13445
rect 10785 13411 10843 13445
rect 10918 13411 10935 13445
rect 10969 13411 11027 13445
rect 11061 13411 11119 13445
rect 11153 13411 11211 13445
rect 11245 13411 11274 13445
rect 10722 13394 10850 13411
rect 10918 13394 11274 13411
rect 10722 13380 11274 13394
rect 10986 13342 11084 13348
rect 10986 13290 11006 13342
rect 11060 13290 11084 13342
rect 11410 13302 11484 13507
rect 11855 13493 11929 13574
rect 11660 13394 12210 13400
rect 11660 13382 12220 13394
rect 11660 13369 12002 13382
rect 12070 13369 12220 13382
rect 11660 13335 11689 13369
rect 11723 13335 11781 13369
rect 11815 13335 11873 13369
rect 11907 13335 11965 13369
rect 11999 13335 12002 13369
rect 12091 13335 12147 13369
rect 12181 13335 12220 13369
rect 11660 13320 12002 13335
rect 12070 13328 12220 13335
rect 12070 13320 12210 13328
rect 11660 13304 12210 13320
rect 10986 13272 11084 13290
rect 11198 13282 11484 13302
rect 11198 13244 11208 13282
rect 11246 13244 11484 13282
rect 11198 13228 11484 13244
rect 9414 13030 9422 13064
rect 9456 13030 9474 13064
rect 9414 13010 9474 13030
rect 9504 13066 9614 13080
rect 9504 13032 9542 13066
rect 9576 13032 9614 13066
rect 9504 13024 9614 13032
rect 10428 13064 10947 13089
rect 10428 13030 10860 13064
rect 10894 13030 10947 13064
rect 5856 12916 6408 12928
rect 5856 12897 5996 12916
rect 6064 12897 6408 12916
rect 5856 12863 5885 12897
rect 5919 12863 5977 12897
rect 6064 12863 6069 12897
rect 6103 12863 6161 12897
rect 6195 12863 6253 12897
rect 6287 12863 6345 12897
rect 6379 12863 6408 12897
rect 5856 12856 5996 12863
rect 6064 12856 6408 12863
rect 9538 12862 9569 13024
rect 10428 13011 10947 13030
rect 11042 13086 11124 13158
rect 11042 13032 11062 13086
rect 11114 13032 11124 13086
rect 5856 12832 6408 12856
rect 9244 12848 9980 12862
rect 9244 12831 9856 12848
rect 9928 12831 9980 12848
rect 9244 12797 9273 12831
rect 9307 12797 9365 12831
rect 9399 12797 9457 12831
rect 9491 12797 9549 12831
rect 9583 12797 9641 12831
rect 9675 12797 9733 12831
rect 9767 12797 9825 12831
rect 9951 12797 9980 12831
rect 9244 12782 9856 12797
rect 9928 12782 9980 12797
rect 9244 12766 9980 12782
rect 9342 12646 9894 12662
rect 9342 12631 9500 12646
rect 9574 12631 9894 12646
rect 9342 12597 9371 12631
rect 9405 12597 9463 12631
rect 9497 12597 9500 12631
rect 9589 12597 9647 12631
rect 9681 12597 9739 12631
rect 9773 12597 9831 12631
rect 9865 12597 9894 12631
rect 9342 12580 9500 12597
rect 9574 12580 9894 12597
rect 9342 12566 9894 12580
rect 5852 12432 6404 12452
rect 5852 12421 6280 12432
rect 6348 12421 6404 12432
rect 5852 12387 5881 12421
rect 5915 12387 5973 12421
rect 6007 12387 6065 12421
rect 6099 12387 6157 12421
rect 6191 12387 6249 12421
rect 6375 12387 6404 12421
rect 5852 12370 6280 12387
rect 6348 12370 6404 12387
rect 5852 12356 6404 12370
rect 9442 12342 9518 12368
rect 9642 12342 9692 12566
rect 9826 12394 9976 12408
rect 9826 12374 9872 12394
rect 9442 12302 9456 12342
rect 9498 12302 9518 12342
rect 9442 12286 9518 12302
rect 9634 12332 9702 12342
rect 9634 12292 9646 12332
rect 9688 12292 9702 12332
rect 9826 12340 9836 12374
rect 9826 12326 9872 12340
rect 9934 12326 9976 12394
rect 9826 12310 9976 12326
rect 6334 12208 6402 12218
rect 6334 12156 6340 12208
rect 6392 12156 6402 12208
rect 6334 12150 6402 12156
rect 4478 12100 5028 12114
rect 4478 12083 4906 12100
rect 4980 12083 5028 12100
rect 4478 12049 4507 12083
rect 4541 12049 4597 12083
rect 4631 12049 4689 12083
rect 4723 12049 4781 12083
rect 4815 12049 4873 12083
rect 4999 12049 5028 12083
rect 4478 12034 4906 12049
rect 4980 12034 5028 12049
rect 4478 12018 5028 12034
rect 5562 12112 6095 12121
rect 5562 12078 6018 12112
rect 6054 12078 6095 12112
rect 5562 12043 6095 12078
rect 6142 12118 6212 12126
rect 9456 12118 9508 12286
rect 9634 12280 9702 12292
rect 10428 12125 10506 13011
rect 11042 12974 11124 13032
rect 10722 12920 11274 12932
rect 10722 12901 10862 12920
rect 10930 12901 11274 12920
rect 10722 12867 10751 12901
rect 10785 12867 10843 12901
rect 10930 12867 10935 12901
rect 10969 12867 11027 12901
rect 11061 12867 11119 12901
rect 11153 12867 11211 12901
rect 11245 12867 11274 12901
rect 10722 12860 10862 12867
rect 10930 12860 11274 12867
rect 10722 12836 11274 12860
rect 10718 12436 11270 12456
rect 10718 12432 11146 12436
rect 10706 12425 11146 12432
rect 11214 12425 11270 12436
rect 10706 12391 10747 12425
rect 10781 12391 10839 12425
rect 10873 12391 10931 12425
rect 10965 12391 11023 12425
rect 11057 12391 11115 12425
rect 11241 12391 11270 12425
rect 10706 12374 11146 12391
rect 11214 12374 11270 12391
rect 10706 12366 11270 12374
rect 10718 12360 11270 12366
rect 11200 12212 11268 12222
rect 11200 12160 11206 12212
rect 11258 12160 11268 12212
rect 11200 12154 11268 12160
rect 6142 12066 6150 12118
rect 6202 12066 6212 12118
rect 6142 12060 6212 12066
rect 9342 12104 9894 12118
rect 9342 12087 9772 12104
rect 9846 12087 9894 12104
rect 9342 12053 9371 12087
rect 9405 12053 9463 12087
rect 9497 12053 9555 12087
rect 9589 12053 9647 12087
rect 9681 12053 9739 12087
rect 9865 12053 9894 12087
rect 4388 11820 5124 11838
rect 4388 11807 4560 11820
rect 4640 11807 5124 11820
rect 4388 11773 4417 11807
rect 4451 11773 4509 11807
rect 4543 11773 4560 11807
rect 4640 11773 4693 11807
rect 4727 11773 4785 11807
rect 4819 11773 4877 11807
rect 4911 11773 4969 11807
rect 5003 11773 5061 11807
rect 5095 11773 5124 11807
rect 4388 11756 4560 11773
rect 4640 11756 5124 11773
rect 4388 11742 5124 11756
rect 4558 11496 4618 11742
rect 5562 11670 5640 12043
rect 9342 12038 9772 12053
rect 9846 12038 9894 12053
rect 9342 12022 9894 12038
rect 10428 12116 10961 12125
rect 10428 12082 10884 12116
rect 10920 12082 10961 12116
rect 10428 12047 10961 12082
rect 11008 12122 11078 12130
rect 11008 12070 11016 12122
rect 11068 12070 11078 12122
rect 11008 12064 11078 12070
rect 5852 11892 6404 11908
rect 5852 11888 6002 11892
rect 5844 11877 6002 11888
rect 6070 11877 6404 11892
rect 5844 11843 5881 11877
rect 5915 11843 5973 11877
rect 6099 11843 6157 11877
rect 6191 11843 6249 11877
rect 6283 11843 6341 11877
rect 6375 11843 6404 11877
rect 5844 11830 6002 11843
rect 6070 11830 6404 11843
rect 5844 11822 6404 11830
rect 5852 11812 6404 11822
rect 9254 11824 9990 11842
rect 9254 11811 9426 11824
rect 9506 11811 9990 11824
rect 9254 11777 9283 11811
rect 9317 11777 9375 11811
rect 9409 11777 9426 11811
rect 9506 11777 9559 11811
rect 9593 11777 9651 11811
rect 9685 11777 9743 11811
rect 9777 11777 9835 11811
rect 9869 11777 9927 11811
rect 9961 11777 9990 11811
rect 9254 11760 9426 11777
rect 9506 11760 9990 11777
rect 9254 11746 9990 11760
rect 5042 11656 5640 11670
rect 5042 11622 5048 11656
rect 5084 11622 5640 11656
rect 5042 11592 5640 11622
rect 4558 11462 4566 11496
rect 4600 11462 4618 11496
rect 4558 11442 4618 11462
rect 4648 11498 4758 11512
rect 4648 11464 4686 11498
rect 4720 11464 4758 11498
rect 4648 11456 4758 11464
rect 9424 11500 9484 11746
rect 10428 11674 10506 12047
rect 10718 11898 11270 11912
rect 10714 11896 11270 11898
rect 10714 11881 10868 11896
rect 10936 11881 11270 11896
rect 10714 11847 10747 11881
rect 10781 11847 10839 11881
rect 10965 11847 11023 11881
rect 11057 11847 11115 11881
rect 11149 11847 11207 11881
rect 11241 11847 11270 11881
rect 10714 11834 10868 11847
rect 10936 11834 11270 11847
rect 10714 11832 11270 11834
rect 10718 11816 11270 11832
rect 9908 11660 10506 11674
rect 9908 11626 9914 11660
rect 9950 11626 10506 11660
rect 9908 11596 10506 11626
rect 9424 11466 9432 11500
rect 9466 11466 9484 11500
rect 4682 11294 4713 11456
rect 9424 11446 9484 11466
rect 9514 11502 9624 11516
rect 9514 11468 9552 11502
rect 9586 11468 9624 11502
rect 9514 11460 9624 11468
rect 9548 11298 9579 11460
rect 4388 11278 5124 11294
rect 4388 11263 4994 11278
rect 5074 11263 5124 11278
rect 4388 11229 4417 11263
rect 4451 11229 4509 11263
rect 4543 11229 4601 11263
rect 4635 11229 4693 11263
rect 4727 11229 4785 11263
rect 4819 11229 4877 11263
rect 4911 11229 4969 11263
rect 5095 11229 5124 11263
rect 4388 11214 4994 11229
rect 5074 11214 5124 11229
rect 4388 11198 5124 11214
rect 9254 11282 9990 11298
rect 9254 11267 9860 11282
rect 9940 11267 9990 11282
rect 9254 11233 9283 11267
rect 9317 11233 9375 11267
rect 9409 11233 9467 11267
rect 9501 11233 9559 11267
rect 9593 11233 9651 11267
rect 9685 11233 9743 11267
rect 9777 11233 9835 11267
rect 9961 11233 9990 11267
rect 9254 11218 9860 11233
rect 9940 11218 9990 11233
rect 9254 11202 9990 11218
rect 4486 11074 5038 11094
rect 4486 11063 4626 11074
rect 4706 11063 5038 11074
rect 4486 11029 4515 11063
rect 4549 11029 4607 11063
rect 4733 11029 4791 11063
rect 4825 11029 4883 11063
rect 4917 11029 4975 11063
rect 5009 11029 5038 11063
rect 4486 11010 4626 11029
rect 4706 11010 5038 11029
rect 4486 10998 5038 11010
rect 9352 11078 9904 11098
rect 9352 11067 9492 11078
rect 9572 11067 9904 11078
rect 9352 11033 9381 11067
rect 9415 11033 9473 11067
rect 9599 11033 9657 11067
rect 9691 11033 9749 11067
rect 9783 11033 9841 11067
rect 9875 11033 9904 11067
rect 9352 11014 9492 11033
rect 9572 11014 9904 11033
rect 9352 11002 9904 11014
rect 4586 10774 4662 10786
rect 4586 10734 4600 10774
rect 4642 10734 4662 10774
rect 4586 10718 4662 10734
rect 4776 10764 4848 10998
rect 4776 10730 4790 10764
rect 4778 10724 4790 10730
rect 4832 10730 4848 10764
rect 9452 10778 9528 10790
rect 4970 10732 5202 10762
rect 4970 10730 5054 10732
rect 4832 10724 4846 10730
rect 4606 10550 4656 10718
rect 4778 10708 4846 10724
rect 4970 10694 4982 10730
rect 5016 10694 5054 10730
rect 4970 10676 5054 10694
rect 5108 10676 5202 10732
rect 9452 10738 9466 10778
rect 9508 10738 9528 10778
rect 9452 10722 9528 10738
rect 9642 10768 9714 11002
rect 9642 10734 9656 10768
rect 9644 10728 9656 10734
rect 9698 10734 9714 10768
rect 9836 10736 10068 10766
rect 9836 10734 9920 10736
rect 9698 10728 9712 10734
rect 4970 10652 5202 10676
rect 9472 10554 9522 10722
rect 9644 10712 9712 10728
rect 9836 10698 9848 10734
rect 9882 10698 9920 10734
rect 9836 10680 9920 10698
rect 9974 10680 10068 10736
rect 9836 10656 10068 10680
rect 9644 10554 9712 10558
rect 4778 10550 4846 10554
rect 4486 10540 5038 10550
rect 4486 10519 4904 10540
rect 4984 10519 5038 10540
rect 4486 10485 4515 10519
rect 4549 10485 4607 10519
rect 4641 10485 4699 10519
rect 4733 10485 4791 10519
rect 4825 10485 4883 10519
rect 5009 10485 5038 10519
rect 4486 10476 4904 10485
rect 4984 10476 5038 10485
rect 4486 10454 5038 10476
rect 9352 10544 9904 10554
rect 9352 10523 9770 10544
rect 9850 10523 9904 10544
rect 9352 10489 9381 10523
rect 9415 10489 9473 10523
rect 9507 10489 9565 10523
rect 9599 10489 9657 10523
rect 9691 10489 9749 10523
rect 9875 10489 9904 10523
rect 9352 10480 9770 10489
rect 9850 10480 9904 10489
rect 9352 10458 9904 10480
rect 6112 6638 6470 6648
rect 6112 6617 6226 6638
rect 6282 6628 6470 6638
rect 6282 6617 6484 6628
rect 6112 6583 6141 6617
rect 6175 6583 6226 6617
rect 6282 6583 6325 6617
rect 6359 6583 6407 6617
rect 6441 6583 6484 6617
rect 6112 6580 6226 6583
rect 6282 6580 6484 6583
rect 6112 6562 6484 6580
rect 6112 6552 6470 6562
rect 6134 6390 6228 6398
rect 6134 6338 6168 6390
rect 6220 6338 6228 6390
rect 6262 6396 6328 6398
rect 6262 6344 6268 6396
rect 6320 6344 6328 6396
rect 6262 6338 6328 6344
rect 6134 6332 6228 6338
rect 6112 6088 6470 6104
rect 6112 6073 6170 6088
rect 6226 6073 6470 6088
rect 6112 6039 6141 6073
rect 6226 6039 6233 6073
rect 6267 6039 6325 6073
rect 6359 6039 6407 6073
rect 6441 6039 6470 6073
rect 6112 6030 6170 6039
rect 6226 6030 6470 6039
rect 6112 6008 6470 6030
rect 9928 6002 11490 6016
rect 9928 5985 10406 6002
rect 10464 6000 11490 6002
rect 10464 5985 10774 6000
rect 10832 5985 11490 6000
rect 9928 5951 9957 5985
rect 9991 5951 10047 5985
rect 10081 5951 10139 5985
rect 10173 5951 10231 5985
rect 10265 5951 10323 5985
rect 10357 5951 10406 5985
rect 10464 5951 10507 5985
rect 10541 5951 10599 5985
rect 10633 5951 10691 5985
rect 10725 5951 10774 5985
rect 10832 5951 10875 5985
rect 10909 5951 10967 5985
rect 11001 5951 11059 5985
rect 11093 5951 11151 5985
rect 11185 5951 11243 5985
rect 11277 5951 11335 5985
rect 11369 5951 11427 5985
rect 11461 5951 11490 5985
rect 9928 5940 10406 5951
rect 10464 5940 10774 5951
rect 9928 5936 10774 5940
rect 10832 5936 11490 5951
rect 9928 5920 11490 5936
rect 11988 5986 13552 6004
rect 13946 5996 15510 6012
rect 15942 6008 17504 6018
rect 11988 5973 12796 5986
rect 12852 5973 13552 5986
rect 11988 5939 12017 5973
rect 12051 5939 12109 5973
rect 12143 5939 12201 5973
rect 12235 5939 12293 5973
rect 12327 5939 12385 5973
rect 12419 5939 12477 5973
rect 12511 5939 12569 5973
rect 12603 5939 12661 5973
rect 12695 5939 12753 5973
rect 12787 5939 12796 5973
rect 12879 5939 12937 5973
rect 12971 5939 13029 5973
rect 13063 5939 13121 5973
rect 13155 5939 13213 5973
rect 13247 5939 13305 5973
rect 13339 5939 13397 5973
rect 13431 5939 13489 5973
rect 13523 5939 13552 5973
rect 11988 5928 12796 5939
rect 12852 5928 13552 5939
rect 13944 5994 15510 5996
rect 13944 5981 14754 5994
rect 14810 5981 15510 5994
rect 13944 5947 13975 5981
rect 14009 5947 14067 5981
rect 14101 5947 14159 5981
rect 14193 5947 14251 5981
rect 14285 5947 14343 5981
rect 14377 5947 14435 5981
rect 14469 5947 14527 5981
rect 14561 5947 14619 5981
rect 14653 5947 14711 5981
rect 14745 5947 14754 5981
rect 14837 5947 14895 5981
rect 14929 5947 14987 5981
rect 15021 5947 15079 5981
rect 15113 5947 15171 5981
rect 15205 5947 15263 5981
rect 15297 5947 15355 5981
rect 15389 5947 15447 5981
rect 15481 5947 15510 5981
rect 13944 5936 14754 5947
rect 14810 5936 15510 5947
rect 15938 6000 17504 6008
rect 15938 5987 16748 6000
rect 16804 5987 17504 6000
rect 15938 5953 15971 5987
rect 16005 5953 16061 5987
rect 16095 5953 16153 5987
rect 16187 5953 16245 5987
rect 16279 5953 16337 5987
rect 16371 5953 16429 5987
rect 16463 5953 16521 5987
rect 16555 5953 16613 5987
rect 16647 5953 16705 5987
rect 16739 5953 16748 5987
rect 16831 5953 16889 5987
rect 16923 5953 16981 5987
rect 17015 5953 17073 5987
rect 17107 5953 17165 5987
rect 17199 5953 17257 5987
rect 17291 5953 17349 5987
rect 17383 5953 17441 5987
rect 17475 5953 17504 5987
rect 15938 5942 16748 5953
rect 16804 5942 17504 5953
rect 13944 5930 15510 5936
rect 10214 5747 10272 5753
rect 10214 5713 10226 5747
rect 10260 5744 10272 5747
rect 10300 5744 10328 5920
rect 11988 5908 13552 5928
rect 13946 5916 15510 5930
rect 15942 5922 17504 5942
rect 10398 5815 10456 5821
rect 10398 5781 10410 5815
rect 10444 5812 10456 5815
rect 11138 5815 11196 5821
rect 11138 5812 11150 5815
rect 10444 5784 11150 5812
rect 10444 5781 10456 5784
rect 10398 5775 10456 5781
rect 11138 5781 11150 5784
rect 11184 5781 11196 5815
rect 11138 5775 11196 5781
rect 10582 5747 10640 5753
rect 10582 5744 10594 5747
rect 10260 5716 10594 5744
rect 10260 5713 10272 5716
rect 10214 5707 10272 5713
rect 10582 5713 10594 5716
rect 10628 5744 10640 5747
rect 10954 5747 11012 5753
rect 10954 5744 10966 5747
rect 10628 5716 10966 5744
rect 10628 5713 10640 5716
rect 10582 5707 10640 5713
rect 10954 5713 10966 5716
rect 11000 5744 11012 5747
rect 11230 5747 11288 5753
rect 11230 5744 11242 5747
rect 11000 5716 11242 5744
rect 11000 5713 11012 5716
rect 10954 5707 11012 5713
rect 11230 5713 11242 5716
rect 11276 5713 11288 5747
rect 11230 5707 11288 5713
rect 12276 5735 12334 5741
rect 12276 5701 12288 5735
rect 12322 5732 12334 5735
rect 12362 5732 12390 5908
rect 12460 5803 12518 5809
rect 12460 5769 12472 5803
rect 12506 5800 12518 5803
rect 13200 5803 13258 5809
rect 13200 5800 13212 5803
rect 12506 5772 13212 5800
rect 12506 5769 12518 5772
rect 12460 5763 12518 5769
rect 13200 5769 13212 5772
rect 13246 5769 13258 5803
rect 13200 5763 13258 5769
rect 14234 5743 14292 5749
rect 12644 5735 12702 5741
rect 12644 5732 12656 5735
rect 12322 5704 12656 5732
rect 12322 5701 12334 5704
rect 12276 5695 12334 5701
rect 12644 5701 12656 5704
rect 12690 5732 12702 5735
rect 13016 5735 13074 5741
rect 13016 5732 13028 5735
rect 12690 5704 13028 5732
rect 12690 5701 12702 5704
rect 12644 5695 12702 5701
rect 13016 5701 13028 5704
rect 13062 5732 13074 5735
rect 13292 5735 13350 5741
rect 13292 5732 13304 5735
rect 13062 5704 13304 5732
rect 13062 5701 13074 5704
rect 13016 5695 13074 5701
rect 13292 5701 13304 5704
rect 13338 5701 13350 5735
rect 14234 5709 14246 5743
rect 14280 5740 14292 5743
rect 14320 5740 14348 5916
rect 14418 5811 14476 5817
rect 14418 5777 14430 5811
rect 14464 5808 14476 5811
rect 15158 5811 15216 5817
rect 15158 5808 15170 5811
rect 14464 5780 15170 5808
rect 14464 5777 14476 5780
rect 14418 5771 14476 5777
rect 15158 5777 15170 5780
rect 15204 5777 15216 5811
rect 15158 5771 15216 5777
rect 16228 5749 16286 5755
rect 14602 5743 14660 5749
rect 14602 5740 14614 5743
rect 14280 5712 14614 5740
rect 14280 5709 14292 5712
rect 14234 5703 14292 5709
rect 14602 5709 14614 5712
rect 14648 5740 14660 5743
rect 14974 5743 15032 5749
rect 14974 5740 14986 5743
rect 14648 5712 14986 5740
rect 14648 5709 14660 5712
rect 14602 5703 14660 5709
rect 14974 5709 14986 5712
rect 15020 5740 15032 5743
rect 15250 5743 15308 5749
rect 15250 5740 15262 5743
rect 15020 5712 15262 5740
rect 15020 5709 15032 5712
rect 14974 5703 15032 5709
rect 15250 5709 15262 5712
rect 15296 5709 15308 5743
rect 16228 5715 16240 5749
rect 16274 5746 16286 5749
rect 16314 5746 16342 5922
rect 16412 5817 16470 5823
rect 16412 5783 16424 5817
rect 16458 5814 16470 5817
rect 17152 5817 17210 5823
rect 17152 5814 17164 5817
rect 16458 5786 17164 5814
rect 16458 5783 16470 5786
rect 16412 5777 16470 5783
rect 17152 5783 17164 5786
rect 17198 5783 17210 5817
rect 17152 5777 17210 5783
rect 16596 5749 16654 5755
rect 16596 5746 16608 5749
rect 16274 5718 16608 5746
rect 16274 5715 16286 5718
rect 16228 5709 16286 5715
rect 16596 5715 16608 5718
rect 16642 5746 16654 5749
rect 16968 5749 17026 5755
rect 16968 5746 16980 5749
rect 16642 5718 16980 5746
rect 16642 5715 16654 5718
rect 16596 5709 16654 5715
rect 16968 5715 16980 5718
rect 17014 5746 17026 5749
rect 17244 5749 17302 5755
rect 17244 5746 17256 5749
rect 17014 5718 17256 5746
rect 17014 5715 17026 5718
rect 16968 5709 17026 5715
rect 17244 5715 17256 5718
rect 17290 5715 17302 5749
rect 17244 5709 17302 5715
rect 15250 5703 15308 5709
rect 13292 5695 13350 5701
rect 10306 5679 10364 5685
rect 10306 5645 10318 5679
rect 10352 5676 10364 5679
rect 10766 5679 10824 5685
rect 10766 5676 10778 5679
rect 10352 5648 10778 5676
rect 10352 5645 10364 5648
rect 10306 5639 10364 5645
rect 10766 5645 10778 5648
rect 10812 5676 10824 5679
rect 11138 5679 11196 5685
rect 16320 5681 16378 5687
rect 11138 5676 11150 5679
rect 10812 5648 11150 5676
rect 10812 5645 10824 5648
rect 10766 5639 10824 5645
rect 10404 5618 10470 5620
rect 1746 5590 3308 5596
rect 1736 5578 3308 5590
rect 1736 5565 2564 5578
rect 2620 5565 3308 5578
rect 1736 5531 1775 5565
rect 1809 5531 1865 5565
rect 1899 5531 1957 5565
rect 1991 5531 2049 5565
rect 2083 5531 2141 5565
rect 2175 5531 2233 5565
rect 2267 5531 2325 5565
rect 2359 5531 2417 5565
rect 2451 5531 2509 5565
rect 2543 5531 2564 5565
rect 2635 5531 2693 5565
rect 2727 5531 2785 5565
rect 2819 5531 2877 5565
rect 2911 5531 2969 5565
rect 3003 5531 3061 5565
rect 3095 5531 3153 5565
rect 3187 5531 3245 5565
rect 3279 5531 3308 5565
rect 1736 5524 2564 5531
rect 1746 5520 2564 5524
rect 2620 5520 3308 5531
rect 1746 5500 3308 5520
rect 3880 5570 5442 5588
rect 3880 5557 4686 5570
rect 4742 5557 5442 5570
rect 3880 5523 3909 5557
rect 3943 5523 3999 5557
rect 4033 5523 4091 5557
rect 4125 5523 4183 5557
rect 4217 5523 4275 5557
rect 4309 5523 4367 5557
rect 4401 5523 4459 5557
rect 4493 5523 4551 5557
rect 4585 5523 4643 5557
rect 4677 5523 4686 5557
rect 4769 5523 4827 5557
rect 4861 5523 4919 5557
rect 4953 5523 5011 5557
rect 5045 5523 5103 5557
rect 5137 5523 5195 5557
rect 5229 5523 5287 5557
rect 5321 5523 5379 5557
rect 5413 5523 5442 5557
rect 3880 5512 4686 5523
rect 4742 5512 5442 5523
rect 2032 5327 2090 5333
rect 2032 5293 2044 5327
rect 2078 5324 2090 5327
rect 2118 5324 2146 5500
rect 3880 5492 5442 5512
rect 5830 5570 7394 5588
rect 5830 5557 6638 5570
rect 6694 5557 7394 5570
rect 5830 5523 5859 5557
rect 5893 5523 5951 5557
rect 5985 5523 6043 5557
rect 6077 5523 6135 5557
rect 6169 5523 6227 5557
rect 6261 5523 6319 5557
rect 6353 5523 6411 5557
rect 6445 5523 6503 5557
rect 6537 5523 6595 5557
rect 6629 5523 6638 5557
rect 6721 5523 6779 5557
rect 6813 5523 6871 5557
rect 6905 5523 6963 5557
rect 6997 5523 7055 5557
rect 7089 5523 7147 5557
rect 7181 5523 7239 5557
rect 7273 5523 7331 5557
rect 7365 5523 7394 5557
rect 5830 5512 6638 5523
rect 6694 5512 7394 5523
rect 5830 5492 7394 5512
rect 7832 5576 9396 5594
rect 7832 5563 8640 5576
rect 8696 5563 9396 5576
rect 7832 5529 7861 5563
rect 7895 5529 7953 5563
rect 7987 5529 8045 5563
rect 8079 5529 8137 5563
rect 8171 5529 8229 5563
rect 8263 5529 8321 5563
rect 8355 5529 8413 5563
rect 8447 5529 8505 5563
rect 8539 5529 8597 5563
rect 8631 5529 8640 5563
rect 8723 5529 8781 5563
rect 8815 5529 8873 5563
rect 8907 5529 8965 5563
rect 8999 5529 9057 5563
rect 9091 5529 9149 5563
rect 9183 5529 9241 5563
rect 9275 5529 9333 5563
rect 9367 5529 9396 5563
rect 10404 5566 10410 5618
rect 10462 5566 10470 5618
rect 10404 5562 10470 5566
rect 7832 5518 8640 5529
rect 8696 5518 9396 5529
rect 7832 5498 9396 5518
rect 2216 5395 2274 5401
rect 2216 5361 2228 5395
rect 2262 5392 2274 5395
rect 2956 5395 3014 5401
rect 2956 5392 2968 5395
rect 2262 5364 2968 5392
rect 2262 5361 2274 5364
rect 2216 5355 2274 5361
rect 2956 5361 2968 5364
rect 3002 5361 3014 5395
rect 2956 5355 3014 5361
rect 2400 5327 2458 5333
rect 2400 5324 2412 5327
rect 2078 5296 2412 5324
rect 2078 5293 2090 5296
rect 2032 5287 2090 5293
rect 2400 5293 2412 5296
rect 2446 5324 2458 5327
rect 2772 5327 2830 5333
rect 2772 5324 2784 5327
rect 2446 5296 2784 5324
rect 2446 5293 2458 5296
rect 2400 5287 2458 5293
rect 2772 5293 2784 5296
rect 2818 5324 2830 5327
rect 3048 5327 3106 5333
rect 3048 5324 3060 5327
rect 2818 5296 3060 5324
rect 2818 5293 2830 5296
rect 2772 5287 2830 5293
rect 3048 5293 3060 5296
rect 3094 5293 3106 5327
rect 3048 5287 3106 5293
rect 4166 5319 4224 5325
rect 4166 5285 4178 5319
rect 4212 5316 4224 5319
rect 4252 5316 4280 5492
rect 4350 5387 4408 5393
rect 4350 5353 4362 5387
rect 4396 5384 4408 5387
rect 5090 5387 5148 5393
rect 5090 5384 5102 5387
rect 4396 5356 5102 5384
rect 4396 5353 4408 5356
rect 4350 5347 4408 5353
rect 5090 5353 5102 5356
rect 5136 5353 5148 5387
rect 5090 5347 5148 5353
rect 4534 5319 4592 5325
rect 4534 5316 4546 5319
rect 4212 5288 4546 5316
rect 4212 5285 4224 5288
rect 4166 5279 4224 5285
rect 4534 5285 4546 5288
rect 4580 5316 4592 5319
rect 4906 5319 4964 5325
rect 4906 5316 4918 5319
rect 4580 5288 4918 5316
rect 4580 5285 4592 5288
rect 4534 5279 4592 5285
rect 4906 5285 4918 5288
rect 4952 5316 4964 5319
rect 5182 5319 5240 5325
rect 5182 5316 5194 5319
rect 4952 5288 5194 5316
rect 4952 5285 4964 5288
rect 4906 5279 4964 5285
rect 5182 5285 5194 5288
rect 5228 5285 5240 5319
rect 5182 5279 5240 5285
rect 6118 5319 6176 5325
rect 6118 5285 6130 5319
rect 6164 5316 6176 5319
rect 6204 5316 6232 5492
rect 6302 5387 6360 5393
rect 6302 5353 6314 5387
rect 6348 5384 6360 5387
rect 7042 5387 7100 5393
rect 7042 5384 7054 5387
rect 6348 5356 7054 5384
rect 6348 5353 6360 5356
rect 6302 5347 6360 5353
rect 7042 5353 7054 5356
rect 7088 5353 7100 5387
rect 7042 5347 7100 5353
rect 8120 5325 8178 5331
rect 6486 5319 6544 5325
rect 6486 5316 6498 5319
rect 6164 5288 6498 5316
rect 6164 5285 6176 5288
rect 6118 5279 6176 5285
rect 6486 5285 6498 5288
rect 6532 5316 6544 5319
rect 6858 5319 6916 5325
rect 6858 5316 6870 5319
rect 6532 5288 6870 5316
rect 6532 5285 6544 5288
rect 6486 5279 6544 5285
rect 6858 5285 6870 5288
rect 6904 5316 6916 5319
rect 7134 5319 7192 5325
rect 7134 5316 7146 5319
rect 6904 5288 7146 5316
rect 6904 5285 6916 5288
rect 6858 5279 6916 5285
rect 7134 5285 7146 5288
rect 7180 5285 7192 5319
rect 8120 5291 8132 5325
rect 8166 5322 8178 5325
rect 8206 5322 8234 5498
rect 10860 5472 10888 5648
rect 11138 5645 11150 5648
rect 11184 5645 11196 5679
rect 14326 5675 14384 5681
rect 11138 5639 11196 5645
rect 12368 5667 12426 5673
rect 12368 5633 12380 5667
rect 12414 5664 12426 5667
rect 12828 5667 12886 5673
rect 12828 5664 12840 5667
rect 12414 5636 12840 5664
rect 12414 5633 12426 5636
rect 11412 5606 11472 5630
rect 12368 5627 12426 5633
rect 12828 5633 12840 5636
rect 12874 5664 12886 5667
rect 13200 5667 13258 5673
rect 13200 5664 13212 5667
rect 12874 5636 13212 5664
rect 12874 5633 12886 5636
rect 12828 5627 12886 5633
rect 11412 5570 11426 5606
rect 11466 5604 11472 5606
rect 11466 5596 11818 5604
rect 12464 5600 12524 5606
rect 12464 5596 12478 5600
rect 11466 5570 12478 5596
rect 11412 5566 12478 5570
rect 12512 5566 12524 5600
rect 11412 5554 11472 5566
rect 11804 5562 12524 5566
rect 11896 5558 12524 5562
rect 12464 5544 12524 5558
rect 9928 5452 11490 5472
rect 12922 5460 12950 5636
rect 13200 5633 13212 5636
rect 13246 5633 13258 5667
rect 14326 5641 14338 5675
rect 14372 5672 14384 5675
rect 14786 5675 14844 5681
rect 14786 5672 14798 5675
rect 14372 5644 14798 5672
rect 14372 5641 14384 5644
rect 14326 5635 14384 5641
rect 14786 5641 14798 5644
rect 14832 5672 14844 5675
rect 15158 5675 15216 5681
rect 15158 5672 15170 5675
rect 14832 5644 15170 5672
rect 14832 5641 14844 5644
rect 14786 5635 14844 5641
rect 13200 5627 13258 5633
rect 13482 5594 13534 5612
rect 14422 5608 14482 5614
rect 14422 5604 14436 5608
rect 13565 5594 14436 5604
rect 13480 5558 13494 5594
rect 13528 5574 14436 5594
rect 14470 5574 14482 5608
rect 13528 5566 14482 5574
rect 13528 5558 13588 5566
rect 13480 5556 13588 5558
rect 13482 5546 13534 5556
rect 14422 5552 14482 5566
rect 14880 5468 14908 5644
rect 15158 5641 15170 5644
rect 15204 5641 15216 5675
rect 16320 5647 16332 5681
rect 16366 5678 16378 5681
rect 16780 5681 16838 5687
rect 16780 5678 16792 5681
rect 16366 5650 16792 5678
rect 16366 5647 16378 5650
rect 16320 5641 16378 5647
rect 16780 5647 16792 5650
rect 16826 5678 16838 5681
rect 17152 5681 17210 5687
rect 17152 5678 17164 5681
rect 16826 5650 17164 5678
rect 16826 5647 16838 5650
rect 16780 5641 16838 5647
rect 15158 5635 15216 5641
rect 15440 5602 15492 5620
rect 16416 5614 16476 5620
rect 16416 5610 16430 5614
rect 15848 5606 16430 5610
rect 15524 5602 16430 5606
rect 15438 5566 15452 5602
rect 15486 5580 16430 5602
rect 16464 5580 16476 5614
rect 15486 5572 16476 5580
rect 15486 5566 15884 5572
rect 15438 5564 15884 5566
rect 15440 5554 15492 5564
rect 16416 5558 16476 5572
rect 16874 5474 16902 5650
rect 17152 5647 17164 5650
rect 17198 5647 17210 5681
rect 17152 5641 17210 5647
rect 17434 5608 17486 5626
rect 17432 5572 17446 5608
rect 17480 5596 17540 5608
rect 17480 5572 17822 5596
rect 17432 5570 17822 5572
rect 17434 5564 17822 5570
rect 17434 5560 17514 5564
rect 9928 5441 11214 5452
rect 11270 5441 11490 5452
rect 9928 5407 9957 5441
rect 9991 5407 10047 5441
rect 10081 5407 10139 5441
rect 10173 5407 10231 5441
rect 10265 5407 10323 5441
rect 10357 5407 10415 5441
rect 10449 5407 10507 5441
rect 10541 5407 10599 5441
rect 10633 5407 10691 5441
rect 10725 5407 10783 5441
rect 10817 5407 10875 5441
rect 10909 5407 10967 5441
rect 11001 5407 11059 5441
rect 11093 5407 11151 5441
rect 11185 5407 11214 5441
rect 11277 5407 11335 5441
rect 11369 5407 11427 5441
rect 11461 5407 11490 5441
rect 8304 5393 8362 5399
rect 8304 5359 8316 5393
rect 8350 5390 8362 5393
rect 9044 5393 9102 5399
rect 9044 5390 9056 5393
rect 8350 5362 9056 5390
rect 8350 5359 8362 5362
rect 8304 5353 8362 5359
rect 9044 5359 9056 5362
rect 9090 5359 9102 5393
rect 9928 5394 11214 5407
rect 11270 5394 11490 5407
rect 9928 5376 11490 5394
rect 11988 5440 13552 5460
rect 11988 5429 12800 5440
rect 12856 5429 13552 5440
rect 11988 5395 12017 5429
rect 12051 5395 12109 5429
rect 12143 5395 12201 5429
rect 12235 5395 12293 5429
rect 12327 5395 12385 5429
rect 12419 5395 12477 5429
rect 12511 5395 12569 5429
rect 12603 5395 12661 5429
rect 12695 5395 12753 5429
rect 12787 5395 12800 5429
rect 12879 5395 12937 5429
rect 12971 5395 13029 5429
rect 13063 5395 13121 5429
rect 13155 5395 13213 5429
rect 13247 5395 13305 5429
rect 13339 5395 13397 5429
rect 13431 5395 13489 5429
rect 13523 5395 13552 5429
rect 11988 5382 12800 5395
rect 12856 5382 13552 5395
rect 11988 5364 13552 5382
rect 13946 5448 15510 5468
rect 13946 5437 14758 5448
rect 14814 5437 15510 5448
rect 13946 5403 13975 5437
rect 14009 5403 14067 5437
rect 14101 5403 14159 5437
rect 14193 5403 14251 5437
rect 14285 5403 14343 5437
rect 14377 5403 14435 5437
rect 14469 5403 14527 5437
rect 14561 5403 14619 5437
rect 14653 5403 14711 5437
rect 14745 5403 14758 5437
rect 14837 5403 14895 5437
rect 14929 5403 14987 5437
rect 15021 5403 15079 5437
rect 15113 5403 15171 5437
rect 15205 5403 15263 5437
rect 15297 5403 15355 5437
rect 15389 5403 15447 5437
rect 15481 5403 15510 5437
rect 13946 5390 14758 5403
rect 14814 5390 15510 5403
rect 13946 5372 15510 5390
rect 15942 5454 17504 5474
rect 15942 5443 16752 5454
rect 16808 5443 17504 5454
rect 15942 5409 15971 5443
rect 16005 5409 16061 5443
rect 16095 5409 16153 5443
rect 16187 5409 16245 5443
rect 16279 5409 16337 5443
rect 16371 5409 16429 5443
rect 16463 5409 16521 5443
rect 16555 5409 16613 5443
rect 16647 5409 16705 5443
rect 16739 5409 16752 5443
rect 16831 5409 16889 5443
rect 16923 5409 16981 5443
rect 17015 5409 17073 5443
rect 17107 5409 17165 5443
rect 17199 5409 17257 5443
rect 17291 5409 17349 5443
rect 17383 5409 17441 5443
rect 17475 5409 17504 5443
rect 15942 5396 16752 5409
rect 16808 5396 17504 5409
rect 15942 5378 17504 5396
rect 9044 5353 9102 5359
rect 8488 5325 8546 5331
rect 8488 5322 8500 5325
rect 8166 5294 8500 5322
rect 8166 5291 8178 5294
rect 8120 5285 8178 5291
rect 8488 5291 8500 5294
rect 8534 5322 8546 5325
rect 8860 5325 8918 5331
rect 8860 5322 8872 5325
rect 8534 5294 8872 5322
rect 8534 5291 8546 5294
rect 8488 5285 8546 5291
rect 8860 5291 8872 5294
rect 8906 5322 8918 5325
rect 9136 5325 9194 5331
rect 9136 5322 9148 5325
rect 8906 5294 9148 5322
rect 8906 5291 8918 5294
rect 8860 5285 8918 5291
rect 9136 5291 9148 5294
rect 9182 5291 9194 5325
rect 9136 5285 9194 5291
rect 17790 5302 17822 5564
rect 18302 5440 19222 5444
rect 18302 5428 19226 5440
rect 18302 5413 18726 5428
rect 18784 5413 19226 5428
rect 18302 5379 18331 5413
rect 18365 5379 18423 5413
rect 18457 5379 18515 5413
rect 18549 5379 18607 5413
rect 18641 5379 18699 5413
rect 18784 5379 18791 5413
rect 18825 5379 18883 5413
rect 18917 5379 18975 5413
rect 19009 5379 19067 5413
rect 19101 5379 19159 5413
rect 19193 5379 19226 5413
rect 18302 5364 18726 5379
rect 18784 5374 19226 5379
rect 18784 5364 19222 5374
rect 18302 5348 19222 5364
rect 7134 5279 7192 5285
rect 17790 5270 18732 5302
rect 2124 5259 2182 5265
rect 2124 5225 2136 5259
rect 2170 5256 2182 5259
rect 2584 5259 2642 5265
rect 2584 5256 2596 5259
rect 2170 5228 2596 5256
rect 2170 5225 2182 5228
rect 2124 5219 2182 5225
rect 2584 5225 2596 5228
rect 2630 5256 2642 5259
rect 2956 5259 3014 5265
rect 2956 5256 2968 5259
rect 2630 5228 2968 5256
rect 2630 5225 2642 5228
rect 2584 5219 2642 5225
rect 2222 5198 2288 5200
rect 2222 5146 2228 5198
rect 2280 5146 2288 5198
rect 2222 5142 2288 5146
rect 2678 5052 2706 5228
rect 2956 5225 2968 5228
rect 3002 5225 3014 5259
rect 8212 5257 8270 5263
rect 2956 5219 3014 5225
rect 4258 5251 4316 5257
rect 4258 5217 4270 5251
rect 4304 5248 4316 5251
rect 4718 5251 4776 5257
rect 4718 5248 4730 5251
rect 4304 5220 4730 5248
rect 4304 5217 4316 5220
rect 4258 5211 4316 5217
rect 4718 5217 4730 5220
rect 4764 5248 4776 5251
rect 5090 5251 5148 5257
rect 5090 5248 5102 5251
rect 4764 5220 5102 5248
rect 4764 5217 4776 5220
rect 4718 5211 4776 5217
rect 3230 5186 3290 5210
rect 3230 5150 3244 5186
rect 3284 5184 3290 5186
rect 4354 5184 4414 5190
rect 3284 5180 3837 5184
rect 4354 5180 4368 5184
rect 3284 5150 4368 5180
rect 4402 5150 4414 5184
rect 3230 5146 4414 5150
rect 3230 5134 3290 5146
rect 3636 5142 4414 5146
rect 4354 5128 4414 5142
rect 1746 5040 3308 5052
rect 4812 5044 4840 5220
rect 5090 5217 5102 5220
rect 5136 5217 5148 5251
rect 5090 5211 5148 5217
rect 6210 5251 6268 5257
rect 6210 5217 6222 5251
rect 6256 5248 6268 5251
rect 6670 5251 6728 5257
rect 6670 5248 6682 5251
rect 6256 5220 6682 5248
rect 6256 5217 6268 5220
rect 6210 5211 6268 5217
rect 6670 5217 6682 5220
rect 6716 5248 6728 5251
rect 7042 5251 7100 5257
rect 7042 5248 7054 5251
rect 6716 5220 7054 5248
rect 6716 5217 6728 5220
rect 6670 5211 6728 5217
rect 5372 5178 5424 5196
rect 6306 5184 6366 5190
rect 6306 5180 6320 5184
rect 5612 5178 6320 5180
rect 5370 5142 5384 5178
rect 5418 5150 6320 5178
rect 6354 5150 6366 5184
rect 5418 5142 6366 5150
rect 5370 5140 5659 5142
rect 5372 5130 5424 5140
rect 6306 5128 6366 5142
rect 6764 5044 6792 5220
rect 7042 5217 7054 5220
rect 7088 5217 7100 5251
rect 8212 5223 8224 5257
rect 8258 5254 8270 5257
rect 8672 5257 8730 5263
rect 8672 5254 8684 5257
rect 8258 5226 8684 5254
rect 8258 5223 8270 5226
rect 8212 5217 8270 5223
rect 8672 5223 8684 5226
rect 8718 5254 8730 5257
rect 9044 5257 9102 5263
rect 9044 5254 9056 5257
rect 8718 5226 9056 5254
rect 8718 5223 8730 5226
rect 8672 5217 8730 5223
rect 7042 5211 7100 5217
rect 7324 5178 7376 5196
rect 8308 5190 8368 5196
rect 8308 5186 8322 5190
rect 7550 5178 8322 5186
rect 7322 5142 7336 5178
rect 7370 5156 8322 5178
rect 8356 5156 8368 5190
rect 7370 5148 8368 5156
rect 7370 5142 7611 5148
rect 7322 5140 7611 5142
rect 7324 5130 7376 5140
rect 8308 5134 8368 5148
rect 8766 5050 8794 5226
rect 9044 5223 9056 5226
rect 9090 5223 9102 5257
rect 9044 5217 9102 5223
rect 9906 5210 17524 5242
rect 9326 5184 9378 5202
rect 9906 5184 9938 5210
rect 9324 5148 9338 5184
rect 9372 5148 9938 5184
rect 9324 5146 9938 5148
rect 9326 5136 9378 5146
rect 9762 5144 9938 5146
rect 17492 5146 17524 5210
rect 18598 5222 18648 5242
rect 18598 5188 18608 5222
rect 18642 5188 18648 5222
rect 10046 5138 11610 5142
rect 10046 5120 11614 5138
rect 10046 5111 10188 5120
rect 10244 5111 11614 5120
rect 17492 5114 18178 5146
rect 18598 5134 18648 5188
rect 18678 5194 18732 5270
rect 18678 5160 18690 5194
rect 18724 5160 18732 5194
rect 10046 5077 10075 5111
rect 10109 5077 10167 5111
rect 10244 5077 10259 5111
rect 10293 5077 10351 5111
rect 10385 5077 10443 5111
rect 10477 5077 10535 5111
rect 10569 5077 10627 5111
rect 10661 5077 10719 5111
rect 10753 5077 10811 5111
rect 10845 5077 10903 5111
rect 10937 5077 10995 5111
rect 11029 5077 11087 5111
rect 11121 5077 11179 5111
rect 11213 5077 11271 5111
rect 11305 5077 11363 5111
rect 11397 5077 11455 5111
rect 11489 5077 11547 5111
rect 11581 5077 11614 5111
rect 18146 5102 18178 5114
rect 18426 5108 18480 5120
rect 18250 5102 18432 5108
rect 10046 5062 10188 5077
rect 10244 5072 11614 5077
rect 12228 5080 13788 5098
rect 10244 5062 11610 5072
rect 1746 5021 2584 5040
rect 2640 5021 3308 5040
rect 1746 4987 1775 5021
rect 1809 4987 1865 5021
rect 1899 4987 1957 5021
rect 1991 4987 2049 5021
rect 2083 4987 2141 5021
rect 2175 4987 2233 5021
rect 2267 4987 2325 5021
rect 2359 4987 2417 5021
rect 2451 4987 2509 5021
rect 2543 4987 2584 5021
rect 2640 4987 2693 5021
rect 2727 4987 2785 5021
rect 2819 4987 2877 5021
rect 2911 4987 2969 5021
rect 3003 4987 3061 5021
rect 3095 4987 3153 5021
rect 3187 4987 3245 5021
rect 3279 4987 3308 5021
rect 1746 4982 2584 4987
rect 2640 4982 3308 4987
rect 1746 4956 3308 4982
rect 3880 5024 5442 5044
rect 3880 5013 4690 5024
rect 4746 5013 5442 5024
rect 3880 4979 3909 5013
rect 3943 4979 3999 5013
rect 4033 4979 4091 5013
rect 4125 4979 4183 5013
rect 4217 4979 4275 5013
rect 4309 4979 4367 5013
rect 4401 4979 4459 5013
rect 4493 4979 4551 5013
rect 4585 4979 4643 5013
rect 4677 4979 4690 5013
rect 4769 4979 4827 5013
rect 4861 4979 4919 5013
rect 4953 4979 5011 5013
rect 5045 4979 5103 5013
rect 5137 4979 5195 5013
rect 5229 4979 5287 5013
rect 5321 4979 5379 5013
rect 5413 4979 5442 5013
rect 3880 4966 4690 4979
rect 4746 4966 5442 4979
rect 3880 4948 5442 4966
rect 5830 5024 7394 5044
rect 5830 5013 6642 5024
rect 6698 5013 7394 5024
rect 5830 4979 5859 5013
rect 5893 4979 5951 5013
rect 5985 4979 6043 5013
rect 6077 4979 6135 5013
rect 6169 4979 6227 5013
rect 6261 4979 6319 5013
rect 6353 4979 6411 5013
rect 6445 4979 6503 5013
rect 6537 4979 6595 5013
rect 6629 4979 6642 5013
rect 6721 4979 6779 5013
rect 6813 4979 6871 5013
rect 6905 4979 6963 5013
rect 6997 4979 7055 5013
rect 7089 4979 7147 5013
rect 7181 4979 7239 5013
rect 7273 4979 7331 5013
rect 7365 4979 7394 5013
rect 5830 4966 6642 4979
rect 6698 4966 7394 4979
rect 5830 4948 7394 4966
rect 7832 5030 9396 5050
rect 10046 5046 11610 5062
rect 12228 5067 13032 5080
rect 13088 5067 13788 5080
rect 7832 5019 8644 5030
rect 8700 5019 9396 5030
rect 7832 4985 7861 5019
rect 7895 4985 7953 5019
rect 7987 4985 8045 5019
rect 8079 4985 8137 5019
rect 8171 4985 8229 5019
rect 8263 4985 8321 5019
rect 8355 4985 8413 5019
rect 8447 4985 8505 5019
rect 8539 4985 8597 5019
rect 8631 4985 8644 5019
rect 8723 4985 8781 5019
rect 8815 4985 8873 5019
rect 8907 4985 8965 5019
rect 8999 4985 9057 5019
rect 9091 4985 9149 5019
rect 9183 4985 9241 5019
rect 9275 4985 9333 5019
rect 9367 4985 9396 5019
rect 7832 4972 8644 4985
rect 8700 4972 9396 4985
rect 7832 4954 9396 4972
rect 10242 4873 10300 4879
rect 10242 4839 10254 4873
rect 10288 4870 10300 4873
rect 10328 4870 10356 5046
rect 12228 5033 12257 5067
rect 12291 5033 12345 5067
rect 12379 5033 12437 5067
rect 12471 5033 12529 5067
rect 12563 5033 12621 5067
rect 12655 5033 12713 5067
rect 12747 5033 12805 5067
rect 12839 5033 12897 5067
rect 12931 5033 12989 5067
rect 13023 5033 13032 5067
rect 13115 5033 13173 5067
rect 13207 5033 13265 5067
rect 13299 5033 13357 5067
rect 13391 5033 13449 5067
rect 13483 5033 13541 5067
rect 13575 5033 13633 5067
rect 13667 5033 13725 5067
rect 13759 5033 13788 5067
rect 12228 5022 13032 5033
rect 13088 5022 13788 5033
rect 12228 5002 13788 5022
rect 14228 5074 15790 5092
rect 14228 5061 15034 5074
rect 15090 5061 15790 5074
rect 14228 5027 14257 5061
rect 14291 5027 14347 5061
rect 14381 5027 14439 5061
rect 14473 5027 14531 5061
rect 14565 5027 14623 5061
rect 14657 5027 14715 5061
rect 14749 5027 14807 5061
rect 14841 5027 14899 5061
rect 14933 5027 14991 5061
rect 15025 5027 15034 5061
rect 15117 5027 15175 5061
rect 15209 5027 15267 5061
rect 15301 5027 15359 5061
rect 15393 5027 15451 5061
rect 15485 5027 15543 5061
rect 15577 5027 15635 5061
rect 15669 5027 15727 5061
rect 15761 5027 15790 5061
rect 14228 5016 15034 5027
rect 15090 5016 15790 5027
rect 10426 4941 10484 4947
rect 10426 4907 10438 4941
rect 10472 4938 10484 4941
rect 11166 4941 11224 4947
rect 11166 4938 11178 4941
rect 10472 4910 11178 4938
rect 10472 4907 10484 4910
rect 10426 4901 10484 4907
rect 11166 4907 11178 4910
rect 11212 4907 11224 4941
rect 11166 4901 11224 4907
rect 10610 4873 10668 4879
rect 10610 4870 10622 4873
rect 10288 4842 10622 4870
rect 10288 4839 10300 4842
rect 10242 4833 10300 4839
rect 10610 4839 10622 4842
rect 10656 4870 10668 4873
rect 10982 4873 11040 4879
rect 10982 4870 10994 4873
rect 10656 4842 10994 4870
rect 10656 4839 10668 4842
rect 10610 4833 10668 4839
rect 10982 4839 10994 4842
rect 11028 4870 11040 4873
rect 11258 4873 11316 4879
rect 11258 4870 11270 4873
rect 11028 4842 11270 4870
rect 11028 4839 11040 4842
rect 10982 4833 11040 4839
rect 11258 4839 11270 4842
rect 11304 4839 11316 4873
rect 11258 4833 11316 4839
rect 12512 4829 12570 4835
rect 10334 4805 10392 4811
rect 10334 4771 10346 4805
rect 10380 4802 10392 4805
rect 10794 4805 10852 4811
rect 10794 4802 10806 4805
rect 10380 4774 10806 4802
rect 10380 4771 10392 4774
rect 10334 4765 10392 4771
rect 10794 4771 10806 4774
rect 10840 4802 10852 4805
rect 11166 4805 11224 4811
rect 11166 4802 11178 4805
rect 10840 4774 11178 4802
rect 10840 4771 10852 4774
rect 10794 4765 10852 4771
rect 10432 4744 10498 4746
rect 10432 4692 10438 4744
rect 10490 4692 10498 4744
rect 10432 4688 10498 4692
rect 10888 4598 10916 4774
rect 11166 4771 11178 4774
rect 11212 4771 11224 4805
rect 12512 4795 12524 4829
rect 12558 4826 12570 4829
rect 12598 4826 12626 5002
rect 14228 4996 15790 5016
rect 16252 5056 17812 5074
rect 18146 5070 18432 5102
rect 18470 5070 18572 5108
rect 16252 5043 17056 5056
rect 17112 5043 17812 5056
rect 18426 5054 18480 5070
rect 16252 5009 16281 5043
rect 16315 5009 16369 5043
rect 16403 5009 16461 5043
rect 16495 5009 16553 5043
rect 16587 5009 16645 5043
rect 16679 5009 16737 5043
rect 16771 5009 16829 5043
rect 16863 5009 16921 5043
rect 16955 5009 17013 5043
rect 17047 5009 17056 5043
rect 17139 5009 17197 5043
rect 17231 5009 17289 5043
rect 17323 5009 17381 5043
rect 17415 5009 17473 5043
rect 17507 5009 17565 5043
rect 17599 5009 17657 5043
rect 17691 5009 17749 5043
rect 17783 5009 17812 5043
rect 18608 5024 18640 5134
rect 18678 5114 18732 5160
rect 18678 5110 18716 5114
rect 18250 5023 18640 5024
rect 16252 4998 17056 5009
rect 17112 4998 17812 5009
rect 12696 4897 12754 4903
rect 12696 4863 12708 4897
rect 12742 4894 12754 4897
rect 13436 4897 13494 4903
rect 13436 4894 13448 4897
rect 12742 4866 13448 4894
rect 12742 4863 12754 4866
rect 12696 4857 12754 4863
rect 13436 4863 13448 4866
rect 13482 4863 13494 4897
rect 13436 4857 13494 4863
rect 12880 4829 12938 4835
rect 12880 4826 12892 4829
rect 12558 4798 12892 4826
rect 12558 4795 12570 4798
rect 12512 4789 12570 4795
rect 12880 4795 12892 4798
rect 12926 4826 12938 4829
rect 13252 4829 13310 4835
rect 13252 4826 13264 4829
rect 12926 4798 13264 4826
rect 12926 4795 12938 4798
rect 12880 4789 12938 4795
rect 13252 4795 13264 4798
rect 13298 4826 13310 4829
rect 13528 4829 13586 4835
rect 13528 4826 13540 4829
rect 13298 4798 13540 4826
rect 13298 4795 13310 4798
rect 13252 4789 13310 4795
rect 13528 4795 13540 4798
rect 13574 4795 13586 4829
rect 13528 4789 13586 4795
rect 14514 4823 14572 4829
rect 14514 4789 14526 4823
rect 14560 4820 14572 4823
rect 14600 4820 14628 4996
rect 16252 4978 17812 4998
rect 18169 4992 18640 5023
rect 19046 5050 19112 5098
rect 19046 4998 19056 5050
rect 19108 4998 19112 5050
rect 18169 4985 18277 4992
rect 14698 4891 14756 4897
rect 14698 4857 14710 4891
rect 14744 4888 14756 4891
rect 15438 4891 15496 4897
rect 15438 4888 15450 4891
rect 14744 4860 15450 4888
rect 14744 4857 14756 4860
rect 14698 4851 14756 4857
rect 15438 4857 15450 4860
rect 15484 4857 15496 4891
rect 15438 4851 15496 4857
rect 14882 4823 14940 4829
rect 14882 4820 14894 4823
rect 14560 4792 14894 4820
rect 14560 4789 14572 4792
rect 14514 4783 14572 4789
rect 14882 4789 14894 4792
rect 14928 4820 14940 4823
rect 15254 4823 15312 4829
rect 15254 4820 15266 4823
rect 14928 4792 15266 4820
rect 14928 4789 14940 4792
rect 14882 4783 14940 4789
rect 15254 4789 15266 4792
rect 15300 4820 15312 4823
rect 15530 4823 15588 4829
rect 15530 4820 15542 4823
rect 15300 4792 15542 4820
rect 15300 4789 15312 4792
rect 15254 4783 15312 4789
rect 15530 4789 15542 4792
rect 15576 4789 15588 4823
rect 15530 4783 15588 4789
rect 16536 4805 16594 4811
rect 11166 4765 11224 4771
rect 16536 4771 16548 4805
rect 16582 4802 16594 4805
rect 16622 4802 16650 4978
rect 16720 4873 16778 4879
rect 16720 4839 16732 4873
rect 16766 4870 16778 4873
rect 17460 4873 17518 4879
rect 17460 4870 17472 4873
rect 16766 4842 17472 4870
rect 16766 4839 16778 4842
rect 16720 4833 16778 4839
rect 17460 4839 17472 4842
rect 17506 4839 17518 4873
rect 17460 4833 17518 4839
rect 16904 4805 16962 4811
rect 16904 4802 16916 4805
rect 16582 4774 16916 4802
rect 16582 4771 16594 4774
rect 12604 4761 12662 4767
rect 11440 4732 11500 4756
rect 11440 4696 11454 4732
rect 11494 4730 11500 4732
rect 11494 4712 11818 4730
rect 12604 4727 12616 4761
rect 12650 4758 12662 4761
rect 13064 4761 13122 4767
rect 13064 4758 13076 4761
rect 12650 4730 13076 4758
rect 12650 4727 12662 4730
rect 12604 4721 12662 4727
rect 13064 4727 13076 4730
rect 13110 4758 13122 4761
rect 13436 4761 13494 4767
rect 16536 4765 16594 4771
rect 16904 4771 16916 4774
rect 16950 4802 16962 4805
rect 17276 4805 17334 4811
rect 17276 4802 17288 4805
rect 16950 4774 17288 4802
rect 16950 4771 16962 4774
rect 16904 4765 16962 4771
rect 17276 4771 17288 4774
rect 17322 4802 17334 4805
rect 17552 4805 17610 4811
rect 17552 4802 17564 4805
rect 17322 4774 17564 4802
rect 17322 4771 17334 4774
rect 17276 4765 17334 4771
rect 17552 4771 17564 4774
rect 17598 4771 17610 4805
rect 17552 4765 17610 4771
rect 13436 4758 13448 4761
rect 13110 4730 13448 4758
rect 13110 4727 13122 4730
rect 13064 4721 13122 4727
rect 11494 4696 12102 4712
rect 11440 4692 12102 4696
rect 11440 4680 11500 4692
rect 11774 4690 12102 4692
rect 12700 4694 12760 4700
rect 12700 4690 12714 4694
rect 11774 4660 12714 4690
rect 12748 4660 12760 4694
rect 11774 4652 12760 4660
rect 12700 4638 12760 4652
rect 10046 4590 11610 4598
rect 10046 4580 11612 4590
rect 10046 4567 10788 4580
rect 10844 4567 11612 4580
rect 10046 4533 10075 4567
rect 10109 4533 10167 4567
rect 10201 4533 10259 4567
rect 10293 4533 10351 4567
rect 10385 4566 10443 4567
rect 10477 4566 10535 4567
rect 10385 4533 10440 4566
rect 10492 4533 10535 4566
rect 10569 4533 10627 4567
rect 10661 4533 10719 4567
rect 10753 4533 10788 4567
rect 10845 4533 10903 4567
rect 10937 4533 10995 4567
rect 11029 4533 11087 4567
rect 11121 4533 11179 4567
rect 11213 4533 11271 4567
rect 11305 4533 11363 4567
rect 11397 4533 11455 4567
rect 11489 4533 11547 4567
rect 11581 4533 11612 4567
rect 13158 4554 13186 4730
rect 13436 4727 13448 4730
rect 13482 4727 13494 4761
rect 13436 4721 13494 4727
rect 14606 4755 14664 4761
rect 14606 4721 14618 4755
rect 14652 4752 14664 4755
rect 15066 4755 15124 4761
rect 15066 4752 15078 4755
rect 14652 4724 15078 4752
rect 14652 4721 14664 4724
rect 14606 4715 14664 4721
rect 15066 4721 15078 4724
rect 15112 4752 15124 4755
rect 15438 4755 15496 4761
rect 15438 4752 15450 4755
rect 15112 4724 15450 4752
rect 15112 4721 15124 4724
rect 15066 4715 15124 4721
rect 13718 4688 13770 4706
rect 14702 4688 14762 4694
rect 13716 4652 13730 4688
rect 13764 4684 14105 4688
rect 14702 4684 14716 4688
rect 13764 4654 14716 4684
rect 14750 4654 14762 4688
rect 13764 4652 14762 4654
rect 13716 4650 14762 4652
rect 13718 4640 13770 4650
rect 14082 4646 14762 4650
rect 14702 4632 14762 4646
rect 10046 4512 10440 4533
rect 10492 4522 10788 4533
rect 10844 4524 11612 4533
rect 12228 4534 13788 4554
rect 15160 4548 15188 4724
rect 15438 4721 15450 4724
rect 15484 4721 15496 4755
rect 15438 4715 15496 4721
rect 16628 4737 16686 4743
rect 16628 4703 16640 4737
rect 16674 4734 16686 4737
rect 17088 4737 17146 4743
rect 17088 4734 17100 4737
rect 16674 4706 17100 4734
rect 16674 4703 16686 4706
rect 15720 4682 15772 4700
rect 16628 4697 16686 4703
rect 17088 4703 17100 4706
rect 17134 4734 17146 4737
rect 17460 4737 17518 4743
rect 17460 4734 17472 4737
rect 17134 4706 17472 4734
rect 17134 4703 17146 4706
rect 17088 4697 17146 4703
rect 15718 4646 15732 4682
rect 15766 4666 15870 4682
rect 16724 4670 16784 4676
rect 16724 4666 16738 4670
rect 15766 4646 16738 4666
rect 15718 4644 16738 4646
rect 15720 4634 15772 4644
rect 15845 4636 16738 4644
rect 16772 4636 16784 4670
rect 15845 4628 16784 4636
rect 16724 4614 16784 4628
rect 10844 4522 11610 4524
rect 10492 4512 11610 4522
rect 10046 4502 11610 4512
rect 12228 4523 13036 4534
rect 13092 4523 13788 4534
rect 12228 4489 12257 4523
rect 12291 4489 12345 4523
rect 12379 4489 12437 4523
rect 12471 4489 12529 4523
rect 12563 4489 12621 4523
rect 12655 4489 12713 4523
rect 12747 4489 12805 4523
rect 12839 4489 12897 4523
rect 12931 4489 12989 4523
rect 13023 4489 13036 4523
rect 13115 4489 13173 4523
rect 13207 4489 13265 4523
rect 13299 4489 13357 4523
rect 13391 4489 13449 4523
rect 13483 4489 13541 4523
rect 13575 4489 13633 4523
rect 13667 4489 13725 4523
rect 13759 4489 13788 4523
rect 12228 4476 13036 4489
rect 13092 4476 13788 4489
rect 12228 4458 13788 4476
rect 14228 4528 15790 4548
rect 17182 4530 17210 4706
rect 17460 4703 17472 4706
rect 17506 4703 17518 4737
rect 17460 4697 17518 4703
rect 17742 4664 17794 4682
rect 18169 4664 18207 4985
rect 19046 4944 19112 4998
rect 18302 4894 19222 4900
rect 18302 4880 19226 4894
rect 18302 4869 18720 4880
rect 18778 4869 19226 4880
rect 18302 4835 18331 4869
rect 18365 4835 18423 4869
rect 18457 4835 18515 4869
rect 18549 4835 18607 4869
rect 18641 4835 18699 4869
rect 18778 4835 18791 4869
rect 18825 4835 18883 4869
rect 18917 4835 18975 4869
rect 19009 4835 19067 4869
rect 19101 4835 19159 4869
rect 19193 4835 19226 4869
rect 18302 4816 18720 4835
rect 18778 4828 19226 4835
rect 18778 4816 19222 4828
rect 18302 4804 19222 4816
rect 17740 4628 17754 4664
rect 17788 4628 18207 4664
rect 17740 4626 18207 4628
rect 17742 4616 17794 4626
rect 14228 4517 15038 4528
rect 15094 4517 15790 4528
rect 14228 4483 14257 4517
rect 14291 4483 14347 4517
rect 14381 4483 14439 4517
rect 14473 4483 14531 4517
rect 14565 4483 14623 4517
rect 14657 4483 14715 4517
rect 14749 4483 14807 4517
rect 14841 4483 14899 4517
rect 14933 4483 14991 4517
rect 15025 4483 15038 4517
rect 15117 4483 15175 4517
rect 15209 4483 15267 4517
rect 15301 4483 15359 4517
rect 15393 4483 15451 4517
rect 15485 4483 15543 4517
rect 15577 4483 15635 4517
rect 15669 4483 15727 4517
rect 15761 4483 15790 4517
rect 14228 4470 15038 4483
rect 15094 4470 15790 4483
rect 14228 4452 15790 4470
rect 16252 4510 17812 4530
rect 16252 4499 17060 4510
rect 17116 4499 17812 4510
rect 16252 4465 16281 4499
rect 16315 4465 16369 4499
rect 16403 4465 16461 4499
rect 16495 4465 16553 4499
rect 16587 4465 16645 4499
rect 16679 4465 16737 4499
rect 16771 4465 16829 4499
rect 16863 4465 16921 4499
rect 16955 4465 17013 4499
rect 17047 4465 17060 4499
rect 17139 4465 17197 4499
rect 17231 4465 17289 4499
rect 17323 4465 17381 4499
rect 17415 4465 17473 4499
rect 17507 4465 17565 4499
rect 17599 4465 17657 4499
rect 17691 4465 17749 4499
rect 17783 4465 17812 4499
rect 16252 4452 17060 4465
rect 17116 4452 17812 4465
rect 16252 4434 17812 4452
rect 5994 3382 6358 3388
rect 5994 3357 6194 3382
rect 6254 3357 6358 3382
rect 5994 3323 6023 3357
rect 6057 3323 6111 3357
rect 6145 3323 6194 3357
rect 6254 3323 6295 3357
rect 6329 3323 6358 3357
rect 5994 3320 6194 3323
rect 6254 3320 6358 3323
rect 5994 3292 6358 3320
rect 6104 3130 6198 3138
rect 6104 3078 6138 3130
rect 6190 3078 6198 3130
rect 6232 3136 6298 3138
rect 6232 3084 6238 3136
rect 6290 3084 6298 3136
rect 6232 3078 6298 3084
rect 6104 3072 6198 3078
rect 5994 2828 6358 2844
rect 5994 2813 6176 2828
rect 6236 2813 6358 2828
rect 5994 2779 6023 2813
rect 6057 2779 6111 2813
rect 6145 2779 6176 2813
rect 6237 2779 6295 2813
rect 6329 2779 6358 2813
rect 5994 2766 6176 2779
rect 6236 2766 6358 2779
rect 5994 2748 6358 2766
rect 7733 2338 7899 2340
rect 9700 2338 9883 2340
rect 11684 2338 11827 2340
rect 13613 2338 13829 2340
rect 15706 2338 15935 2340
rect 1716 2332 3278 2336
rect 3788 2332 3961 2334
rect 5747 2332 5875 2334
rect 1695 2318 3278 2332
rect 1695 2305 2604 2318
rect 2660 2305 3278 2318
rect 1695 2301 1745 2305
rect 1716 2271 1745 2301
rect 1779 2271 1835 2305
rect 1869 2271 1927 2305
rect 1961 2271 2019 2305
rect 2053 2271 2111 2305
rect 2145 2271 2203 2305
rect 2237 2271 2295 2305
rect 2329 2271 2387 2305
rect 2421 2271 2479 2305
rect 2513 2271 2571 2305
rect 2660 2271 2663 2305
rect 2697 2271 2755 2305
rect 2789 2271 2847 2305
rect 2881 2271 2939 2305
rect 2973 2271 3031 2305
rect 3065 2271 3123 2305
rect 3157 2271 3215 2305
rect 3249 2271 3278 2305
rect 1716 2260 2604 2271
rect 2660 2260 3278 2271
rect 1716 2240 3278 2260
rect 3786 2314 5348 2332
rect 3786 2301 4592 2314
rect 4648 2301 5348 2314
rect 3786 2267 3815 2301
rect 3849 2267 3905 2301
rect 3939 2267 3997 2301
rect 4031 2267 4089 2301
rect 4123 2267 4181 2301
rect 4215 2267 4273 2301
rect 4307 2267 4365 2301
rect 4399 2267 4457 2301
rect 4491 2267 4549 2301
rect 4583 2267 4592 2301
rect 4675 2267 4733 2301
rect 4767 2267 4825 2301
rect 4859 2267 4917 2301
rect 4951 2267 5009 2301
rect 5043 2267 5101 2301
rect 5135 2267 5193 2301
rect 5227 2267 5285 2301
rect 5319 2267 5348 2301
rect 3786 2256 4592 2267
rect 4648 2256 5348 2267
rect 2002 2067 2060 2073
rect 2002 2033 2014 2067
rect 2048 2064 2060 2067
rect 2088 2064 2116 2240
rect 3786 2236 5348 2256
rect 5742 2314 7300 2332
rect 5742 2301 6544 2314
rect 6600 2301 7300 2314
rect 7733 2320 9302 2338
rect 7733 2309 8546 2320
rect 5742 2267 5771 2301
rect 5805 2267 5857 2301
rect 5891 2267 5949 2301
rect 5983 2267 6041 2301
rect 6075 2267 6133 2301
rect 6167 2267 6225 2301
rect 6259 2267 6317 2301
rect 6351 2267 6409 2301
rect 6443 2267 6501 2301
rect 6535 2267 6544 2301
rect 6627 2267 6685 2301
rect 6719 2267 6777 2301
rect 6811 2267 6869 2301
rect 6903 2267 6961 2301
rect 6995 2267 7053 2301
rect 7087 2267 7145 2301
rect 7179 2267 7237 2301
rect 7271 2267 7300 2301
rect 5742 2256 6544 2267
rect 6600 2256 7300 2267
rect 5742 2236 7300 2256
rect 7740 2307 8546 2309
rect 8602 2307 9302 2320
rect 7740 2273 7769 2307
rect 7803 2273 7859 2307
rect 7893 2273 7951 2307
rect 7985 2273 8043 2307
rect 8077 2273 8135 2307
rect 8169 2273 8227 2307
rect 8261 2273 8319 2307
rect 8353 2273 8411 2307
rect 8445 2273 8503 2307
rect 8537 2273 8546 2307
rect 8629 2273 8687 2307
rect 8721 2273 8779 2307
rect 8813 2273 8871 2307
rect 8905 2273 8963 2307
rect 8997 2273 9055 2307
rect 9089 2273 9147 2307
rect 9181 2273 9239 2307
rect 9273 2273 9302 2307
rect 7740 2262 8546 2273
rect 8602 2262 9302 2273
rect 7740 2242 9302 2262
rect 9696 2320 11254 2338
rect 9696 2307 10498 2320
rect 10554 2307 11254 2320
rect 9696 2273 9725 2307
rect 9759 2273 9811 2307
rect 9845 2273 9903 2307
rect 9937 2273 9995 2307
rect 10029 2273 10087 2307
rect 10121 2273 10179 2307
rect 10213 2273 10271 2307
rect 10305 2273 10363 2307
rect 10397 2273 10455 2307
rect 10489 2273 10498 2307
rect 10581 2273 10639 2307
rect 10673 2273 10731 2307
rect 10765 2273 10823 2307
rect 10857 2273 10915 2307
rect 10949 2273 11007 2307
rect 11041 2273 11099 2307
rect 11133 2273 11191 2307
rect 11225 2273 11254 2307
rect 9696 2262 10498 2273
rect 10554 2262 11254 2273
rect 9696 2242 11254 2262
rect 11684 2320 13246 2338
rect 11684 2307 12490 2320
rect 12546 2307 13246 2320
rect 13613 2320 15198 2338
rect 13613 2309 14442 2320
rect 11684 2273 11713 2307
rect 11747 2273 11803 2307
rect 11837 2273 11895 2307
rect 11929 2273 11987 2307
rect 12021 2273 12079 2307
rect 12113 2273 12171 2307
rect 12205 2273 12263 2307
rect 12297 2273 12355 2307
rect 12389 2273 12447 2307
rect 12481 2273 12490 2307
rect 12573 2273 12631 2307
rect 12665 2273 12723 2307
rect 12757 2273 12815 2307
rect 12849 2273 12907 2307
rect 12941 2273 12999 2307
rect 13033 2273 13091 2307
rect 13125 2273 13183 2307
rect 13217 2273 13246 2307
rect 11684 2262 12490 2273
rect 12546 2262 13246 2273
rect 11684 2242 13246 2262
rect 13638 2307 14442 2309
rect 14498 2307 15198 2320
rect 13638 2273 13667 2307
rect 13701 2273 13755 2307
rect 13789 2273 13847 2307
rect 13881 2273 13939 2307
rect 13973 2273 14031 2307
rect 14065 2273 14123 2307
rect 14157 2273 14215 2307
rect 14249 2273 14307 2307
rect 14341 2273 14399 2307
rect 14433 2273 14442 2307
rect 14525 2273 14583 2307
rect 14617 2273 14675 2307
rect 14709 2273 14767 2307
rect 14801 2273 14859 2307
rect 14893 2273 14951 2307
rect 14985 2273 15043 2307
rect 15077 2273 15135 2307
rect 15169 2273 15198 2307
rect 13638 2262 14442 2273
rect 14498 2262 15198 2273
rect 13638 2242 15198 2262
rect 15700 2320 17262 2338
rect 15700 2307 16506 2320
rect 16562 2307 17262 2320
rect 15700 2273 15729 2307
rect 15763 2273 15819 2307
rect 15853 2273 15911 2307
rect 15945 2273 16003 2307
rect 16037 2273 16095 2307
rect 16129 2273 16187 2307
rect 16221 2273 16279 2307
rect 16313 2273 16371 2307
rect 16405 2273 16463 2307
rect 16497 2273 16506 2307
rect 16589 2273 16647 2307
rect 16681 2273 16739 2307
rect 16773 2273 16831 2307
rect 16865 2273 16923 2307
rect 16957 2273 17015 2307
rect 17049 2273 17107 2307
rect 17141 2273 17199 2307
rect 17233 2273 17262 2307
rect 15700 2262 16506 2273
rect 16562 2262 17262 2273
rect 15700 2242 17262 2262
rect 2186 2135 2244 2141
rect 2186 2101 2198 2135
rect 2232 2132 2244 2135
rect 2926 2135 2984 2141
rect 2926 2132 2938 2135
rect 2232 2104 2938 2132
rect 2232 2101 2244 2104
rect 2186 2095 2244 2101
rect 2926 2101 2938 2104
rect 2972 2101 2984 2135
rect 2926 2095 2984 2101
rect 2370 2067 2428 2073
rect 2370 2064 2382 2067
rect 2048 2036 2382 2064
rect 2048 2033 2060 2036
rect 2002 2027 2060 2033
rect 2370 2033 2382 2036
rect 2416 2064 2428 2067
rect 2742 2067 2800 2073
rect 2742 2064 2754 2067
rect 2416 2036 2754 2064
rect 2416 2033 2428 2036
rect 2370 2027 2428 2033
rect 2742 2033 2754 2036
rect 2788 2064 2800 2067
rect 3018 2067 3076 2073
rect 3018 2064 3030 2067
rect 2788 2036 3030 2064
rect 2788 2033 2800 2036
rect 2742 2027 2800 2033
rect 3018 2033 3030 2036
rect 3064 2033 3076 2067
rect 3018 2027 3076 2033
rect 4072 2063 4130 2069
rect 4072 2029 4084 2063
rect 4118 2060 4130 2063
rect 4158 2060 4186 2236
rect 4256 2131 4314 2137
rect 4256 2097 4268 2131
rect 4302 2128 4314 2131
rect 4996 2131 5054 2137
rect 4996 2128 5008 2131
rect 4302 2100 5008 2128
rect 4302 2097 4314 2100
rect 4256 2091 4314 2097
rect 4996 2097 5008 2100
rect 5042 2097 5054 2131
rect 4996 2091 5054 2097
rect 4440 2063 4498 2069
rect 4440 2060 4452 2063
rect 4118 2032 4452 2060
rect 4118 2029 4130 2032
rect 4072 2023 4130 2029
rect 4440 2029 4452 2032
rect 4486 2060 4498 2063
rect 4812 2063 4870 2069
rect 4812 2060 4824 2063
rect 4486 2032 4824 2060
rect 4486 2029 4498 2032
rect 4440 2023 4498 2029
rect 4812 2029 4824 2032
rect 4858 2060 4870 2063
rect 5088 2063 5146 2069
rect 5088 2060 5100 2063
rect 4858 2032 5100 2060
rect 4858 2029 4870 2032
rect 4812 2023 4870 2029
rect 5088 2029 5100 2032
rect 5134 2029 5146 2063
rect 5088 2023 5146 2029
rect 6024 2063 6082 2069
rect 6024 2029 6036 2063
rect 6070 2060 6082 2063
rect 6110 2060 6138 2236
rect 6208 2131 6266 2137
rect 6208 2097 6220 2131
rect 6254 2128 6266 2131
rect 6948 2131 7006 2137
rect 6948 2128 6960 2131
rect 6254 2100 6960 2128
rect 6254 2097 6266 2100
rect 6208 2091 6266 2097
rect 6948 2097 6960 2100
rect 6994 2097 7006 2131
rect 6948 2091 7006 2097
rect 8026 2069 8084 2075
rect 6392 2063 6450 2069
rect 6392 2060 6404 2063
rect 6070 2032 6404 2060
rect 6070 2029 6082 2032
rect 6024 2023 6082 2029
rect 6392 2029 6404 2032
rect 6438 2060 6450 2063
rect 6764 2063 6822 2069
rect 6764 2060 6776 2063
rect 6438 2032 6776 2060
rect 6438 2029 6450 2032
rect 6392 2023 6450 2029
rect 6764 2029 6776 2032
rect 6810 2060 6822 2063
rect 7040 2063 7098 2069
rect 7040 2060 7052 2063
rect 6810 2032 7052 2060
rect 6810 2029 6822 2032
rect 6764 2023 6822 2029
rect 7040 2029 7052 2032
rect 7086 2029 7098 2063
rect 8026 2035 8038 2069
rect 8072 2066 8084 2069
rect 8112 2066 8140 2242
rect 8210 2137 8268 2143
rect 8210 2103 8222 2137
rect 8256 2134 8268 2137
rect 8950 2137 9008 2143
rect 8950 2134 8962 2137
rect 8256 2106 8962 2134
rect 8256 2103 8268 2106
rect 8210 2097 8268 2103
rect 8950 2103 8962 2106
rect 8996 2103 9008 2137
rect 8950 2097 9008 2103
rect 8394 2069 8452 2075
rect 8394 2066 8406 2069
rect 8072 2038 8406 2066
rect 8072 2035 8084 2038
rect 8026 2029 8084 2035
rect 8394 2035 8406 2038
rect 8440 2066 8452 2069
rect 8766 2069 8824 2075
rect 8766 2066 8778 2069
rect 8440 2038 8778 2066
rect 8440 2035 8452 2038
rect 8394 2029 8452 2035
rect 8766 2035 8778 2038
rect 8812 2066 8824 2069
rect 9042 2069 9100 2075
rect 9042 2066 9054 2069
rect 8812 2038 9054 2066
rect 8812 2035 8824 2038
rect 8766 2029 8824 2035
rect 9042 2035 9054 2038
rect 9088 2035 9100 2069
rect 9042 2029 9100 2035
rect 9978 2069 10036 2075
rect 9978 2035 9990 2069
rect 10024 2066 10036 2069
rect 10064 2066 10092 2242
rect 10162 2137 10220 2143
rect 10162 2103 10174 2137
rect 10208 2134 10220 2137
rect 10902 2137 10960 2143
rect 10902 2134 10914 2137
rect 10208 2106 10914 2134
rect 10208 2103 10220 2106
rect 10162 2097 10220 2103
rect 10902 2103 10914 2106
rect 10948 2103 10960 2137
rect 10902 2097 10960 2103
rect 10346 2069 10404 2075
rect 10346 2066 10358 2069
rect 10024 2038 10358 2066
rect 10024 2035 10036 2038
rect 9978 2029 10036 2035
rect 10346 2035 10358 2038
rect 10392 2066 10404 2069
rect 10718 2069 10776 2075
rect 10718 2066 10730 2069
rect 10392 2038 10730 2066
rect 10392 2035 10404 2038
rect 10346 2029 10404 2035
rect 10718 2035 10730 2038
rect 10764 2066 10776 2069
rect 10994 2069 11052 2075
rect 10994 2066 11006 2069
rect 10764 2038 11006 2066
rect 10764 2035 10776 2038
rect 10718 2029 10776 2035
rect 10994 2035 11006 2038
rect 11040 2035 11052 2069
rect 10994 2029 11052 2035
rect 11970 2069 12028 2075
rect 11970 2035 11982 2069
rect 12016 2066 12028 2069
rect 12056 2066 12084 2242
rect 12154 2137 12212 2143
rect 12154 2103 12166 2137
rect 12200 2134 12212 2137
rect 12894 2137 12952 2143
rect 12894 2134 12906 2137
rect 12200 2106 12906 2134
rect 12200 2103 12212 2106
rect 12154 2097 12212 2103
rect 12894 2103 12906 2106
rect 12940 2103 12952 2137
rect 12894 2097 12952 2103
rect 12338 2069 12396 2075
rect 12338 2066 12350 2069
rect 12016 2038 12350 2066
rect 12016 2035 12028 2038
rect 11970 2029 12028 2035
rect 12338 2035 12350 2038
rect 12384 2066 12396 2069
rect 12710 2069 12768 2075
rect 12710 2066 12722 2069
rect 12384 2038 12722 2066
rect 12384 2035 12396 2038
rect 12338 2029 12396 2035
rect 12710 2035 12722 2038
rect 12756 2066 12768 2069
rect 12986 2069 13044 2075
rect 12986 2066 12998 2069
rect 12756 2038 12998 2066
rect 12756 2035 12768 2038
rect 12710 2029 12768 2035
rect 12986 2035 12998 2038
rect 13032 2035 13044 2069
rect 12986 2029 13044 2035
rect 13922 2069 13980 2075
rect 13922 2035 13934 2069
rect 13968 2066 13980 2069
rect 14008 2066 14036 2242
rect 14106 2137 14164 2143
rect 14106 2103 14118 2137
rect 14152 2134 14164 2137
rect 14846 2137 14904 2143
rect 14846 2134 14858 2137
rect 14152 2106 14858 2134
rect 14152 2103 14164 2106
rect 14106 2097 14164 2103
rect 14846 2103 14858 2106
rect 14892 2103 14904 2137
rect 14846 2097 14904 2103
rect 14290 2069 14348 2075
rect 14290 2066 14302 2069
rect 13968 2038 14302 2066
rect 13968 2035 13980 2038
rect 13922 2029 13980 2035
rect 14290 2035 14302 2038
rect 14336 2066 14348 2069
rect 14662 2069 14720 2075
rect 14662 2066 14674 2069
rect 14336 2038 14674 2066
rect 14336 2035 14348 2038
rect 14290 2029 14348 2035
rect 14662 2035 14674 2038
rect 14708 2066 14720 2069
rect 14938 2069 14996 2075
rect 14938 2066 14950 2069
rect 14708 2038 14950 2066
rect 14708 2035 14720 2038
rect 14662 2029 14720 2035
rect 14938 2035 14950 2038
rect 14984 2035 14996 2069
rect 14938 2029 14996 2035
rect 15986 2069 16044 2075
rect 15986 2035 15998 2069
rect 16032 2066 16044 2069
rect 16072 2066 16100 2242
rect 16170 2137 16228 2143
rect 16170 2103 16182 2137
rect 16216 2134 16228 2137
rect 16910 2137 16968 2143
rect 16910 2134 16922 2137
rect 16216 2106 16922 2134
rect 16216 2103 16228 2106
rect 16170 2097 16228 2103
rect 16910 2103 16922 2106
rect 16956 2103 16968 2137
rect 16910 2097 16968 2103
rect 16354 2069 16412 2075
rect 16354 2066 16366 2069
rect 16032 2038 16366 2066
rect 16032 2035 16044 2038
rect 15986 2029 16044 2035
rect 16354 2035 16366 2038
rect 16400 2066 16412 2069
rect 16726 2069 16784 2075
rect 16726 2066 16738 2069
rect 16400 2038 16738 2066
rect 16400 2035 16412 2038
rect 16354 2029 16412 2035
rect 16726 2035 16738 2038
rect 16772 2066 16784 2069
rect 17002 2069 17060 2075
rect 17002 2066 17014 2069
rect 16772 2038 17014 2066
rect 16772 2035 16784 2038
rect 16726 2029 16784 2035
rect 17002 2035 17014 2038
rect 17048 2035 17060 2069
rect 17002 2029 17060 2035
rect 7040 2023 7098 2029
rect 2094 1999 2152 2005
rect 2094 1965 2106 1999
rect 2140 1996 2152 1999
rect 2554 1999 2612 2005
rect 2554 1996 2566 1999
rect 2140 1968 2566 1996
rect 2140 1965 2152 1968
rect 2094 1959 2152 1965
rect 2554 1965 2566 1968
rect 2600 1996 2612 1999
rect 2926 1999 2984 2005
rect 8118 2001 8176 2007
rect 2926 1996 2938 1999
rect 2600 1968 2938 1996
rect 2600 1965 2612 1968
rect 2554 1959 2612 1965
rect 2192 1938 2258 1940
rect 2192 1886 2198 1938
rect 2250 1886 2258 1938
rect 2192 1882 2258 1886
rect 2648 1792 2676 1968
rect 2926 1965 2938 1968
rect 2972 1965 2984 1999
rect 2926 1959 2984 1965
rect 4164 1995 4222 2001
rect 4164 1961 4176 1995
rect 4210 1992 4222 1995
rect 4624 1995 4682 2001
rect 4624 1992 4636 1995
rect 4210 1964 4636 1992
rect 4210 1961 4222 1964
rect 4164 1955 4222 1961
rect 4624 1961 4636 1964
rect 4670 1992 4682 1995
rect 4996 1995 5054 2001
rect 4996 1992 5008 1995
rect 4670 1964 5008 1992
rect 4670 1961 4682 1964
rect 4624 1955 4682 1961
rect 3200 1926 3260 1950
rect 3200 1890 3214 1926
rect 3254 1924 3260 1926
rect 4260 1928 4320 1934
rect 4260 1924 4274 1928
rect 3254 1894 4274 1924
rect 4308 1894 4320 1928
rect 3254 1890 4320 1894
rect 3200 1886 4320 1890
rect 3200 1874 3260 1886
rect 4260 1872 4320 1886
rect 1716 1778 3278 1792
rect 4718 1788 4746 1964
rect 4996 1961 5008 1964
rect 5042 1961 5054 1995
rect 4996 1955 5054 1961
rect 6116 1995 6174 2001
rect 6116 1961 6128 1995
rect 6162 1992 6174 1995
rect 6576 1995 6634 2001
rect 6576 1992 6588 1995
rect 6162 1964 6588 1992
rect 6162 1961 6174 1964
rect 6116 1955 6174 1961
rect 6576 1961 6588 1964
rect 6622 1992 6634 1995
rect 6948 1995 7006 2001
rect 6948 1992 6960 1995
rect 6622 1964 6960 1992
rect 6622 1961 6634 1964
rect 6576 1955 6634 1961
rect 5278 1922 5330 1940
rect 6212 1928 6272 1934
rect 6212 1924 6226 1928
rect 5518 1922 6226 1924
rect 5276 1886 5290 1922
rect 5324 1894 6226 1922
rect 6260 1894 6272 1928
rect 5324 1886 6272 1894
rect 5276 1884 5565 1886
rect 5278 1874 5330 1884
rect 6212 1872 6272 1886
rect 6670 1788 6698 1964
rect 6948 1961 6960 1964
rect 6994 1961 7006 1995
rect 8118 1967 8130 2001
rect 8164 1998 8176 2001
rect 8578 2001 8636 2007
rect 8578 1998 8590 2001
rect 8164 1970 8590 1998
rect 8164 1967 8176 1970
rect 8118 1961 8176 1967
rect 8578 1967 8590 1970
rect 8624 1998 8636 2001
rect 8950 2001 9008 2007
rect 8950 1998 8962 2001
rect 8624 1970 8962 1998
rect 8624 1967 8636 1970
rect 8578 1961 8636 1967
rect 6948 1955 7006 1961
rect 7230 1922 7282 1940
rect 8214 1934 8274 1940
rect 8214 1930 8228 1934
rect 7456 1922 8228 1930
rect 7228 1886 7242 1922
rect 7276 1900 8228 1922
rect 8262 1900 8274 1934
rect 7276 1892 8274 1900
rect 7276 1886 7517 1892
rect 7228 1884 7517 1886
rect 7230 1874 7282 1884
rect 8214 1878 8274 1892
rect 8672 1794 8700 1970
rect 8950 1967 8962 1970
rect 8996 1967 9008 2001
rect 8950 1961 9008 1967
rect 10070 2001 10128 2007
rect 10070 1967 10082 2001
rect 10116 1998 10128 2001
rect 10530 2001 10588 2007
rect 10530 1998 10542 2001
rect 10116 1970 10542 1998
rect 10116 1967 10128 1970
rect 10070 1961 10128 1967
rect 10530 1967 10542 1970
rect 10576 1998 10588 2001
rect 10902 2001 10960 2007
rect 10902 1998 10914 2001
rect 10576 1970 10914 1998
rect 10576 1967 10588 1970
rect 10530 1961 10588 1967
rect 9232 1928 9284 1946
rect 10166 1934 10226 1940
rect 10166 1930 10180 1934
rect 9472 1928 10180 1930
rect 9230 1892 9244 1928
rect 9278 1900 10180 1928
rect 10214 1900 10226 1934
rect 9278 1892 10226 1900
rect 9230 1890 9519 1892
rect 9232 1880 9284 1890
rect 10166 1878 10226 1892
rect 10624 1794 10652 1970
rect 10902 1967 10914 1970
rect 10948 1967 10960 2001
rect 10902 1961 10960 1967
rect 12062 2001 12120 2007
rect 12062 1967 12074 2001
rect 12108 1998 12120 2001
rect 12522 2001 12580 2007
rect 12522 1998 12534 2001
rect 12108 1970 12534 1998
rect 12108 1967 12120 1970
rect 12062 1961 12120 1967
rect 12522 1967 12534 1970
rect 12568 1998 12580 2001
rect 12894 2001 12952 2007
rect 12894 1998 12906 2001
rect 12568 1970 12906 1998
rect 12568 1967 12580 1970
rect 12522 1961 12580 1967
rect 11184 1928 11236 1946
rect 12158 1934 12218 1940
rect 12158 1930 12172 1934
rect 11317 1928 12172 1930
rect 11182 1892 11196 1928
rect 11230 1900 12172 1928
rect 12206 1900 12218 1934
rect 11230 1892 12218 1900
rect 11182 1890 11382 1892
rect 11184 1880 11236 1890
rect 12158 1878 12218 1892
rect 12616 1794 12644 1970
rect 12894 1967 12906 1970
rect 12940 1967 12952 2001
rect 12894 1961 12952 1967
rect 14014 2001 14072 2007
rect 14014 1967 14026 2001
rect 14060 1998 14072 2001
rect 14474 2001 14532 2007
rect 14474 1998 14486 2001
rect 14060 1970 14486 1998
rect 14060 1967 14072 1970
rect 14014 1961 14072 1967
rect 14474 1967 14486 1970
rect 14520 1998 14532 2001
rect 14846 2001 14904 2007
rect 14846 1998 14858 2001
rect 14520 1970 14858 1998
rect 14520 1967 14532 1970
rect 14474 1961 14532 1967
rect 13176 1928 13228 1946
rect 14110 1934 14170 1940
rect 14110 1930 14124 1934
rect 13416 1928 14124 1930
rect 13174 1892 13188 1928
rect 13222 1900 14124 1928
rect 14158 1900 14170 1934
rect 13222 1892 14170 1900
rect 13174 1890 13463 1892
rect 13176 1880 13228 1890
rect 14110 1878 14170 1892
rect 14568 1794 14596 1970
rect 14846 1967 14858 1970
rect 14892 1967 14904 2001
rect 14846 1961 14904 1967
rect 16078 2001 16136 2007
rect 16078 1967 16090 2001
rect 16124 1998 16136 2001
rect 16538 2001 16596 2007
rect 16538 1998 16550 2001
rect 16124 1970 16550 1998
rect 16124 1967 16136 1970
rect 16078 1961 16136 1967
rect 16538 1967 16550 1970
rect 16584 1998 16596 2001
rect 16910 2001 16968 2007
rect 16910 1998 16922 2001
rect 16584 1970 16922 1998
rect 16584 1967 16596 1970
rect 16538 1961 16596 1967
rect 15128 1928 15180 1946
rect 16174 1934 16234 1940
rect 16174 1930 16188 1934
rect 15538 1928 16188 1930
rect 15126 1892 15140 1928
rect 15174 1900 16188 1928
rect 16222 1900 16234 1934
rect 15174 1892 16234 1900
rect 15126 1890 15575 1892
rect 15128 1880 15180 1890
rect 16174 1878 16234 1892
rect 16632 1794 16660 1970
rect 16910 1967 16922 1970
rect 16956 1967 16968 2001
rect 16910 1961 16968 1967
rect 17192 1928 17244 1946
rect 17362 1930 17488 1982
rect 17362 1928 17402 1930
rect 17190 1892 17204 1928
rect 17238 1892 17402 1928
rect 17190 1890 17402 1892
rect 17192 1880 17244 1890
rect 17362 1876 17402 1890
rect 17454 1876 17488 1930
rect 17362 1828 17488 1876
rect 1716 1761 2604 1778
rect 2656 1761 3278 1778
rect 1716 1727 1745 1761
rect 1779 1727 1835 1761
rect 1869 1727 1927 1761
rect 1961 1727 2019 1761
rect 2053 1727 2111 1761
rect 2145 1727 2203 1761
rect 2237 1727 2295 1761
rect 2329 1727 2387 1761
rect 2421 1727 2479 1761
rect 2513 1727 2571 1761
rect 2656 1727 2663 1761
rect 2697 1727 2755 1761
rect 2789 1727 2847 1761
rect 2881 1727 2939 1761
rect 2973 1727 3031 1761
rect 3065 1727 3123 1761
rect 3157 1727 3215 1761
rect 3249 1727 3278 1761
rect 1716 1720 2604 1727
rect 2656 1720 3278 1727
rect 3786 1768 5348 1788
rect 3786 1757 4596 1768
rect 4652 1757 5348 1768
rect 3786 1725 3815 1757
rect 1716 1696 3278 1720
rect 3783 1723 3815 1725
rect 3849 1723 3905 1757
rect 3939 1723 3997 1757
rect 4031 1723 4089 1757
rect 4123 1723 4181 1757
rect 4215 1723 4273 1757
rect 4307 1723 4365 1757
rect 4399 1723 4457 1757
rect 4491 1723 4549 1757
rect 4583 1723 4596 1757
rect 4675 1723 4733 1757
rect 4767 1723 4825 1757
rect 4859 1723 4917 1757
rect 4951 1723 5009 1757
rect 5043 1723 5101 1757
rect 5135 1723 5193 1757
rect 5227 1723 5285 1757
rect 5319 1723 5348 1757
rect 5742 1768 7300 1788
rect 5742 1757 6548 1768
rect 6604 1757 7300 1768
rect 5742 1725 5771 1757
rect 3783 1710 4596 1723
rect 4652 1710 5348 1723
rect 1719 1692 1849 1696
rect 3783 1694 5348 1710
rect 5738 1723 5771 1725
rect 5805 1723 5857 1757
rect 5891 1723 5949 1757
rect 5983 1723 6041 1757
rect 6075 1723 6133 1757
rect 6167 1723 6225 1757
rect 6259 1723 6317 1757
rect 6351 1723 6409 1757
rect 6443 1723 6501 1757
rect 6535 1723 6548 1757
rect 6627 1723 6685 1757
rect 6719 1723 6777 1757
rect 6811 1723 6869 1757
rect 6903 1723 6961 1757
rect 6995 1723 7053 1757
rect 7087 1723 7145 1757
rect 7179 1723 7237 1757
rect 7271 1723 7300 1757
rect 5738 1710 6548 1723
rect 6604 1710 7300 1723
rect 5738 1694 7300 1710
rect 7740 1774 9302 1794
rect 7740 1763 8550 1774
rect 8606 1763 9302 1774
rect 7740 1729 7769 1763
rect 7803 1729 7859 1763
rect 7893 1729 7951 1763
rect 7985 1729 8043 1763
rect 8077 1729 8135 1763
rect 8169 1729 8227 1763
rect 8261 1729 8319 1763
rect 8353 1729 8411 1763
rect 8445 1729 8503 1763
rect 8537 1729 8550 1763
rect 8629 1729 8687 1763
rect 8721 1729 8779 1763
rect 8813 1729 8871 1763
rect 8905 1729 8963 1763
rect 8997 1729 9055 1763
rect 9089 1729 9147 1763
rect 9181 1729 9239 1763
rect 9273 1729 9302 1763
rect 7740 1716 8550 1729
rect 8606 1716 9302 1729
rect 7740 1698 9302 1716
rect 9696 1774 11254 1794
rect 9696 1763 10502 1774
rect 10558 1763 11254 1774
rect 9696 1729 9725 1763
rect 9759 1729 9811 1763
rect 9845 1729 9903 1763
rect 9937 1729 9995 1763
rect 10029 1729 10087 1763
rect 10121 1729 10179 1763
rect 10213 1729 10271 1763
rect 10305 1729 10363 1763
rect 10397 1729 10455 1763
rect 10489 1729 10502 1763
rect 10581 1729 10639 1763
rect 10673 1729 10731 1763
rect 10765 1729 10823 1763
rect 10857 1729 10915 1763
rect 10949 1729 11007 1763
rect 11041 1729 11099 1763
rect 11133 1729 11191 1763
rect 11225 1729 11254 1763
rect 9696 1716 10502 1729
rect 10558 1716 11254 1729
rect 9696 1698 11254 1716
rect 11684 1774 13246 1794
rect 11684 1763 12494 1774
rect 12550 1763 13246 1774
rect 11684 1729 11713 1763
rect 11747 1729 11803 1763
rect 11837 1729 11895 1763
rect 11929 1729 11987 1763
rect 12021 1729 12079 1763
rect 12113 1729 12171 1763
rect 12205 1729 12263 1763
rect 12297 1729 12355 1763
rect 12389 1729 12447 1763
rect 12481 1729 12494 1763
rect 12573 1729 12631 1763
rect 12665 1729 12723 1763
rect 12757 1729 12815 1763
rect 12849 1729 12907 1763
rect 12941 1729 12999 1763
rect 13033 1729 13091 1763
rect 13125 1729 13183 1763
rect 13217 1729 13246 1763
rect 11684 1716 12494 1729
rect 12550 1716 13246 1729
rect 11684 1698 13246 1716
rect 13638 1774 15198 1794
rect 13638 1763 14446 1774
rect 14502 1763 15198 1774
rect 13638 1729 13667 1763
rect 13701 1729 13755 1763
rect 13789 1729 13847 1763
rect 13881 1729 13939 1763
rect 13973 1729 14031 1763
rect 14065 1729 14123 1763
rect 14157 1729 14215 1763
rect 14249 1729 14307 1763
rect 14341 1729 14399 1763
rect 14433 1729 14446 1763
rect 14525 1729 14583 1763
rect 14617 1729 14675 1763
rect 14709 1729 14767 1763
rect 14801 1729 14859 1763
rect 14893 1729 14951 1763
rect 14985 1729 15043 1763
rect 15077 1729 15135 1763
rect 15169 1729 15198 1763
rect 15700 1774 17262 1794
rect 15700 1763 16510 1774
rect 16566 1763 17262 1774
rect 15700 1731 15729 1763
rect 13638 1716 14446 1729
rect 14502 1716 15198 1729
rect 13638 1698 15198 1716
rect 15681 1729 15729 1731
rect 15763 1729 15819 1763
rect 15853 1729 15911 1763
rect 15945 1729 16003 1763
rect 16037 1729 16095 1763
rect 16129 1729 16187 1763
rect 16221 1729 16279 1763
rect 16313 1729 16371 1763
rect 16405 1729 16463 1763
rect 16497 1729 16510 1763
rect 16589 1729 16647 1763
rect 16681 1729 16739 1763
rect 16773 1729 16831 1763
rect 16865 1729 16923 1763
rect 16957 1729 17015 1763
rect 17049 1729 17107 1763
rect 17141 1729 17199 1763
rect 17233 1729 17262 1763
rect 15681 1716 16510 1729
rect 16566 1716 17262 1729
rect 15681 1700 17262 1716
rect 15700 1698 17262 1700
rect 3786 1692 5348 1694
rect 5742 1692 7300 1694
<< via1 >>
rect 18768 43898 18962 44096
rect 18562 42805 18579 42820
rect 18579 42805 18613 42820
rect 18613 42805 18624 42820
rect 18562 42762 18624 42805
rect 19124 42747 19186 42782
rect 19124 42724 19157 42747
rect 19157 42724 19186 42747
rect 18540 40943 18602 40948
rect 18540 40909 18563 40943
rect 18563 40909 18597 40943
rect 18597 40909 18602 40943
rect 18540 40890 18602 40909
rect 19106 40909 19107 40940
rect 19107 40909 19141 40940
rect 19141 40909 19168 40940
rect 19106 40882 19168 40909
rect 18564 39297 18571 39320
rect 18571 39297 18605 39320
rect 18605 39297 18626 39320
rect 18564 39262 18626 39297
rect 19106 39297 19115 39316
rect 19115 39297 19149 39316
rect 19149 39297 19168 39316
rect 19106 39258 19168 39297
rect 18572 38069 18634 38124
rect 18572 38066 18585 38069
rect 18585 38066 18619 38069
rect 18619 38066 18634 38069
rect 19122 38127 19129 38140
rect 19129 38127 19163 38140
rect 19163 38127 19184 38140
rect 19122 38082 19184 38127
rect 18580 37011 18642 37054
rect 18580 36996 18597 37011
rect 18597 36996 18631 37011
rect 18631 36996 18642 37011
rect 19128 37011 19190 37044
rect 19128 36986 19141 37011
rect 19141 36986 19175 37011
rect 19175 36986 19190 37011
rect 18598 36215 18652 36256
rect 18598 36200 18605 36215
rect 18605 36200 18639 36215
rect 18639 36200 18652 36215
rect 19142 36273 19149 36284
rect 19149 36273 19183 36284
rect 19183 36273 19200 36284
rect 19142 36228 19200 36273
rect 18618 34091 18684 34132
rect 18618 34066 18629 34091
rect 18629 34066 18663 34091
rect 18663 34066 18684 34091
rect 19160 34091 19226 34142
rect 19160 34076 19173 34091
rect 19173 34076 19207 34091
rect 19207 34076 19226 34091
rect 18618 31809 18684 31850
rect 18618 31784 18629 31809
rect 18629 31784 18663 31809
rect 18663 31784 18684 31809
rect 19160 31809 19226 31860
rect 19160 31794 19173 31809
rect 19173 31794 19207 31809
rect 19207 31794 19226 31809
rect 18622 29563 18688 29604
rect 18622 29538 18633 29563
rect 18633 29538 18667 29563
rect 18667 29538 18688 29563
rect 19164 29563 19230 29614
rect 19164 29548 19177 29563
rect 19177 29548 19211 29563
rect 19211 29548 19230 29563
rect 18614 27377 18680 27418
rect 18614 27352 18625 27377
rect 18625 27352 18659 27377
rect 18659 27352 18680 27377
rect 19156 27377 19222 27428
rect 19156 27362 19169 27377
rect 19169 27362 19203 27377
rect 19203 27362 19222 27377
rect 18618 25131 18684 25172
rect 18618 25106 18629 25131
rect 18629 25106 18663 25131
rect 18663 25106 18684 25131
rect 19160 25131 19226 25182
rect 19160 25116 19173 25131
rect 19173 25116 19207 25131
rect 19207 25116 19226 25131
rect 8536 23389 8602 23400
rect 8536 23355 8561 23389
rect 8561 23355 8602 23389
rect 8536 23334 8602 23355
rect 10782 23393 10848 23404
rect 10782 23359 10807 23393
rect 10807 23359 10848 23393
rect 10782 23338 10848 23359
rect 12968 23385 13034 23396
rect 12968 23351 12993 23385
rect 12993 23351 13034 23385
rect 12968 23330 13034 23351
rect 15214 23389 15280 23400
rect 15214 23355 15239 23389
rect 15239 23355 15280 23389
rect 15214 23334 15280 23355
rect 17496 23389 17562 23400
rect 17496 23355 17521 23389
rect 17521 23355 17562 23389
rect 17496 23334 17562 23355
rect 8546 22845 8612 22858
rect 8546 22811 8561 22845
rect 8561 22811 8612 22845
rect 8546 22792 8612 22811
rect 10792 22849 10858 22862
rect 10792 22815 10807 22849
rect 10807 22815 10858 22849
rect 10792 22796 10858 22815
rect 12978 22841 13044 22854
rect 12978 22807 12993 22841
rect 12993 22807 13044 22841
rect 12978 22788 13044 22807
rect 15224 22845 15290 22858
rect 15224 22811 15239 22845
rect 15239 22811 15290 22845
rect 15224 22792 15290 22811
rect 17506 22845 17572 22858
rect 17506 22811 17521 22845
rect 17521 22811 17572 22845
rect 17506 22792 17572 22811
rect 9540 17811 9600 17822
rect 9540 17777 9551 17811
rect 9551 17777 9585 17811
rect 9585 17777 9600 17811
rect 9540 17762 9600 17777
rect 16455 17701 16523 17714
rect 15683 17663 15751 17674
rect 15683 17629 15688 17663
rect 15688 17629 15722 17663
rect 15722 17629 15751 17663
rect 16455 17667 16466 17701
rect 16466 17667 16500 17701
rect 16500 17667 16523 17701
rect 16455 17652 16523 17667
rect 17335 17703 17403 17714
rect 17335 17669 17340 17703
rect 17340 17669 17374 17703
rect 17374 17669 17403 17703
rect 17335 17652 17403 17669
rect 18121 17693 18189 17704
rect 18121 17659 18142 17693
rect 18142 17659 18189 17693
rect 18121 17642 18189 17659
rect 19219 17695 19287 17708
rect 19219 17661 19230 17695
rect 19230 17661 19264 17695
rect 19264 17661 19287 17695
rect 19219 17646 19287 17661
rect 15683 17612 15751 17629
rect 20099 17697 20167 17708
rect 20099 17663 20104 17697
rect 20104 17663 20138 17697
rect 20138 17663 20167 17697
rect 20099 17646 20167 17663
rect 20885 17687 20953 17698
rect 20885 17653 20906 17687
rect 20906 17653 20953 17687
rect 20885 17636 20953 17653
rect 21475 17685 21543 17698
rect 21475 17651 21486 17685
rect 21486 17651 21520 17685
rect 21520 17651 21543 17685
rect 21475 17636 21543 17651
rect 22355 17687 22423 17698
rect 22355 17653 22360 17687
rect 22360 17653 22394 17687
rect 22394 17653 22423 17687
rect 22355 17636 22423 17653
rect 23141 17677 23209 17688
rect 23141 17643 23162 17677
rect 23162 17643 23209 17677
rect 23141 17626 23209 17643
rect 6646 17504 6722 17576
rect 9536 17267 9594 17278
rect 9536 17233 9551 17267
rect 9551 17233 9585 17267
rect 9585 17233 9594 17267
rect 9536 17218 9594 17233
rect 11414 16986 11474 17042
rect 4590 16603 4642 16624
rect 4590 16570 4623 16603
rect 4623 16570 4642 16603
rect 6006 16340 6076 16406
rect 4976 16059 5034 16074
rect 4976 16025 4991 16059
rect 4991 16025 5034 16059
rect 4976 16020 5034 16025
rect 4746 15859 4808 15874
rect 4746 15825 4779 15859
rect 4779 15825 4808 15859
rect 4746 15814 4808 15825
rect 6712 15749 6780 15768
rect 6712 15715 6729 15749
rect 6729 15715 6763 15749
rect 6763 15715 6780 15749
rect 6712 15706 6780 15715
rect 4976 15490 5030 15502
rect 4976 15456 5006 15490
rect 5006 15456 5030 15490
rect 4976 15448 5030 15456
rect 4898 15315 4966 15332
rect 4898 15281 4905 15315
rect 4905 15281 4963 15315
rect 4963 15281 4966 15315
rect 4898 15270 4966 15281
rect 4582 15039 4648 15052
rect 4582 15005 4599 15039
rect 4599 15005 4633 15039
rect 4633 15005 4648 15039
rect 4582 14986 4648 15005
rect 6608 15400 6660 15408
rect 6608 15364 6632 15400
rect 6632 15364 6660 15400
rect 6608 15356 6660 15364
rect 6130 15249 6198 15264
rect 6130 15215 6147 15249
rect 6147 15215 6181 15249
rect 6181 15215 6198 15249
rect 6130 15202 6198 15215
rect 7114 15205 7182 15218
rect 7114 15171 7131 15205
rect 7131 15171 7182 15205
rect 7114 15156 7182 15171
rect 5012 14495 5078 14508
rect 5012 14461 5059 14495
rect 5059 14461 5078 14495
rect 5012 14442 5078 14461
rect 4682 14295 4754 14314
rect 4682 14261 4697 14295
rect 4697 14261 4731 14295
rect 4731 14261 4754 14295
rect 4682 14244 4754 14261
rect 5030 13838 5090 13900
rect 4884 13751 4956 13770
rect 4884 13717 4915 13751
rect 4915 13717 4956 13751
rect 4884 13700 4956 13717
rect 4576 13371 4648 13384
rect 4576 13337 4591 13371
rect 4591 13337 4625 13371
rect 4625 13337 4648 13371
rect 4576 13318 4648 13337
rect 5794 14705 5862 14716
rect 5794 14671 5813 14705
rect 5813 14671 5862 14705
rect 5794 14654 5862 14671
rect 6350 14283 6418 14294
rect 6350 14249 6405 14283
rect 6405 14249 6418 14283
rect 6350 14232 6418 14249
rect 7916 14267 7984 14284
rect 7916 14233 7935 14267
rect 7935 14233 7969 14267
rect 7969 14233 7984 14267
rect 7916 14222 7984 14233
rect 9456 16607 9508 16628
rect 9456 16574 9489 16607
rect 9489 16574 9508 16607
rect 10872 16344 10942 16410
rect 9842 16063 9900 16078
rect 9842 16029 9857 16063
rect 9857 16029 9900 16063
rect 9842 16024 9900 16029
rect 9612 15863 9674 15878
rect 9612 15829 9645 15863
rect 9645 15829 9674 15863
rect 9612 15818 9674 15829
rect 11578 15753 11646 15772
rect 11578 15719 11595 15753
rect 11595 15719 11629 15753
rect 11629 15719 11646 15753
rect 11578 15710 11646 15719
rect 9842 15494 9896 15506
rect 9842 15460 9872 15494
rect 9872 15460 9896 15494
rect 9842 15452 9896 15460
rect 9764 15319 9832 15336
rect 9764 15285 9771 15319
rect 9771 15285 9829 15319
rect 9829 15285 9832 15319
rect 9764 15274 9832 15285
rect 9448 15043 9514 15056
rect 9448 15009 9465 15043
rect 9465 15009 9499 15043
rect 9499 15009 9514 15043
rect 9448 14990 9514 15009
rect 11474 15404 11526 15412
rect 11474 15368 11498 15404
rect 11498 15368 11526 15404
rect 11474 15360 11526 15368
rect 10996 15253 11064 15268
rect 10996 15219 11013 15253
rect 11013 15219 11047 15253
rect 11047 15219 11064 15253
rect 10996 15206 11064 15219
rect 11980 15209 12048 15222
rect 11980 15175 11997 15209
rect 11997 15175 12048 15209
rect 11980 15160 12048 15175
rect 9878 14499 9944 14512
rect 9878 14465 9925 14499
rect 9925 14465 9944 14499
rect 9878 14446 9944 14465
rect 9548 14299 9620 14318
rect 9548 14265 9563 14299
rect 9563 14265 9597 14299
rect 9597 14265 9620 14299
rect 9548 14248 9620 14265
rect 5298 13304 5360 13356
rect 6012 13880 6064 13890
rect 6012 13846 6020 13880
rect 6020 13846 6054 13880
rect 6054 13846 6064 13880
rect 6012 13838 6064 13846
rect 6110 13920 6162 13930
rect 6110 13886 6118 13920
rect 6118 13886 6152 13920
rect 6152 13886 6162 13920
rect 6110 13878 6162 13886
rect 6208 13830 6260 13886
rect 6828 13909 6896 13918
rect 6828 13875 6857 13909
rect 6857 13875 6896 13909
rect 6828 13856 6896 13875
rect 7652 13882 7704 13936
rect 7866 13960 7946 13980
rect 7866 13918 7880 13960
rect 7880 13918 7930 13960
rect 7930 13918 7946 13960
rect 7866 13904 7946 13918
rect 9896 13842 9956 13904
rect 5862 13739 5930 13754
rect 5862 13705 5887 13739
rect 5887 13705 5930 13739
rect 9750 13755 9822 13774
rect 5862 13692 5930 13705
rect 7656 13676 7724 13738
rect 9750 13721 9781 13755
rect 9781 13721 9822 13755
rect 9750 13704 9822 13721
rect 5984 13441 6052 13450
rect 5984 13407 6011 13441
rect 6011 13407 6052 13441
rect 5984 13390 6052 13407
rect 6140 13334 6194 13338
rect 6140 13298 6146 13334
rect 6146 13298 6182 13334
rect 6182 13298 6194 13334
rect 6140 13286 6194 13298
rect 7136 13365 7204 13378
rect 7136 13331 7191 13365
rect 7191 13331 7204 13365
rect 7136 13316 7204 13331
rect 9442 13375 9514 13388
rect 9442 13341 9457 13375
rect 9457 13341 9491 13375
rect 9491 13341 9514 13375
rect 9442 13322 9514 13341
rect 10660 14709 10728 14720
rect 10660 14675 10679 14709
rect 10679 14675 10728 14709
rect 16453 17157 16521 17172
rect 15691 17119 15759 17134
rect 15691 17085 15722 17119
rect 15722 17085 15759 17119
rect 16453 17123 16466 17157
rect 16466 17123 16500 17157
rect 16500 17123 16521 17157
rect 16453 17110 16521 17123
rect 17343 17159 17411 17174
rect 17343 17125 17374 17159
rect 17374 17125 17411 17159
rect 17343 17112 17411 17125
rect 18101 17149 18169 17166
rect 18101 17115 18108 17149
rect 18108 17115 18142 17149
rect 18142 17115 18169 17149
rect 18101 17104 18169 17115
rect 15691 17072 15759 17085
rect 19217 17151 19285 17166
rect 19217 17117 19230 17151
rect 19230 17117 19264 17151
rect 19264 17117 19285 17151
rect 19217 17104 19285 17117
rect 20107 17153 20175 17168
rect 20107 17119 20138 17153
rect 20138 17119 20175 17153
rect 20107 17106 20175 17119
rect 20865 17143 20933 17160
rect 20865 17109 20872 17143
rect 20872 17109 20906 17143
rect 20906 17109 20933 17143
rect 20865 17098 20933 17109
rect 21473 17141 21541 17156
rect 21473 17107 21486 17141
rect 21486 17107 21520 17141
rect 21520 17107 21541 17141
rect 21473 17094 21541 17107
rect 22363 17143 22431 17158
rect 22363 17109 22394 17143
rect 22394 17109 22431 17143
rect 22363 17096 22431 17109
rect 23121 17133 23189 17150
rect 23121 17099 23128 17133
rect 23128 17099 23162 17133
rect 23162 17099 23189 17133
rect 23121 17088 23189 17099
rect 16430 16711 16498 16722
rect 16430 16677 16457 16711
rect 16457 16677 16491 16711
rect 16491 16677 16498 16711
rect 16430 16660 16498 16677
rect 17188 16701 17256 16714
rect 17188 16667 17225 16701
rect 17225 16667 17256 16701
rect 17188 16652 17256 16667
rect 18078 16703 18146 16716
rect 18078 16669 18099 16703
rect 18099 16669 18133 16703
rect 18133 16669 18146 16703
rect 18078 16654 18146 16669
rect 18686 16701 18754 16712
rect 18686 16667 18713 16701
rect 18713 16667 18747 16701
rect 18747 16667 18754 16701
rect 18686 16650 18754 16667
rect 19444 16691 19512 16704
rect 19444 16657 19481 16691
rect 19481 16657 19512 16691
rect 19444 16642 19512 16657
rect 20334 16693 20402 16706
rect 20334 16659 20355 16693
rect 20355 16659 20389 16693
rect 20389 16659 20402 16693
rect 20334 16644 20402 16659
rect 21450 16695 21518 16706
rect 21450 16661 21477 16695
rect 21477 16661 21511 16695
rect 21511 16661 21518 16695
rect 21450 16644 21518 16661
rect 22208 16685 22276 16698
rect 22208 16651 22245 16685
rect 22245 16651 22276 16685
rect 22208 16636 22276 16651
rect 23098 16687 23166 16700
rect 23098 16653 23119 16687
rect 23119 16653 23153 16687
rect 23153 16653 23166 16687
rect 23098 16638 23166 16653
rect 16410 16167 16478 16184
rect 16410 16133 16457 16167
rect 16457 16133 16478 16167
rect 16410 16122 16478 16133
rect 17196 16157 17264 16174
rect 17196 16123 17225 16157
rect 17225 16123 17259 16157
rect 17259 16123 17264 16157
rect 17196 16112 17264 16123
rect 18076 16159 18144 16174
rect 18076 16125 18099 16159
rect 18099 16125 18133 16159
rect 18133 16125 18144 16159
rect 18076 16112 18144 16125
rect 18666 16157 18734 16174
rect 18666 16123 18713 16157
rect 18713 16123 18734 16157
rect 18666 16112 18734 16123
rect 19452 16147 19520 16164
rect 19452 16113 19481 16147
rect 19481 16113 19515 16147
rect 19515 16113 19520 16147
rect 19452 16102 19520 16113
rect 20332 16149 20400 16164
rect 20332 16115 20355 16149
rect 20355 16115 20389 16149
rect 20389 16115 20400 16149
rect 20332 16102 20400 16115
rect 21430 16151 21498 16168
rect 21430 16117 21477 16151
rect 21477 16117 21498 16151
rect 21430 16106 21498 16117
rect 22216 16141 22284 16158
rect 22216 16107 22245 16141
rect 22245 16107 22279 16141
rect 22279 16107 22284 16141
rect 22216 16096 22284 16107
rect 23096 16143 23164 16158
rect 23096 16109 23119 16143
rect 23119 16109 23153 16143
rect 23153 16109 23164 16143
rect 23096 16096 23164 16109
rect 24400 14849 24462 14870
rect 24400 14815 24433 14849
rect 24433 14815 24462 14849
rect 24400 14810 24462 14815
rect 10660 14658 10728 14675
rect 11216 14287 11284 14298
rect 11216 14253 11271 14287
rect 11271 14253 11284 14287
rect 11216 14236 11284 14253
rect 24144 14662 24196 14714
rect 12782 14271 12850 14288
rect 12782 14237 12801 14271
rect 12801 14237 12835 14271
rect 12835 14237 12850 14271
rect 12782 14226 12850 14237
rect 24452 14552 24504 14564
rect 24452 14518 24456 14552
rect 24456 14518 24492 14552
rect 24492 14518 24504 14552
rect 24452 14512 24504 14518
rect 24552 14554 24556 14578
rect 24556 14554 24592 14578
rect 24592 14554 24604 14578
rect 24552 14526 24604 14554
rect 24698 14562 24750 14602
rect 24698 14550 24712 14562
rect 24712 14550 24746 14562
rect 24746 14550 24750 14562
rect 23992 14305 24054 14318
rect 23992 14271 24007 14305
rect 24007 14271 24054 14305
rect 23992 14258 24054 14271
rect 6196 13066 6248 13082
rect 6196 13032 6232 13066
rect 6232 13032 6248 13066
rect 6196 13028 6248 13032
rect 4990 12827 5062 12844
rect 4990 12793 4993 12827
rect 4993 12793 5051 12827
rect 5051 12793 5062 12827
rect 4990 12778 5062 12793
rect 4634 12627 4708 12642
rect 4634 12593 4689 12627
rect 4689 12593 4708 12627
rect 4634 12576 4708 12593
rect 5006 12322 5068 12390
rect 10164 13308 10226 13360
rect 10878 13884 10930 13894
rect 10878 13850 10886 13884
rect 10886 13850 10920 13884
rect 10920 13850 10930 13884
rect 10878 13842 10930 13850
rect 10976 13924 11028 13934
rect 10976 13890 10984 13924
rect 10984 13890 11018 13924
rect 11018 13890 11028 13924
rect 10976 13882 11028 13890
rect 11074 13834 11126 13890
rect 11694 13913 11762 13922
rect 11694 13879 11723 13913
rect 11723 13879 11762 13913
rect 11694 13860 11762 13879
rect 12518 13886 12570 13940
rect 12732 13964 12812 13984
rect 12732 13922 12746 13964
rect 12746 13922 12796 13964
rect 12796 13922 12812 13964
rect 12732 13908 12812 13922
rect 10728 13743 10796 13758
rect 10728 13709 10753 13743
rect 10753 13709 10796 13743
rect 10728 13696 10796 13709
rect 12522 13680 12590 13742
rect 10850 13445 10918 13454
rect 10850 13411 10877 13445
rect 10877 13411 10918 13445
rect 10850 13394 10918 13411
rect 11006 13338 11060 13342
rect 11006 13302 11012 13338
rect 11012 13302 11048 13338
rect 11048 13302 11060 13338
rect 11006 13290 11060 13302
rect 12002 13369 12070 13382
rect 12002 13335 12057 13369
rect 12057 13335 12070 13369
rect 12002 13320 12070 13335
rect 5996 12897 6064 12916
rect 5996 12863 6011 12897
rect 6011 12863 6064 12897
rect 5996 12856 6064 12863
rect 11062 13070 11114 13086
rect 11062 13036 11098 13070
rect 11098 13036 11114 13070
rect 11062 13032 11114 13036
rect 9856 12831 9928 12848
rect 9856 12797 9859 12831
rect 9859 12797 9917 12831
rect 9917 12797 9928 12831
rect 9856 12782 9928 12797
rect 9500 12631 9574 12646
rect 9500 12597 9555 12631
rect 9555 12597 9574 12631
rect 9500 12580 9574 12597
rect 6280 12421 6348 12432
rect 6280 12387 6283 12421
rect 6283 12387 6341 12421
rect 6341 12387 6348 12421
rect 6280 12370 6348 12387
rect 9872 12326 9934 12394
rect 6340 12196 6392 12208
rect 6340 12162 6346 12196
rect 6346 12162 6380 12196
rect 6380 12162 6392 12196
rect 6340 12156 6392 12162
rect 4906 12083 4980 12100
rect 4906 12049 4907 12083
rect 4907 12049 4965 12083
rect 4965 12049 4980 12083
rect 4906 12034 4980 12049
rect 10862 12901 10930 12920
rect 10862 12867 10877 12901
rect 10877 12867 10930 12901
rect 10862 12860 10930 12867
rect 11146 12425 11214 12436
rect 11146 12391 11149 12425
rect 11149 12391 11207 12425
rect 11207 12391 11214 12425
rect 11146 12374 11214 12391
rect 11206 12200 11258 12212
rect 11206 12166 11212 12200
rect 11212 12166 11246 12200
rect 11246 12166 11258 12200
rect 11206 12160 11258 12166
rect 6150 12110 6202 12118
rect 6150 12076 6158 12110
rect 6158 12076 6194 12110
rect 6194 12076 6202 12110
rect 6150 12066 6202 12076
rect 9772 12087 9846 12104
rect 9772 12053 9773 12087
rect 9773 12053 9831 12087
rect 9831 12053 9846 12087
rect 4560 11807 4640 11820
rect 4560 11773 4601 11807
rect 4601 11773 4635 11807
rect 4635 11773 4640 11807
rect 4560 11756 4640 11773
rect 9772 12038 9846 12053
rect 11016 12114 11068 12122
rect 11016 12080 11024 12114
rect 11024 12080 11060 12114
rect 11060 12080 11068 12114
rect 11016 12070 11068 12080
rect 6002 11877 6070 11892
rect 6002 11843 6007 11877
rect 6007 11843 6065 11877
rect 6065 11843 6070 11877
rect 6002 11830 6070 11843
rect 9426 11811 9506 11824
rect 9426 11777 9467 11811
rect 9467 11777 9501 11811
rect 9501 11777 9506 11811
rect 9426 11760 9506 11777
rect 10868 11881 10936 11896
rect 10868 11847 10873 11881
rect 10873 11847 10931 11881
rect 10931 11847 10936 11881
rect 10868 11834 10936 11847
rect 4994 11263 5074 11278
rect 4994 11229 5003 11263
rect 5003 11229 5061 11263
rect 5061 11229 5074 11263
rect 4994 11214 5074 11229
rect 9860 11267 9940 11282
rect 9860 11233 9869 11267
rect 9869 11233 9927 11267
rect 9927 11233 9940 11267
rect 9860 11218 9940 11233
rect 4626 11063 4706 11074
rect 4626 11029 4641 11063
rect 4641 11029 4699 11063
rect 4699 11029 4706 11063
rect 4626 11010 4706 11029
rect 9492 11067 9572 11078
rect 9492 11033 9507 11067
rect 9507 11033 9565 11067
rect 9565 11033 9572 11067
rect 9492 11014 9572 11033
rect 5054 10676 5108 10732
rect 9920 10680 9974 10736
rect 4904 10519 4984 10540
rect 4904 10485 4917 10519
rect 4917 10485 4975 10519
rect 4975 10485 4984 10519
rect 4904 10476 4984 10485
rect 9770 10523 9850 10544
rect 9770 10489 9783 10523
rect 9783 10489 9841 10523
rect 9841 10489 9850 10523
rect 9770 10480 9850 10489
rect 6226 6617 6282 6638
rect 6226 6583 6233 6617
rect 6233 6583 6267 6617
rect 6267 6583 6282 6617
rect 6226 6580 6282 6583
rect 6168 6382 6220 6390
rect 6168 6348 6178 6382
rect 6178 6348 6212 6382
rect 6212 6348 6220 6382
rect 6168 6338 6220 6348
rect 6268 6384 6320 6396
rect 6268 6350 6274 6384
rect 6274 6350 6308 6384
rect 6308 6350 6320 6384
rect 6268 6344 6320 6350
rect 6170 6073 6226 6088
rect 6170 6039 6175 6073
rect 6175 6039 6226 6073
rect 6170 6030 6226 6039
rect 10406 5985 10464 6002
rect 10774 5985 10832 6000
rect 10406 5951 10415 5985
rect 10415 5951 10449 5985
rect 10449 5951 10464 5985
rect 10774 5951 10783 5985
rect 10783 5951 10817 5985
rect 10817 5951 10832 5985
rect 10406 5940 10464 5951
rect 10774 5936 10832 5951
rect 12796 5973 12852 5986
rect 12796 5939 12845 5973
rect 12845 5939 12852 5973
rect 12796 5928 12852 5939
rect 14754 5981 14810 5994
rect 14754 5947 14803 5981
rect 14803 5947 14810 5981
rect 14754 5936 14810 5947
rect 16748 5987 16804 6000
rect 16748 5953 16797 5987
rect 16797 5953 16804 5987
rect 16748 5942 16804 5953
rect 2564 5565 2620 5578
rect 2564 5531 2601 5565
rect 2601 5531 2620 5565
rect 2564 5520 2620 5531
rect 4686 5557 4742 5570
rect 4686 5523 4735 5557
rect 4735 5523 4742 5557
rect 4686 5512 4742 5523
rect 6638 5557 6694 5570
rect 6638 5523 6687 5557
rect 6687 5523 6694 5557
rect 6638 5512 6694 5523
rect 8640 5563 8696 5576
rect 8640 5529 8689 5563
rect 8689 5529 8696 5563
rect 10410 5614 10462 5618
rect 10410 5580 10418 5614
rect 10418 5580 10452 5614
rect 10452 5580 10462 5614
rect 10410 5566 10462 5580
rect 8640 5518 8696 5529
rect 11214 5441 11270 5452
rect 11214 5407 11243 5441
rect 11243 5407 11270 5441
rect 11214 5394 11270 5407
rect 12800 5429 12856 5440
rect 12800 5395 12845 5429
rect 12845 5395 12856 5429
rect 12800 5382 12856 5395
rect 14758 5437 14814 5448
rect 14758 5403 14803 5437
rect 14803 5403 14814 5437
rect 14758 5390 14814 5403
rect 16752 5443 16808 5454
rect 16752 5409 16797 5443
rect 16797 5409 16808 5443
rect 16752 5396 16808 5409
rect 18726 5413 18784 5428
rect 18726 5379 18733 5413
rect 18733 5379 18784 5413
rect 18726 5364 18784 5379
rect 2228 5194 2280 5198
rect 2228 5160 2236 5194
rect 2236 5160 2270 5194
rect 2270 5160 2280 5194
rect 2228 5146 2280 5160
rect 10188 5111 10244 5120
rect 10188 5077 10201 5111
rect 10201 5077 10244 5111
rect 10188 5062 10244 5077
rect 2584 5021 2640 5040
rect 2584 4987 2601 5021
rect 2601 4987 2635 5021
rect 2635 4987 2640 5021
rect 2584 4982 2640 4987
rect 4690 5013 4746 5024
rect 4690 4979 4735 5013
rect 4735 4979 4746 5013
rect 4690 4966 4746 4979
rect 6642 5013 6698 5024
rect 6642 4979 6687 5013
rect 6687 4979 6698 5013
rect 6642 4966 6698 4979
rect 13032 5067 13088 5080
rect 8644 5019 8700 5030
rect 8644 4985 8689 5019
rect 8689 4985 8700 5019
rect 8644 4972 8700 4985
rect 13032 5033 13081 5067
rect 13081 5033 13088 5067
rect 13032 5022 13088 5033
rect 15034 5061 15090 5074
rect 15034 5027 15083 5061
rect 15083 5027 15090 5061
rect 15034 5016 15090 5027
rect 10438 4740 10490 4744
rect 10438 4706 10446 4740
rect 10446 4706 10480 4740
rect 10480 4706 10490 4740
rect 10438 4692 10490 4706
rect 17056 5043 17112 5056
rect 17056 5009 17105 5043
rect 17105 5009 17112 5043
rect 17056 4998 17112 5009
rect 19056 5042 19108 5050
rect 19056 5004 19064 5042
rect 19064 5004 19102 5042
rect 19102 5004 19108 5042
rect 19056 4998 19108 5004
rect 10788 4567 10844 4580
rect 10440 4533 10443 4566
rect 10443 4533 10477 4566
rect 10477 4533 10492 4566
rect 10788 4533 10811 4567
rect 10811 4533 10844 4567
rect 10440 4512 10492 4533
rect 10788 4522 10844 4533
rect 13036 4523 13092 4534
rect 13036 4489 13081 4523
rect 13081 4489 13092 4523
rect 13036 4476 13092 4489
rect 18720 4869 18778 4880
rect 18720 4835 18733 4869
rect 18733 4835 18778 4869
rect 18720 4816 18778 4835
rect 15038 4517 15094 4528
rect 15038 4483 15083 4517
rect 15083 4483 15094 4517
rect 15038 4470 15094 4483
rect 17060 4499 17116 4510
rect 17060 4465 17105 4499
rect 17105 4465 17116 4499
rect 17060 4452 17116 4465
rect 6194 3357 6254 3382
rect 6194 3323 6203 3357
rect 6203 3323 6237 3357
rect 6237 3323 6254 3357
rect 6194 3320 6254 3323
rect 6138 3122 6190 3130
rect 6138 3088 6148 3122
rect 6148 3088 6182 3122
rect 6182 3088 6190 3122
rect 6138 3078 6190 3088
rect 6238 3124 6290 3136
rect 6238 3090 6244 3124
rect 6244 3090 6278 3124
rect 6278 3090 6290 3124
rect 6238 3084 6290 3090
rect 6176 2813 6236 2828
rect 6176 2779 6203 2813
rect 6203 2779 6236 2813
rect 6176 2766 6236 2779
rect 2604 2305 2660 2318
rect 2604 2271 2605 2305
rect 2605 2271 2660 2305
rect 2604 2260 2660 2271
rect 4592 2301 4648 2314
rect 4592 2267 4641 2301
rect 4641 2267 4648 2301
rect 4592 2256 4648 2267
rect 6544 2301 6600 2314
rect 6544 2267 6593 2301
rect 6593 2267 6600 2301
rect 6544 2256 6600 2267
rect 8546 2307 8602 2320
rect 8546 2273 8595 2307
rect 8595 2273 8602 2307
rect 8546 2262 8602 2273
rect 10498 2307 10554 2320
rect 10498 2273 10547 2307
rect 10547 2273 10554 2307
rect 10498 2262 10554 2273
rect 12490 2307 12546 2320
rect 12490 2273 12539 2307
rect 12539 2273 12546 2307
rect 12490 2262 12546 2273
rect 14442 2307 14498 2320
rect 14442 2273 14491 2307
rect 14491 2273 14498 2307
rect 14442 2262 14498 2273
rect 16506 2307 16562 2320
rect 16506 2273 16555 2307
rect 16555 2273 16562 2307
rect 16506 2262 16562 2273
rect 2198 1934 2250 1938
rect 2198 1900 2206 1934
rect 2206 1900 2240 1934
rect 2240 1900 2250 1934
rect 2198 1886 2250 1900
rect 17402 1876 17454 1930
rect 2604 1761 2656 1778
rect 2604 1727 2605 1761
rect 2605 1727 2656 1761
rect 2604 1720 2656 1727
rect 4596 1757 4652 1768
rect 4596 1723 4641 1757
rect 4641 1723 4652 1757
rect 6548 1757 6604 1768
rect 4596 1710 4652 1723
rect 6548 1723 6593 1757
rect 6593 1723 6604 1757
rect 6548 1710 6604 1723
rect 8550 1763 8606 1774
rect 8550 1729 8595 1763
rect 8595 1729 8606 1763
rect 8550 1716 8606 1729
rect 10502 1763 10558 1774
rect 10502 1729 10547 1763
rect 10547 1729 10558 1763
rect 10502 1716 10558 1729
rect 12494 1763 12550 1774
rect 12494 1729 12539 1763
rect 12539 1729 12550 1763
rect 12494 1716 12550 1729
rect 14446 1763 14502 1774
rect 14446 1729 14491 1763
rect 14491 1729 14502 1763
rect 16510 1763 16566 1774
rect 14446 1716 14502 1729
rect 16510 1729 16555 1763
rect 16555 1729 16566 1763
rect 16510 1716 16566 1729
<< metal2 >>
rect 18590 44096 19128 44168
rect 18590 43898 18768 44096
rect 18962 43898 19128 44096
rect 18590 43828 19128 43898
rect 18554 42820 18644 43002
rect 18554 42762 18562 42820
rect 18624 42762 18644 42820
rect 18554 42576 18644 42762
rect 19118 42782 19208 42956
rect 19118 42724 19124 42782
rect 19186 42724 19208 42782
rect 19118 42530 19208 42724
rect 18530 40948 18620 41118
rect 18530 40890 18540 40948
rect 18602 40890 18620 40948
rect 18530 40692 18620 40890
rect 19090 40940 19180 41096
rect 19090 40882 19106 40940
rect 19168 40882 19180 40940
rect 19090 40670 19180 40882
rect 18548 39320 18638 39512
rect 18548 39262 18564 39320
rect 18626 39262 18638 39320
rect 18548 39086 18638 39262
rect 19092 39316 19182 39484
rect 19092 39258 19106 39316
rect 19168 39258 19182 39316
rect 19092 39058 19182 39258
rect 18558 38124 18648 38298
rect 18558 38066 18572 38124
rect 18634 38066 18648 38124
rect 18558 37872 18648 38066
rect 19106 38140 19196 38320
rect 19106 38082 19122 38140
rect 19184 38082 19196 38140
rect 19106 37894 19196 38082
rect 18568 37054 18658 37240
rect 18568 36996 18580 37054
rect 18642 36996 18658 37054
rect 18568 36814 18658 36996
rect 19114 37044 19204 37230
rect 19114 36986 19128 37044
rect 19190 36986 19204 37044
rect 19114 36804 19204 36986
rect 19120 36284 19218 36320
rect 18574 36256 18670 36272
rect 18574 36200 18598 36256
rect 18656 36200 18670 36256
rect 18574 36178 18670 36200
rect 19120 36228 19142 36284
rect 19200 36228 19218 36284
rect 19120 36180 19218 36228
rect 18576 34132 18704 34328
rect 18576 34066 18596 34132
rect 18684 34066 18704 34132
rect 18576 33906 18704 34066
rect 19140 34144 19268 34322
rect 19140 34142 19182 34144
rect 19140 34076 19160 34142
rect 19248 34078 19268 34144
rect 19226 34076 19268 34078
rect 19140 33900 19268 34076
rect 18576 31850 18704 32046
rect 18576 31784 18596 31850
rect 18684 31784 18704 31850
rect 18576 31624 18704 31784
rect 19140 31862 19268 32040
rect 19140 31860 19182 31862
rect 19140 31794 19160 31860
rect 19248 31796 19268 31862
rect 19226 31794 19268 31796
rect 19140 31618 19268 31794
rect 18580 29604 18708 29800
rect 18580 29538 18600 29604
rect 18688 29538 18708 29604
rect 18580 29378 18708 29538
rect 19144 29616 19272 29794
rect 19144 29614 19186 29616
rect 19144 29548 19164 29614
rect 19252 29550 19272 29616
rect 19230 29548 19272 29550
rect 19144 29372 19272 29548
rect 18572 27418 18700 27614
rect 18572 27352 18592 27418
rect 18680 27352 18700 27418
rect 18572 27192 18700 27352
rect 19136 27430 19264 27608
rect 19136 27428 19178 27430
rect 19136 27362 19156 27428
rect 19244 27364 19264 27430
rect 19222 27362 19264 27364
rect 19136 27186 19264 27362
rect 18576 25172 18704 25368
rect 18576 25106 18596 25172
rect 18684 25106 18704 25172
rect 18576 24946 18704 25106
rect 19140 25184 19268 25362
rect 19140 25182 19182 25184
rect 19140 25116 19160 25182
rect 19248 25118 19268 25184
rect 19226 25116 19268 25118
rect 19140 24940 19268 25116
rect 8376 23422 8798 23442
rect 8376 23334 8536 23422
rect 8602 23334 8798 23422
rect 8376 23314 8798 23334
rect 10622 23426 11044 23446
rect 10622 23338 10782 23426
rect 10848 23338 11044 23426
rect 10622 23318 11044 23338
rect 12808 23418 13230 23438
rect 12808 23330 12968 23418
rect 13034 23330 13230 23418
rect 12808 23310 13230 23330
rect 15054 23422 15476 23442
rect 15054 23334 15214 23422
rect 15280 23334 15476 23422
rect 15054 23314 15476 23334
rect 17336 23422 17758 23442
rect 17336 23334 17496 23422
rect 17562 23334 17758 23422
rect 17336 23314 17758 23334
rect 8370 22858 8792 22878
rect 8370 22792 8546 22858
rect 8612 22836 8792 22858
rect 8370 22770 8548 22792
rect 8614 22770 8792 22836
rect 8370 22750 8792 22770
rect 10616 22862 11038 22882
rect 10616 22796 10792 22862
rect 10858 22840 11038 22862
rect 10616 22774 10794 22796
rect 10860 22774 11038 22840
rect 10616 22754 11038 22774
rect 12802 22854 13224 22874
rect 12802 22788 12978 22854
rect 13044 22832 13224 22854
rect 12802 22766 12980 22788
rect 13046 22766 13224 22832
rect 12802 22746 13224 22766
rect 15048 22858 15470 22878
rect 15048 22792 15224 22858
rect 15290 22836 15470 22858
rect 15048 22770 15226 22792
rect 15292 22770 15470 22836
rect 15048 22750 15470 22770
rect 17330 22858 17752 22878
rect 17330 22792 17506 22858
rect 17572 22836 17752 22858
rect 17330 22770 17508 22792
rect 17574 22770 17752 22836
rect 17330 22750 17752 22770
rect 9430 17822 9706 17844
rect 9430 17762 9540 17822
rect 9600 17762 9706 17822
rect 9430 17746 9706 17762
rect 16391 17714 16603 17732
rect 15609 17674 15821 17692
rect 15609 17612 15683 17674
rect 15751 17612 15821 17674
rect 16391 17652 16455 17714
rect 16523 17652 16603 17714
rect 16391 17640 16603 17652
rect 17261 17714 17473 17732
rect 17261 17652 17335 17714
rect 17403 17652 17473 17714
rect 17261 17640 17473 17652
rect 18051 17704 18263 17724
rect 18051 17642 18121 17704
rect 18189 17642 18263 17704
rect 18051 17632 18263 17642
rect 19155 17708 19367 17726
rect 19155 17646 19219 17708
rect 19287 17646 19367 17708
rect 19155 17634 19367 17646
rect 20025 17708 20237 17726
rect 20025 17646 20099 17708
rect 20167 17646 20237 17708
rect 20025 17634 20237 17646
rect 20815 17698 21027 17718
rect 20815 17636 20885 17698
rect 20953 17636 21027 17698
rect 20815 17626 21027 17636
rect 21411 17698 21623 17716
rect 21411 17636 21475 17698
rect 21543 17636 21623 17698
rect 21411 17624 21623 17636
rect 22281 17698 22493 17716
rect 22281 17636 22355 17698
rect 22423 17636 22493 17698
rect 22281 17624 22493 17636
rect 23071 17688 23283 17708
rect 23071 17626 23141 17688
rect 23209 17626 23283 17688
rect 23071 17616 23283 17626
rect 15609 17600 15821 17612
rect 6463 17587 6545 17588
rect 6463 17586 6759 17587
rect 6463 17576 6760 17586
rect 6463 17505 6646 17576
rect 4472 16624 4732 16636
rect 4472 16614 4590 16624
rect 4472 16558 4552 16614
rect 4642 16570 4732 16624
rect 4608 16558 4732 16570
rect 4472 16536 4732 16558
rect 5946 16406 6148 16438
rect 5946 16340 6006 16406
rect 6076 16340 6148 16406
rect 5946 16312 6148 16340
rect 4886 16076 5106 16090
rect 4886 16020 4976 16076
rect 5034 16020 5106 16076
rect 4886 15994 5106 16020
rect 4562 15874 4938 15880
rect 4562 15814 4746 15874
rect 4808 15814 4938 15874
rect 4562 15792 4938 15814
rect 4958 15502 5066 15510
rect 4958 15448 4976 15502
rect 5030 15472 5066 15502
rect 5030 15448 5458 15472
rect 4958 15436 5458 15448
rect 4836 15332 5028 15350
rect 4836 15270 4898 15332
rect 4966 15270 5028 15332
rect 4836 15254 5028 15270
rect 4476 15052 4750 15070
rect 4476 14986 4582 15052
rect 4648 14986 4750 15052
rect 4476 14978 4750 14986
rect 4946 14508 5118 14524
rect 4946 14442 5012 14508
rect 5078 14442 5118 14508
rect 4946 14434 5118 14442
rect 4576 14314 4870 14320
rect 4576 14244 4682 14314
rect 4754 14244 4870 14314
rect 4576 14232 4870 14244
rect 5422 14098 5458 15436
rect 5748 14716 5908 14736
rect 5748 14654 5794 14716
rect 5862 14654 5908 14716
rect 5748 14640 5908 14654
rect 6010 14510 6078 16312
rect 6463 15424 6545 17505
rect 6604 17504 6646 17505
rect 6722 17504 6760 17576
rect 6604 17498 6760 17504
rect 9432 17278 9706 17302
rect 9432 17218 9536 17278
rect 9594 17218 9706 17278
rect 9432 17202 9706 17218
rect 16379 17172 16591 17186
rect 15619 17134 15831 17146
rect 15619 17072 15691 17134
rect 15759 17072 15831 17134
rect 16379 17110 16453 17172
rect 16521 17110 16591 17172
rect 16379 17094 16591 17110
rect 17271 17174 17483 17186
rect 17271 17112 17343 17174
rect 17411 17112 17483 17174
rect 17271 17094 17483 17112
rect 18041 17166 18253 17180
rect 18041 17104 18101 17166
rect 18169 17104 18253 17166
rect 18041 17088 18253 17104
rect 19143 17166 19355 17180
rect 19143 17104 19217 17166
rect 19285 17104 19355 17166
rect 19143 17088 19355 17104
rect 20035 17168 20247 17180
rect 20035 17106 20107 17168
rect 20175 17106 20247 17168
rect 20035 17088 20247 17106
rect 20805 17160 21017 17174
rect 20805 17098 20865 17160
rect 20933 17098 21017 17160
rect 20805 17082 21017 17098
rect 21399 17156 21611 17170
rect 21399 17094 21473 17156
rect 21541 17094 21611 17156
rect 21399 17078 21611 17094
rect 22291 17158 22503 17170
rect 22291 17096 22363 17158
rect 22431 17096 22503 17158
rect 22291 17078 22503 17096
rect 23061 17150 23273 17164
rect 23061 17088 23121 17150
rect 23189 17088 23273 17150
rect 23061 17072 23273 17088
rect 11401 17054 11483 17055
rect 15619 17054 15831 17072
rect 11400 17042 11506 17054
rect 11400 16986 11414 17042
rect 11474 17033 11506 17042
rect 11474 16986 11507 17033
rect 11400 16812 11507 16986
rect 11329 16730 11507 16812
rect 9338 16628 9598 16640
rect 9338 16618 9456 16628
rect 9338 16562 9418 16618
rect 9508 16574 9598 16628
rect 9474 16562 9598 16574
rect 9338 16540 9598 16562
rect 10812 16410 11014 16442
rect 10812 16344 10872 16410
rect 10942 16344 11014 16410
rect 10812 16316 11014 16344
rect 9752 16080 9972 16094
rect 9752 16024 9842 16080
rect 9900 16024 9972 16080
rect 9752 15998 9972 16024
rect 9428 15878 9804 15884
rect 9428 15818 9612 15878
rect 9674 15818 9804 15878
rect 9428 15796 9804 15818
rect 6608 15768 6894 15780
rect 6608 15706 6712 15768
rect 6780 15706 6894 15768
rect 6608 15684 6894 15706
rect 9824 15506 9932 15514
rect 9824 15452 9842 15506
rect 9896 15476 9932 15506
rect 9896 15452 10324 15476
rect 9824 15440 10324 15452
rect 6463 15408 6682 15424
rect 6463 15356 6608 15408
rect 6660 15356 6682 15408
rect 6463 15342 6682 15356
rect 9702 15336 9894 15354
rect 6108 15264 6254 15280
rect 6108 15202 6130 15264
rect 6198 15202 6254 15264
rect 9702 15274 9764 15336
rect 9832 15274 9894 15336
rect 9702 15258 9894 15274
rect 6108 15184 6254 15202
rect 7046 15218 7252 15238
rect 7046 15156 7114 15218
rect 7182 15156 7252 15218
rect 7046 15140 7252 15156
rect 9342 15056 9616 15074
rect 9342 14990 9448 15056
rect 9514 14990 9616 15056
rect 9342 14982 9616 14990
rect 6010 14442 6168 14510
rect 5422 14062 6032 14098
rect 5996 13936 6032 14062
rect 4968 13900 5138 13912
rect 4968 13838 5030 13900
rect 5090 13880 5138 13900
rect 5996 13890 6072 13936
rect 5996 13880 6012 13890
rect 5090 13838 5714 13880
rect 4968 13832 5714 13838
rect 5994 13838 6012 13880
rect 6064 13838 6072 13890
rect 5994 13832 6072 13838
rect 4968 13818 5138 13832
rect 4820 13770 5040 13780
rect 4820 13700 4884 13770
rect 4956 13700 5040 13770
rect 4820 13684 5040 13700
rect 5664 13592 5712 13832
rect 6002 13794 6072 13832
rect 6100 13930 6168 14442
rect 7635 14487 8531 14581
rect 6322 14294 6470 14316
rect 6322 14232 6350 14294
rect 6418 14232 6470 14294
rect 6322 14218 6470 14232
rect 6100 13878 6110 13930
rect 6162 13878 6168 13930
rect 6100 13792 6168 13878
rect 6201 13886 6275 13985
rect 7635 13974 7729 14487
rect 7840 14284 8072 14296
rect 7840 14222 7916 14284
rect 7984 14222 8072 14284
rect 7840 14204 8072 14222
rect 7838 13980 7976 13992
rect 6201 13830 6208 13886
rect 6260 13830 6275 13886
rect 6794 13918 6946 13938
rect 6794 13856 6828 13918
rect 6896 13856 6946 13918
rect 7635 13936 7806 13974
rect 7635 13882 7652 13936
rect 7704 13882 7806 13936
rect 7838 13904 7866 13980
rect 7946 13904 7976 13980
rect 7838 13890 7976 13904
rect 7635 13857 7806 13882
rect 7724 13856 7806 13857
rect 6794 13842 6946 13856
rect 6201 13801 6275 13830
rect 5824 13754 5974 13770
rect 5824 13692 5862 13754
rect 5930 13692 5974 13754
rect 6201 13727 6343 13801
rect 5824 13672 5974 13692
rect 5664 13544 6174 13592
rect 5950 13450 6084 13470
rect 4468 13384 4738 13396
rect 4468 13318 4576 13384
rect 4648 13318 4738 13384
rect 5950 13390 5984 13450
rect 6052 13390 6084 13450
rect 5950 13378 6084 13390
rect 6126 13372 6174 13544
rect 5360 13366 5766 13368
rect 4468 13310 4738 13318
rect 5290 13356 5766 13366
rect 5290 13304 5298 13356
rect 5360 13304 5766 13356
rect 5290 13296 5766 13304
rect 5694 13170 5766 13296
rect 6120 13338 6218 13372
rect 6120 13286 6140 13338
rect 6194 13286 6218 13338
rect 6120 13268 6218 13286
rect 6269 13172 6343 13727
rect 7642 13738 7744 13754
rect 7642 13676 7656 13738
rect 7724 13676 7744 13738
rect 7642 13658 7744 13676
rect 7858 13656 7926 13890
rect 7838 13654 7926 13656
rect 7778 13586 7926 13654
rect 7096 13378 7248 13396
rect 7096 13316 7136 13378
rect 7204 13316 7248 13378
rect 7096 13300 7248 13316
rect 6140 13170 6343 13172
rect 5694 13098 6343 13170
rect 6186 13082 6258 13098
rect 6186 13028 6196 13082
rect 6248 13028 6258 13082
rect 6186 12944 6258 13028
rect 5948 12916 6100 12928
rect 5948 12856 5996 12916
rect 6064 12856 6100 12916
rect 4922 12844 5112 12854
rect 4922 12778 4990 12844
rect 5062 12778 5112 12844
rect 5948 12834 6100 12856
rect 4922 12766 5112 12778
rect 4574 12642 4780 12654
rect 4574 12576 4634 12642
rect 4708 12576 4780 12642
rect 4574 12560 4780 12576
rect 6230 12432 6402 12452
rect 4960 12390 5110 12404
rect 4960 12322 5006 12390
rect 5068 12338 5110 12390
rect 6230 12370 6280 12432
rect 6348 12370 6402 12432
rect 6230 12356 6402 12370
rect 5068 12322 6190 12338
rect 4960 12306 6190 12322
rect 6158 12126 6190 12306
rect 7778 12218 7846 13586
rect 6334 12208 7846 12218
rect 6334 12156 6340 12208
rect 6392 12156 7846 12208
rect 6334 12150 7846 12156
rect 6142 12118 6212 12126
rect 4858 12100 5024 12116
rect 4858 12034 4906 12100
rect 4980 12034 5024 12100
rect 6142 12066 6150 12118
rect 6202 12066 6212 12118
rect 6142 12060 6212 12066
rect 4858 12022 5024 12034
rect 5944 11892 6100 11908
rect 4510 11820 4690 11834
rect 4510 11756 4560 11820
rect 4640 11756 4690 11820
rect 5944 11830 6002 11892
rect 6070 11830 6100 11892
rect 5944 11812 6100 11830
rect 4510 11746 4690 11756
rect 4938 11278 5118 11292
rect 4938 11214 4994 11278
rect 5074 11214 5118 11278
rect 4938 11204 5118 11214
rect 4580 11074 4776 11092
rect 4580 11010 4626 11074
rect 4706 11010 4776 11074
rect 4580 10996 4776 11010
rect 8437 10762 8531 14487
rect 9812 14512 9984 14528
rect 9812 14446 9878 14512
rect 9944 14446 9984 14512
rect 9812 14438 9984 14446
rect 9442 14318 9736 14324
rect 9442 14248 9548 14318
rect 9620 14248 9736 14318
rect 9442 14236 9736 14248
rect 10288 14102 10324 15440
rect 10614 14720 10774 14740
rect 10614 14658 10660 14720
rect 10728 14658 10774 14720
rect 10614 14644 10774 14658
rect 10876 14514 10944 16316
rect 11329 15428 11411 16730
rect 16346 16722 16558 16738
rect 16346 16660 16430 16722
rect 16498 16660 16558 16722
rect 16346 16646 16558 16660
rect 17116 16714 17328 16732
rect 17116 16652 17188 16714
rect 17256 16652 17328 16714
rect 17116 16640 17328 16652
rect 18008 16716 18220 16732
rect 18008 16654 18078 16716
rect 18146 16654 18220 16716
rect 18008 16640 18220 16654
rect 18602 16712 18814 16728
rect 18602 16650 18686 16712
rect 18754 16650 18814 16712
rect 18602 16636 18814 16650
rect 19372 16704 19584 16722
rect 19372 16642 19444 16704
rect 19512 16642 19584 16704
rect 19372 16630 19584 16642
rect 20264 16706 20476 16722
rect 20264 16644 20334 16706
rect 20402 16644 20476 16706
rect 20264 16630 20476 16644
rect 21366 16706 21578 16722
rect 21366 16644 21450 16706
rect 21518 16644 21578 16706
rect 21366 16630 21578 16644
rect 22136 16698 22348 16716
rect 22136 16636 22208 16698
rect 22276 16636 22348 16698
rect 22136 16624 22348 16636
rect 23028 16700 23240 16716
rect 23028 16638 23098 16700
rect 23166 16638 23240 16700
rect 23028 16624 23240 16638
rect 16336 16184 16548 16194
rect 16336 16122 16410 16184
rect 16478 16122 16548 16184
rect 16336 16102 16548 16122
rect 17126 16174 17338 16186
rect 17126 16112 17196 16174
rect 17264 16112 17338 16174
rect 17126 16094 17338 16112
rect 17996 16174 18208 16186
rect 17996 16112 18076 16174
rect 18144 16112 18208 16174
rect 17996 16094 18208 16112
rect 18592 16174 18804 16184
rect 18592 16112 18666 16174
rect 18734 16112 18804 16174
rect 18592 16092 18804 16112
rect 19382 16164 19594 16176
rect 19382 16102 19452 16164
rect 19520 16102 19594 16164
rect 19382 16084 19594 16102
rect 20252 16164 20464 16176
rect 20252 16102 20332 16164
rect 20400 16102 20464 16164
rect 20252 16084 20464 16102
rect 21356 16168 21568 16178
rect 21356 16106 21430 16168
rect 21498 16106 21568 16168
rect 21356 16086 21568 16106
rect 22146 16158 22358 16170
rect 22146 16096 22216 16158
rect 22284 16096 22358 16158
rect 22146 16078 22358 16096
rect 23016 16158 23228 16170
rect 23016 16096 23096 16158
rect 23164 16096 23228 16158
rect 23016 16078 23228 16096
rect 11474 15772 11760 15784
rect 11474 15710 11578 15772
rect 11646 15710 11760 15772
rect 11474 15688 11760 15710
rect 11329 15412 11548 15428
rect 11329 15360 11474 15412
rect 11526 15360 11548 15412
rect 11329 15346 11548 15360
rect 10974 15268 11120 15284
rect 10974 15206 10996 15268
rect 11064 15206 11120 15268
rect 10974 15188 11120 15206
rect 11912 15222 12118 15242
rect 11912 15160 11980 15222
rect 12048 15160 12118 15222
rect 11912 15144 12118 15160
rect 24312 14870 24542 14880
rect 24312 14810 24400 14870
rect 24462 14810 24542 14870
rect 24312 14788 24542 14810
rect 26389 14843 27464 14921
rect 26389 14740 26467 14843
rect 26948 14766 27172 14794
rect 26389 14726 26466 14740
rect 24138 14714 26466 14726
rect 24138 14662 24144 14714
rect 24196 14662 26466 14714
rect 24138 14658 26466 14662
rect 10876 14446 11034 14514
rect 10288 14066 10898 14102
rect 10862 13940 10898 14066
rect 9834 13904 10004 13916
rect 9834 13842 9896 13904
rect 9956 13884 10004 13904
rect 10862 13894 10938 13940
rect 10862 13884 10878 13894
rect 9956 13842 10580 13884
rect 9834 13836 10580 13842
rect 10860 13842 10878 13884
rect 10930 13842 10938 13894
rect 10860 13836 10938 13842
rect 9834 13822 10004 13836
rect 9686 13774 9906 13784
rect 9686 13704 9750 13774
rect 9822 13704 9906 13774
rect 9686 13688 9906 13704
rect 10530 13596 10578 13836
rect 10868 13798 10938 13836
rect 10966 13934 11034 14446
rect 12501 14491 13397 14585
rect 24138 14578 24198 14658
rect 26389 14657 26466 14658
rect 26948 14646 27000 14766
rect 27122 14726 27172 14766
rect 27122 14658 27176 14726
rect 27122 14646 27172 14658
rect 11188 14298 11336 14320
rect 11188 14236 11216 14298
rect 11284 14236 11336 14298
rect 11188 14222 11336 14236
rect 10966 13882 10976 13934
rect 11028 13882 11034 13934
rect 10966 13796 11034 13882
rect 11067 13890 11141 13989
rect 12501 13978 12595 14491
rect 12706 14288 12938 14300
rect 12706 14226 12782 14288
rect 12850 14226 12938 14288
rect 12706 14208 12938 14226
rect 12704 13984 12842 13996
rect 11067 13834 11074 13890
rect 11126 13834 11141 13890
rect 11660 13922 11812 13942
rect 11660 13860 11694 13922
rect 11762 13860 11812 13922
rect 12501 13940 12672 13978
rect 12501 13886 12518 13940
rect 12570 13886 12672 13940
rect 12704 13908 12732 13984
rect 12812 13908 12842 13984
rect 12704 13894 12842 13908
rect 12501 13861 12672 13886
rect 12590 13860 12672 13861
rect 11660 13846 11812 13860
rect 11067 13805 11141 13834
rect 10690 13758 10840 13774
rect 10690 13696 10728 13758
rect 10796 13696 10840 13758
rect 11067 13731 11209 13805
rect 10690 13676 10840 13696
rect 10530 13548 11040 13596
rect 10816 13454 10950 13474
rect 9334 13388 9604 13400
rect 9334 13322 9442 13388
rect 9514 13322 9604 13388
rect 10816 13394 10850 13454
rect 10918 13394 10950 13454
rect 10816 13382 10950 13394
rect 10992 13376 11040 13548
rect 10226 13370 10632 13372
rect 9334 13314 9604 13322
rect 10156 13360 10632 13370
rect 10156 13308 10164 13360
rect 10226 13308 10632 13360
rect 10156 13300 10632 13308
rect 10560 13174 10632 13300
rect 10986 13342 11084 13376
rect 10986 13290 11006 13342
rect 11060 13290 11084 13342
rect 10986 13272 11084 13290
rect 11135 13176 11209 13731
rect 12508 13742 12610 13758
rect 12508 13680 12522 13742
rect 12590 13680 12610 13742
rect 12508 13662 12610 13680
rect 12724 13660 12792 13894
rect 12704 13658 12792 13660
rect 12644 13590 12792 13658
rect 11962 13382 12114 13400
rect 11962 13320 12002 13382
rect 12070 13320 12114 13382
rect 11962 13304 12114 13320
rect 11006 13174 11209 13176
rect 10560 13102 11209 13174
rect 11052 13086 11124 13102
rect 11052 13032 11062 13086
rect 11114 13032 11124 13086
rect 11052 12948 11124 13032
rect 10814 12920 10966 12932
rect 10814 12860 10862 12920
rect 10930 12860 10966 12920
rect 9788 12848 9978 12858
rect 9788 12782 9856 12848
rect 9928 12782 9978 12848
rect 10814 12838 10966 12860
rect 9788 12770 9978 12782
rect 9440 12646 9646 12658
rect 9440 12580 9500 12646
rect 9574 12580 9646 12646
rect 9440 12564 9646 12580
rect 11096 12436 11268 12456
rect 9826 12394 9976 12408
rect 9826 12326 9872 12394
rect 9934 12342 9976 12394
rect 11096 12374 11146 12436
rect 11214 12374 11268 12436
rect 11096 12360 11268 12374
rect 9934 12326 11056 12342
rect 9826 12310 11056 12326
rect 11024 12130 11056 12310
rect 12644 12222 12712 13590
rect 11200 12212 12712 12222
rect 11200 12160 11206 12212
rect 11258 12160 12712 12212
rect 11200 12154 12712 12160
rect 11008 12122 11078 12130
rect 9724 12104 9890 12120
rect 9724 12038 9772 12104
rect 9846 12038 9890 12104
rect 11008 12070 11016 12122
rect 11068 12070 11078 12122
rect 11008 12064 11078 12070
rect 9724 12026 9890 12038
rect 10810 11896 10966 11912
rect 9376 11824 9556 11838
rect 9376 11760 9426 11824
rect 9506 11760 9556 11824
rect 10810 11834 10868 11896
rect 10936 11834 10966 11896
rect 10810 11816 10966 11834
rect 9376 11750 9556 11760
rect 9804 11282 9984 11296
rect 9804 11218 9860 11282
rect 9940 11218 9984 11282
rect 9804 11208 9984 11218
rect 9446 11078 9642 11096
rect 9446 11014 9492 11078
rect 9572 11014 9642 11078
rect 9446 11000 9642 11014
rect 13303 10766 13397 14491
rect 24448 14564 24504 14620
rect 24448 14512 24452 14564
rect 23850 14318 24212 14334
rect 23850 14258 23992 14318
rect 24054 14258 24212 14318
rect 23850 14240 24212 14258
rect 24448 14112 24504 14512
rect 24546 14578 24606 14622
rect 24546 14526 24552 14578
rect 24604 14526 24606 14578
rect 24448 14056 24502 14112
rect 4970 10732 8531 10762
rect 4970 10676 5054 10732
rect 5108 10676 8531 10732
rect 4970 10668 8531 10676
rect 9836 10736 13397 10766
rect 9836 10680 9920 10736
rect 9974 10680 13397 10736
rect 9836 10672 13397 10680
rect 23258 14000 24502 14056
rect 4970 10652 5202 10668
rect 9836 10656 10068 10672
rect 4856 10540 5036 10546
rect 4856 10476 4904 10540
rect 4984 10476 5036 10540
rect 4856 10458 5036 10476
rect 9722 10544 9902 10550
rect 9722 10480 9770 10544
rect 9850 10480 9902 10544
rect 9722 10462 9902 10480
rect 6112 6638 6388 6648
rect 6112 6580 6226 6638
rect 6282 6580 6388 6638
rect 6112 6558 6388 6580
rect 5585 6398 5651 6404
rect 2222 6390 6228 6398
rect 2222 6338 6168 6390
rect 6220 6338 6228 6390
rect 6262 6396 13156 6398
rect 6262 6344 6268 6396
rect 6320 6394 13156 6396
rect 23258 6394 23314 14000
rect 24546 13290 24606 14526
rect 24685 14602 24870 14619
rect 26948 14604 27172 14646
rect 24685 14550 24698 14602
rect 24750 14550 24870 14602
rect 24685 14541 24870 14550
rect 24685 14499 24763 14541
rect 24792 14514 24870 14541
rect 26993 14514 27071 14604
rect 24792 14436 27071 14514
rect 27386 14514 27464 14843
rect 27386 14510 27604 14514
rect 27386 14492 27730 14510
rect 27386 14436 27550 14492
rect 27512 14372 27550 14436
rect 27682 14372 27730 14492
rect 27512 14336 27730 14372
rect 6320 6344 23314 6394
rect 6262 6340 23314 6344
rect 6262 6338 16050 6340
rect 17150 6338 23314 6340
rect 24252 13230 24608 13290
rect 2222 6332 6228 6338
rect 18793 6336 18848 6338
rect 2222 5198 2290 6332
rect 6110 6088 6274 6104
rect 6110 6030 6170 6088
rect 6226 6030 6274 6088
rect 6110 6018 6274 6030
rect 10404 6002 10472 6018
rect 10404 5940 10406 6002
rect 10464 5940 10472 6002
rect 10404 5618 10472 5940
rect 10708 6000 10888 6016
rect 10708 5936 10774 6000
rect 10832 5936 10888 6000
rect 10708 5922 10888 5936
rect 12738 5986 12918 6002
rect 12738 5928 12796 5986
rect 12852 5928 12918 5986
rect 12738 5908 12918 5928
rect 14696 5994 14876 6010
rect 14696 5936 14754 5994
rect 14810 5936 14876 5994
rect 14696 5916 14876 5936
rect 16690 6000 16870 6016
rect 16690 5942 16748 6000
rect 16804 5942 16870 6000
rect 16690 5922 16870 5942
rect 2510 5578 2690 5596
rect 2510 5520 2564 5578
rect 2620 5520 2690 5578
rect 2510 5502 2690 5520
rect 4628 5570 4808 5586
rect 4628 5512 4686 5570
rect 4742 5512 4808 5570
rect 4628 5492 4808 5512
rect 6580 5570 6760 5586
rect 6580 5512 6638 5570
rect 6694 5512 6760 5570
rect 6580 5492 6760 5512
rect 8582 5576 8762 5592
rect 8582 5518 8640 5576
rect 8696 5518 8762 5576
rect 10404 5566 10410 5618
rect 10462 5566 10472 5618
rect 10404 5562 10472 5566
rect 8582 5498 8762 5518
rect 11142 5452 11324 5474
rect 11142 5394 11214 5452
rect 11270 5394 11324 5452
rect 11142 5378 11324 5394
rect 12738 5440 12918 5458
rect 12738 5382 12800 5440
rect 12856 5382 12918 5440
rect 12738 5364 12918 5382
rect 14696 5448 14876 5466
rect 14696 5390 14758 5448
rect 14814 5390 14876 5448
rect 14696 5372 14876 5390
rect 16690 5454 16870 5472
rect 16690 5396 16752 5454
rect 16808 5396 16870 5454
rect 16690 5378 16870 5396
rect 18658 5428 18838 5444
rect 18658 5364 18726 5428
rect 18784 5364 18838 5428
rect 18658 5348 18838 5364
rect 2222 5146 2228 5198
rect 2280 5146 2290 5198
rect 19193 5175 19248 6338
rect 2222 5142 2290 5146
rect 10128 5120 10308 5142
rect 10128 5062 10188 5120
rect 10244 5062 10308 5120
rect 19196 5098 19244 5175
rect 2520 5040 2700 5050
rect 2520 4982 2584 5040
rect 2640 4982 2700 5040
rect 2520 4956 2700 4982
rect 4628 5024 4808 5042
rect 4628 4966 4690 5024
rect 4746 4966 4808 5024
rect 4628 4948 4808 4966
rect 6580 5024 6760 5042
rect 6580 4966 6642 5024
rect 6698 4966 6760 5024
rect 6580 4948 6760 4966
rect 8582 5030 8762 5048
rect 10128 5046 10308 5062
rect 12974 5080 13154 5096
rect 8582 4972 8644 5030
rect 8700 4972 8762 5030
rect 12974 5022 13032 5080
rect 13088 5022 13154 5080
rect 12974 5002 13154 5022
rect 14976 5074 15156 5090
rect 14976 5016 15034 5074
rect 15090 5016 15156 5074
rect 14976 4996 15156 5016
rect 16998 5056 17178 5072
rect 16998 4998 17056 5056
rect 17112 4998 17178 5056
rect 16998 4978 17178 4998
rect 19048 5050 19244 5098
rect 19048 4998 19056 5050
rect 19108 4998 19112 5050
rect 8582 4954 8762 4972
rect 19048 4942 19112 4998
rect 18662 4880 18842 4894
rect 18662 4816 18720 4880
rect 18778 4816 18842 4880
rect 10432 4744 10500 4802
rect 18662 4798 18842 4816
rect 10432 4692 10438 4744
rect 10490 4692 10500 4744
rect 10432 4566 10500 4692
rect 10432 4512 10440 4566
rect 10492 4512 10500 4566
rect 10432 4502 10500 4512
rect 10734 4580 10914 4594
rect 10734 4522 10788 4580
rect 10844 4522 10914 4580
rect 10734 4498 10914 4522
rect 12974 4534 13154 4552
rect 12974 4476 13036 4534
rect 13092 4476 13154 4534
rect 12974 4458 13154 4476
rect 14976 4528 15156 4546
rect 14976 4470 15038 4528
rect 15094 4470 15156 4528
rect 14976 4452 15156 4470
rect 16998 4510 17178 4528
rect 16998 4452 17060 4510
rect 17116 4452 17178 4510
rect 16998 4434 17178 4452
rect 6082 3382 6354 3386
rect 6082 3320 6194 3382
rect 6254 3320 6354 3382
rect 6082 3292 6354 3320
rect 24252 3138 24312 13230
rect 2192 3130 6198 3138
rect 2192 3078 6138 3130
rect 6190 3078 6198 3130
rect 6232 3136 24312 3138
rect 6232 3084 6238 3136
rect 6290 3084 24312 3136
rect 6232 3078 24312 3084
rect 2192 3072 6198 3078
rect 2192 1938 2260 3072
rect 6080 2828 6300 2842
rect 6080 2766 6176 2828
rect 6236 2766 6300 2828
rect 6080 2752 6300 2766
rect 2540 2318 2720 2336
rect 2540 2260 2604 2318
rect 2660 2260 2720 2318
rect 2540 2242 2720 2260
rect 4534 2314 4714 2330
rect 4534 2256 4592 2314
rect 4648 2256 4714 2314
rect 4534 2236 4714 2256
rect 6486 2314 6666 2330
rect 6486 2256 6544 2314
rect 6600 2256 6666 2314
rect 6486 2236 6666 2256
rect 8488 2320 8668 2336
rect 8488 2262 8546 2320
rect 8602 2262 8668 2320
rect 8488 2242 8668 2262
rect 10440 2320 10620 2336
rect 10440 2262 10498 2320
rect 10554 2262 10620 2320
rect 10440 2242 10620 2262
rect 12432 2320 12612 2336
rect 12432 2262 12490 2320
rect 12546 2262 12612 2320
rect 12432 2242 12612 2262
rect 14384 2320 14564 2336
rect 14384 2262 14442 2320
rect 14498 2262 14564 2320
rect 14384 2242 14564 2262
rect 16448 2320 16628 2336
rect 16448 2262 16506 2320
rect 16562 2262 16628 2320
rect 16448 2242 16628 2262
rect 17390 1982 17450 3078
rect 2192 1886 2198 1938
rect 2250 1886 2260 1938
rect 2192 1882 2260 1886
rect 17362 1930 17488 1982
rect 17362 1876 17402 1930
rect 17454 1876 17488 1930
rect 17362 1828 17488 1876
rect 2538 1778 2718 1794
rect 2538 1720 2604 1778
rect 2660 1720 2718 1778
rect 2538 1700 2718 1720
rect 4534 1768 4714 1786
rect 4534 1710 4596 1768
rect 4652 1710 4714 1768
rect 4534 1692 4714 1710
rect 6486 1768 6666 1786
rect 6486 1710 6548 1768
rect 6604 1710 6666 1768
rect 6486 1692 6666 1710
rect 8488 1774 8668 1792
rect 8488 1716 8550 1774
rect 8606 1716 8668 1774
rect 8488 1698 8668 1716
rect 10440 1774 10620 1792
rect 10440 1716 10502 1774
rect 10558 1716 10620 1774
rect 10440 1698 10620 1716
rect 12432 1774 12612 1792
rect 12432 1716 12494 1774
rect 12550 1716 12612 1774
rect 12432 1698 12612 1716
rect 14384 1774 14564 1792
rect 14384 1716 14446 1774
rect 14502 1716 14564 1774
rect 14384 1698 14564 1716
rect 16448 1774 16628 1792
rect 16448 1716 16510 1774
rect 16566 1716 16628 1774
rect 16448 1698 16628 1716
<< via2 >>
rect 18768 43898 18962 44096
rect 18562 42762 18624 42820
rect 19124 42724 19186 42782
rect 18540 40890 18602 40948
rect 19106 40882 19168 40940
rect 18564 39262 18626 39320
rect 19106 39258 19168 39316
rect 18572 38066 18634 38124
rect 19122 38082 19184 38140
rect 18580 36996 18642 37054
rect 19128 36986 19190 37044
rect 18598 36200 18652 36256
rect 18652 36200 18656 36256
rect 19142 36228 19200 36284
rect 18596 34066 18618 34132
rect 18618 34066 18662 34132
rect 19182 34142 19248 34144
rect 19182 34078 19226 34142
rect 19226 34078 19248 34142
rect 18596 31784 18618 31850
rect 18618 31784 18662 31850
rect 19182 31860 19248 31862
rect 19182 31796 19226 31860
rect 19226 31796 19248 31860
rect 18600 29538 18622 29604
rect 18622 29538 18666 29604
rect 19186 29614 19252 29616
rect 19186 29550 19230 29614
rect 19230 29550 19252 29614
rect 18592 27352 18614 27418
rect 18614 27352 18658 27418
rect 19178 27428 19244 27430
rect 19178 27364 19222 27428
rect 19222 27364 19244 27428
rect 18596 25106 18618 25172
rect 18618 25106 18662 25172
rect 19182 25182 19248 25184
rect 19182 25118 19226 25182
rect 19226 25118 19248 25182
rect 8536 23400 8602 23422
rect 8536 23356 8602 23400
rect 10782 23404 10848 23426
rect 10782 23360 10848 23404
rect 12968 23396 13034 23418
rect 12968 23352 13034 23396
rect 15214 23400 15280 23422
rect 15214 23356 15280 23400
rect 17496 23400 17562 23422
rect 17496 23356 17562 23400
rect 8548 22792 8612 22836
rect 8612 22792 8614 22836
rect 8548 22770 8614 22792
rect 10794 22796 10858 22840
rect 10858 22796 10860 22840
rect 10794 22774 10860 22796
rect 12980 22788 13044 22832
rect 13044 22788 13046 22832
rect 12980 22766 13046 22788
rect 15226 22792 15290 22836
rect 15290 22792 15292 22836
rect 15226 22770 15292 22792
rect 17508 22792 17572 22836
rect 17572 22792 17574 22836
rect 17508 22770 17574 22792
rect 9540 17762 9600 17822
rect 15683 17612 15751 17674
rect 16455 17652 16523 17714
rect 17335 17652 17403 17714
rect 18121 17642 18189 17704
rect 19219 17646 19287 17708
rect 20099 17646 20167 17708
rect 20885 17636 20953 17698
rect 21475 17636 21543 17698
rect 22355 17636 22423 17698
rect 23141 17626 23209 17688
rect 4552 16570 4590 16614
rect 4590 16570 4608 16614
rect 4552 16558 4608 16570
rect 4976 16074 5034 16076
rect 4976 16020 5034 16074
rect 4746 15814 4808 15874
rect 4898 15270 4966 15332
rect 4582 14986 4648 15052
rect 5012 14442 5078 14508
rect 4682 14244 4754 14314
rect 5794 14654 5862 14716
rect 9536 17218 9594 17278
rect 15691 17072 15759 17134
rect 16453 17110 16521 17172
rect 17343 17112 17411 17174
rect 18101 17104 18169 17166
rect 19217 17104 19285 17166
rect 20107 17106 20175 17168
rect 20865 17098 20933 17160
rect 21473 17094 21541 17156
rect 22363 17096 22431 17158
rect 23121 17088 23189 17150
rect 9418 16574 9456 16618
rect 9456 16574 9474 16618
rect 9418 16562 9474 16574
rect 9842 16078 9900 16080
rect 9842 16024 9900 16078
rect 9612 15818 9674 15878
rect 6712 15706 6780 15768
rect 6130 15202 6198 15264
rect 9764 15274 9832 15336
rect 7114 15156 7182 15218
rect 9448 14990 9514 15056
rect 4884 13700 4956 13770
rect 6350 14232 6418 14294
rect 7916 14222 7984 14284
rect 6828 13856 6896 13918
rect 5862 13692 5930 13754
rect 4576 13318 4648 13384
rect 5984 13390 6052 13450
rect 7656 13676 7724 13738
rect 7136 13316 7204 13378
rect 5996 12856 6064 12916
rect 4990 12778 5062 12844
rect 4634 12576 4708 12642
rect 6280 12370 6348 12432
rect 4906 12034 4980 12100
rect 4560 11756 4640 11820
rect 6002 11830 6070 11892
rect 4994 11214 5074 11278
rect 4626 11010 4706 11074
rect 9878 14446 9944 14512
rect 9548 14248 9620 14318
rect 10660 14658 10728 14720
rect 16430 16660 16498 16722
rect 17188 16652 17256 16714
rect 18078 16654 18146 16716
rect 18686 16650 18754 16712
rect 19444 16642 19512 16704
rect 20334 16644 20402 16706
rect 21450 16644 21518 16706
rect 22208 16636 22276 16698
rect 23098 16638 23166 16700
rect 16410 16122 16478 16184
rect 17196 16112 17264 16174
rect 18076 16112 18144 16174
rect 18666 16112 18734 16174
rect 19452 16102 19520 16164
rect 20332 16102 20400 16164
rect 21430 16106 21498 16168
rect 22216 16096 22284 16158
rect 23096 16096 23164 16158
rect 11578 15710 11646 15772
rect 10996 15206 11064 15268
rect 11980 15160 12048 15222
rect 24400 14810 24462 14870
rect 9750 13704 9822 13774
rect 27000 14646 27122 14766
rect 11216 14236 11284 14298
rect 12782 14226 12850 14288
rect 11694 13860 11762 13922
rect 10728 13696 10796 13758
rect 9442 13322 9514 13388
rect 10850 13394 10918 13454
rect 12522 13680 12590 13742
rect 12002 13320 12070 13382
rect 10862 12860 10930 12920
rect 9856 12782 9928 12848
rect 9500 12580 9574 12646
rect 11146 12374 11214 12436
rect 9772 12038 9846 12104
rect 9426 11760 9506 11824
rect 10868 11834 10936 11896
rect 9860 11218 9940 11282
rect 9492 11014 9572 11078
rect 23992 14258 24054 14318
rect 4904 10476 4984 10540
rect 9770 10480 9850 10544
rect 6226 6580 6282 6638
rect 27550 14372 27682 14492
rect 6170 6030 6226 6088
rect 10774 5936 10832 6000
rect 12796 5928 12852 5986
rect 14754 5936 14810 5994
rect 16748 5942 16804 6000
rect 2564 5520 2620 5578
rect 4686 5512 4742 5570
rect 6638 5512 6694 5570
rect 8640 5518 8696 5576
rect 11214 5394 11270 5452
rect 12800 5382 12856 5440
rect 14758 5390 14814 5448
rect 16752 5396 16808 5454
rect 18726 5364 18784 5428
rect 10188 5062 10244 5120
rect 2584 4982 2640 5040
rect 4690 4966 4746 5024
rect 6642 4966 6698 5024
rect 8644 4972 8700 5030
rect 13032 5022 13088 5080
rect 15034 5016 15090 5074
rect 17056 4998 17112 5056
rect 18720 4816 18778 4880
rect 10788 4522 10844 4580
rect 13036 4476 13092 4534
rect 15038 4470 15094 4528
rect 17060 4452 17116 4510
rect 6194 3320 6254 3382
rect 6176 2766 6236 2828
rect 2604 2260 2660 2318
rect 4592 2256 4648 2314
rect 6544 2256 6600 2314
rect 8546 2262 8602 2320
rect 10498 2262 10554 2320
rect 12490 2262 12546 2320
rect 14442 2262 14498 2320
rect 16506 2262 16562 2320
rect 2604 1720 2656 1778
rect 2656 1720 2660 1778
rect 4596 1710 4652 1768
rect 6548 1710 6604 1768
rect 8550 1716 8606 1774
rect 10502 1716 10558 1774
rect 12494 1716 12550 1774
rect 14446 1716 14502 1774
rect 16510 1716 16566 1774
<< metal3 >>
rect 18590 44096 19128 44168
rect 18590 43898 18768 44096
rect 18962 43898 19128 44096
rect 18590 43828 19128 43898
rect 17652 43002 18076 43406
rect 17652 42820 18672 43002
rect 19448 42956 19880 43622
rect 17652 42762 18562 42820
rect 18624 42762 18672 42820
rect 17652 42578 18672 42762
rect 19102 42782 19880 42956
rect 19102 42724 19124 42782
rect 19186 42724 19880 42782
rect 17652 41110 18076 42578
rect 19102 42524 19880 42724
rect 18530 41110 18620 41118
rect 17652 40948 18636 41110
rect 19448 41102 19880 42524
rect 19116 41096 19880 41102
rect 17652 40890 18540 40948
rect 18602 40890 18636 40948
rect 17652 40686 18636 40890
rect 19090 40940 19880 41096
rect 19090 40882 19106 40940
rect 19168 40882 19880 40940
rect 17652 39508 18076 40686
rect 19090 40670 19880 40882
rect 17652 39320 18636 39508
rect 19448 39486 19880 40670
rect 19116 39484 19880 39486
rect 17652 39262 18564 39320
rect 18626 39262 18636 39320
rect 17652 39084 18636 39262
rect 19092 39316 19880 39484
rect 19092 39258 19106 39316
rect 19168 39258 19880 39316
rect 17652 38286 18076 39084
rect 19092 39058 19880 39258
rect 19116 39054 19880 39058
rect 19448 38310 19880 39054
rect 18558 38286 18648 38298
rect 17652 38124 18658 38286
rect 17652 38066 18572 38124
rect 18634 38066 18658 38124
rect 17652 37862 18658 38066
rect 19094 38140 19880 38310
rect 19094 38082 19122 38140
rect 19184 38082 19880 38140
rect 19094 37878 19880 38082
rect 17652 37228 18076 37862
rect 17652 37054 18656 37228
rect 19448 37222 19880 37878
rect 17652 36996 18580 37054
rect 18642 36996 18656 37054
rect 17652 36804 18656 36996
rect 19116 37044 19880 37222
rect 19116 36986 19128 37044
rect 19190 36986 19880 37044
rect 17652 36446 18076 36804
rect 19116 36790 19880 36986
rect 19448 36448 19880 36790
rect 17652 36256 18674 36446
rect 17652 36200 18598 36256
rect 18656 36200 18674 36256
rect 17652 36022 18674 36200
rect 19120 36284 19880 36448
rect 19120 36228 19142 36284
rect 19200 36228 19880 36284
rect 17652 34644 18076 36022
rect 19120 36016 19880 36228
rect 17652 34334 18318 34644
rect 19448 34628 19880 36016
rect 17652 34132 18686 34334
rect 19194 34318 19880 34628
rect 17652 34066 18596 34132
rect 18662 34066 18686 34132
rect 17652 33910 18686 34066
rect 19146 34144 19880 34318
rect 19146 34078 19182 34144
rect 19248 34078 19880 34144
rect 17652 33878 18320 33910
rect 19146 33894 19880 34078
rect 17652 33860 18088 33878
rect 19424 33868 19880 33894
rect 17652 32338 18076 33860
rect 17652 32052 18318 32338
rect 19448 32322 19880 33868
rect 17652 31914 18686 32052
rect 19194 32036 19880 32322
rect 17652 31698 17888 31914
rect 18048 31850 18686 31914
rect 18048 31784 18596 31850
rect 18662 31784 18686 31850
rect 18048 31698 18686 31784
rect 17652 31628 18686 31698
rect 19146 31862 19880 32036
rect 19146 31796 19182 31862
rect 19248 31796 19880 31862
rect 17652 31596 18320 31628
rect 19146 31612 19880 31796
rect 17652 30124 18076 31596
rect 17652 29806 18318 30124
rect 19448 30108 19880 31612
rect 17652 29700 18690 29806
rect 19194 29790 19880 30108
rect 17652 29498 17888 29700
rect 18048 29604 18690 29700
rect 18048 29538 18600 29604
rect 18666 29538 18690 29604
rect 18048 29498 18690 29538
rect 17652 29382 18690 29498
rect 19150 29616 19880 29790
rect 19150 29550 19186 29616
rect 19252 29550 19880 29616
rect 17652 27924 18076 29382
rect 19150 29366 19880 29550
rect 17652 27620 18318 27924
rect 19448 27908 19880 29366
rect 17652 27500 18682 27620
rect 19194 27604 19880 27908
rect 17652 27284 17888 27500
rect 18048 27418 18682 27500
rect 18048 27352 18592 27418
rect 18658 27352 18682 27418
rect 18048 27284 18682 27352
rect 17652 27196 18682 27284
rect 19142 27430 19880 27604
rect 19142 27364 19178 27430
rect 19244 27364 19880 27430
rect 17652 27164 18316 27196
rect 19142 27180 19880 27364
rect 17652 25710 18076 27164
rect 19424 27148 19880 27180
rect 17652 25374 18318 25710
rect 19448 25694 19880 27148
rect 17652 25172 18686 25374
rect 19194 25358 19880 25694
rect 17652 25106 18596 25172
rect 18662 25106 18686 25172
rect 17652 24950 18686 25106
rect 19146 25184 19880 25358
rect 19146 25118 19182 25184
rect 19248 25118 19880 25184
rect 17652 24396 18076 24950
rect 19146 24934 19880 25118
rect 228 24272 18076 24396
rect 228 24092 300 24272
rect 488 24092 18076 24272
rect 228 23972 18076 24092
rect 8380 23422 8804 23972
rect 10594 23702 11050 23972
rect 11944 23968 16336 23972
rect 8380 23356 8536 23422
rect 8602 23356 8804 23422
rect 8380 23332 8804 23356
rect 10626 23426 11050 23702
rect 10626 23360 10782 23426
rect 10848 23360 11050 23426
rect 10626 23336 11050 23360
rect 12812 23418 13236 23968
rect 15026 23698 15482 23968
rect 17308 23698 17764 23972
rect 12812 23352 12968 23418
rect 13034 23352 13236 23418
rect 12812 23328 13236 23352
rect 15058 23422 15482 23698
rect 15058 23356 15214 23422
rect 15280 23356 15482 23422
rect 15058 23332 15482 23356
rect 17340 23422 17764 23698
rect 17340 23356 17496 23422
rect 17562 23356 17764 23422
rect 17340 23332 17764 23356
rect 8364 22836 8788 22872
rect 8364 22770 8548 22836
rect 8614 22770 8788 22836
rect 8364 22244 8788 22770
rect 10610 22840 11034 22876
rect 10610 22774 10794 22840
rect 10860 22774 11034 22840
rect 10610 22594 11034 22774
rect 10578 22248 11034 22594
rect 12796 22832 13220 22868
rect 12796 22766 12980 22832
rect 13046 22766 13220 22832
rect 9726 22244 11964 22248
rect 12796 22244 13220 22766
rect 15042 22836 15466 22872
rect 15042 22770 15226 22836
rect 15292 22770 15466 22836
rect 15042 22244 15466 22770
rect 17324 22836 17748 22872
rect 17324 22770 17508 22836
rect 17574 22770 17748 22836
rect 17324 22594 17748 22770
rect 17298 22252 17748 22594
rect 19448 22252 19880 24934
rect 16310 22244 19880 22252
rect 898 22150 19880 22244
rect 898 21970 978 22150
rect 1166 21970 19880 22150
rect 898 21820 19880 21970
rect 814 17848 23871 17936
rect 814 17780 996 17848
rect 1066 17822 23871 17848
rect 1066 17780 9540 17822
rect 814 17762 9540 17780
rect 9600 17762 23871 17822
rect 814 17722 23871 17762
rect 15360 17674 15904 17722
rect 16084 17718 23871 17722
rect 15360 17646 15683 17674
rect 15606 17612 15683 17646
rect 15751 17646 15904 17674
rect 16392 17714 16606 17718
rect 16392 17652 16455 17714
rect 16523 17652 16606 17714
rect 15751 17612 15820 17646
rect 16392 17635 16606 17652
rect 17258 17714 17472 17718
rect 17258 17652 17335 17714
rect 17403 17652 17472 17714
rect 17258 17641 17472 17652
rect 18052 17704 18266 17718
rect 18052 17642 18121 17704
rect 18189 17642 18266 17704
rect 18052 17627 18266 17642
rect 19156 17708 19370 17718
rect 19156 17646 19219 17708
rect 19287 17646 19370 17708
rect 19156 17629 19370 17646
rect 20022 17708 20236 17718
rect 20022 17646 20099 17708
rect 20167 17646 20236 17708
rect 20022 17635 20236 17646
rect 20816 17698 21030 17718
rect 20816 17636 20885 17698
rect 20953 17636 21030 17698
rect 20816 17621 21030 17636
rect 21412 17698 21626 17718
rect 21412 17636 21475 17698
rect 21543 17636 21626 17698
rect 21412 17619 21626 17636
rect 22278 17698 22492 17718
rect 22278 17636 22355 17698
rect 22423 17636 22492 17698
rect 22278 17625 22492 17636
rect 23072 17688 23286 17718
rect 23072 17626 23141 17688
rect 23209 17626 23286 17688
rect 15606 17601 15820 17612
rect 23072 17611 23286 17626
rect 200 17278 13306 17330
rect 200 17218 9536 17278
rect 9594 17218 13306 17278
rect 200 17104 13306 17218
rect 16373 17172 16601 17188
rect 200 16942 322 17104
rect 474 17038 13306 17104
rect 15611 17134 15839 17144
rect 15611 17072 15691 17134
rect 15759 17072 15839 17134
rect 16373 17110 16453 17172
rect 16521 17110 16601 17172
rect 16373 17074 16601 17110
rect 17263 17174 17491 17184
rect 17263 17112 17343 17174
rect 17411 17112 17491 17174
rect 17263 17074 17491 17112
rect 18031 17166 18259 17174
rect 18031 17104 18101 17166
rect 18169 17104 18259 17166
rect 18031 17074 18259 17104
rect 19137 17166 19365 17182
rect 19137 17104 19217 17166
rect 19285 17104 19365 17166
rect 19137 17074 19365 17104
rect 20027 17168 20255 17178
rect 20027 17106 20107 17168
rect 20175 17106 20255 17168
rect 20027 17074 20255 17106
rect 20795 17160 21023 17168
rect 20795 17098 20865 17160
rect 20933 17098 21023 17160
rect 20795 17074 21023 17098
rect 21393 17156 21621 17172
rect 21393 17094 21473 17156
rect 21541 17094 21621 17156
rect 21393 17074 21621 17094
rect 22283 17158 22511 17168
rect 22283 17096 22363 17158
rect 22431 17096 22511 17158
rect 22283 17074 22511 17096
rect 23051 17150 23279 17158
rect 23051 17088 23121 17150
rect 23189 17088 23279 17150
rect 23051 17074 23279 17088
rect 15611 17038 15839 17072
rect 16134 17038 23388 17074
rect 474 16942 23388 17038
rect 200 16810 23388 16942
rect 200 16808 13306 16810
rect 4036 16628 4280 16808
rect 4036 16614 4844 16628
rect 4036 16558 4552 16614
rect 4608 16558 4844 16614
rect 4036 16536 4844 16558
rect 4036 15884 4280 16536
rect 4880 16076 5584 16082
rect 4880 16020 4976 16076
rect 5034 16020 5584 16076
rect 4880 15994 5584 16020
rect 5342 15912 5584 15994
rect 4036 15874 4938 15884
rect 4036 15814 4746 15874
rect 4808 15814 4938 15874
rect 4036 15792 4938 15814
rect 4036 15066 4280 15792
rect 5340 15344 5584 15912
rect 4834 15332 5584 15344
rect 4834 15270 4898 15332
rect 4966 15270 5584 15332
rect 6320 15780 6502 16808
rect 6320 15768 6896 15780
rect 6320 15706 6712 15768
rect 6780 15706 6896 15768
rect 6320 15684 6896 15706
rect 6320 15278 6502 15684
rect 4834 15256 5584 15270
rect 4036 15052 4900 15066
rect 4036 14986 4582 15052
rect 4648 14986 4900 15052
rect 4036 14974 4900 14986
rect 4036 14324 4280 14974
rect 5340 14738 5584 15256
rect 6088 15264 6502 15278
rect 6088 15202 6130 15264
rect 6198 15202 6502 15264
rect 6088 15180 6502 15202
rect 5340 14716 6026 14738
rect 5340 14654 5794 14716
rect 5862 14654 6026 14716
rect 5340 14642 6026 14654
rect 5340 14522 5584 14642
rect 4942 14508 5584 14522
rect 4942 14442 5012 14508
rect 5078 14442 5584 14508
rect 4942 14434 5584 14442
rect 4036 14314 4880 14324
rect 4036 14244 4682 14314
rect 4754 14244 4880 14314
rect 4036 14232 4880 14244
rect 4036 13404 4280 14232
rect 5340 13776 5584 14434
rect 6320 14433 6502 15180
rect 7050 15218 7552 15236
rect 7050 15156 7114 15218
rect 7182 15156 7552 15218
rect 7050 15140 7552 15156
rect 6321 14430 6502 14433
rect 6321 14334 6684 14430
rect 6321 14328 6502 14334
rect 6320 14294 6502 14328
rect 6320 14232 6350 14294
rect 6418 14232 6502 14294
rect 6320 14213 6502 14232
rect 6589 13938 6684 14334
rect 6584 13918 6948 13938
rect 6584 13856 6828 13918
rect 6896 13856 6948 13918
rect 6584 13846 6948 13856
rect 4822 13772 5584 13776
rect 4822 13770 6086 13772
rect 4822 13700 4884 13770
rect 4956 13754 6086 13770
rect 4956 13700 5862 13754
rect 4822 13692 5862 13700
rect 5930 13692 6086 13754
rect 4822 13688 6086 13692
rect 5340 13676 6086 13688
rect 4036 13384 4884 13404
rect 4036 13318 4576 13384
rect 4648 13318 4884 13384
rect 4036 13312 4884 13318
rect 4036 12658 4280 13312
rect 5340 12928 5584 13676
rect 6589 13470 6684 13846
rect 5948 13450 6684 13470
rect 5948 13390 5984 13450
rect 6052 13390 6684 13450
rect 7348 13752 7552 15140
rect 7838 14284 8072 16808
rect 7838 14222 7916 14284
rect 7984 14222 8072 14284
rect 7838 14188 8072 14222
rect 8902 16792 9242 16808
rect 11186 16792 11464 16808
rect 12704 16792 13034 16808
rect 8902 16632 9146 16792
rect 8902 16618 9710 16632
rect 8902 16562 9418 16618
rect 9474 16562 9710 16618
rect 8902 16540 9710 16562
rect 8902 15888 9146 16540
rect 9746 16080 10450 16086
rect 9746 16024 9842 16080
rect 9900 16024 10450 16080
rect 9746 15998 10450 16024
rect 10208 15916 10450 15998
rect 8902 15878 9804 15888
rect 8902 15818 9612 15878
rect 9674 15818 9804 15878
rect 8902 15796 9804 15818
rect 8902 15070 9146 15796
rect 10206 15348 10450 15916
rect 9700 15336 10450 15348
rect 9700 15274 9764 15336
rect 9832 15274 10450 15336
rect 11186 15784 11368 16792
rect 11186 15772 11762 15784
rect 11186 15710 11578 15772
rect 11646 15710 11762 15772
rect 11186 15688 11762 15710
rect 11186 15282 11368 15688
rect 9700 15260 10450 15274
rect 8902 15056 9766 15070
rect 8902 14990 9448 15056
rect 9514 14990 9766 15056
rect 8902 14978 9766 14990
rect 8902 14328 9146 14978
rect 10206 14742 10450 15260
rect 10954 15268 11368 15282
rect 10954 15206 10996 15268
rect 11064 15206 11368 15268
rect 10954 15184 11368 15206
rect 10206 14720 10892 14742
rect 10206 14658 10660 14720
rect 10728 14658 10892 14720
rect 10206 14646 10892 14658
rect 10206 14526 10450 14646
rect 9808 14512 10450 14526
rect 9808 14446 9878 14512
rect 9944 14446 10450 14512
rect 9808 14438 10450 14446
rect 8902 14318 9746 14328
rect 8902 14248 9548 14318
rect 9620 14248 9746 14318
rect 8902 14236 9746 14248
rect 7348 13738 7746 13752
rect 7348 13676 7656 13738
rect 7724 13676 7746 13738
rect 7348 13656 7746 13676
rect 7348 13394 7552 13656
rect 5948 13378 6684 13390
rect 5340 12916 6098 12928
rect 5340 12856 5996 12916
rect 6064 12856 6098 12916
rect 5340 12854 6098 12856
rect 4926 12844 6098 12854
rect 4926 12778 4990 12844
rect 5062 12832 6098 12844
rect 5062 12778 5584 12832
rect 4926 12766 5584 12778
rect 4036 12642 4952 12658
rect 4036 12576 4634 12642
rect 4708 12576 4952 12642
rect 4036 12566 4952 12576
rect 4036 11840 4280 12566
rect 5340 12110 5584 12766
rect 6589 12454 6684 13378
rect 7092 13378 7552 13394
rect 7092 13316 7136 13378
rect 7204 13316 7552 13378
rect 7092 13298 7552 13316
rect 6193 12432 6684 12454
rect 6193 12370 6280 12432
rect 6348 12370 6684 12432
rect 6193 12359 6684 12370
rect 4850 12100 5584 12110
rect 4850 12034 4906 12100
rect 4980 12034 5584 12100
rect 4850 12022 5584 12034
rect 5340 11906 5584 12022
rect 5340 11892 6100 11906
rect 4036 11820 4838 11840
rect 4036 11756 4560 11820
rect 4640 11756 4838 11820
rect 4036 11748 4838 11756
rect 5340 11830 6002 11892
rect 6070 11830 6100 11892
rect 5340 11810 6100 11830
rect 4036 11090 4280 11748
rect 5340 11294 5584 11810
rect 4936 11278 5584 11294
rect 4936 11214 4994 11278
rect 5074 11214 5584 11278
rect 4936 11200 5584 11214
rect 4036 11074 4904 11090
rect 4036 11010 4626 11074
rect 4706 11010 4904 11074
rect 4036 10998 4904 11010
rect 4036 10996 4280 10998
rect 5340 10554 5584 11200
rect 4852 10540 5584 10554
rect 4852 10476 4904 10540
rect 4984 10476 5584 10540
rect 4852 10448 5584 10476
rect 5340 9882 5584 10448
rect 7348 9882 7552 13298
rect 8902 13408 9146 14236
rect 10206 13780 10450 14438
rect 11186 14437 11368 15184
rect 11916 15222 12418 15240
rect 11916 15160 11980 15222
rect 12048 15160 12418 15222
rect 11916 15144 12418 15160
rect 11187 14434 11368 14437
rect 11187 14338 11550 14434
rect 11187 14332 11368 14338
rect 11186 14298 11368 14332
rect 11186 14236 11216 14298
rect 11284 14236 11368 14298
rect 11186 14217 11368 14236
rect 11455 13942 11550 14338
rect 11450 13922 11814 13942
rect 11450 13860 11694 13922
rect 11762 13860 11814 13922
rect 11450 13850 11814 13860
rect 9688 13776 10450 13780
rect 9688 13774 10952 13776
rect 9688 13704 9750 13774
rect 9822 13758 10952 13774
rect 9822 13704 10728 13758
rect 9688 13696 10728 13704
rect 10796 13696 10952 13758
rect 9688 13692 10952 13696
rect 10206 13680 10952 13692
rect 8902 13388 9750 13408
rect 8902 13322 9442 13388
rect 9514 13322 9750 13388
rect 8902 13316 9750 13322
rect 8902 12662 9146 13316
rect 10206 12932 10450 13680
rect 11455 13474 11550 13850
rect 10814 13454 11550 13474
rect 10814 13394 10850 13454
rect 10918 13394 11550 13454
rect 12214 13756 12418 15144
rect 12704 14288 12938 16792
rect 15198 15406 15426 16810
rect 16134 16794 23388 16810
rect 16340 16722 16568 16794
rect 16340 16660 16430 16722
rect 16498 16660 16568 16722
rect 16340 16652 16568 16660
rect 17108 16714 17336 16794
rect 17108 16652 17188 16714
rect 17256 16652 17336 16714
rect 17108 16642 17336 16652
rect 17998 16716 18226 16794
rect 17998 16654 18078 16716
rect 18146 16654 18226 16716
rect 17998 16638 18226 16654
rect 18596 16712 18824 16794
rect 18596 16650 18686 16712
rect 18754 16650 18824 16712
rect 18596 16642 18824 16650
rect 19364 16704 19592 16794
rect 19364 16642 19444 16704
rect 19512 16642 19592 16704
rect 19364 16632 19592 16642
rect 20254 16706 20482 16794
rect 20254 16644 20334 16706
rect 20402 16644 20482 16706
rect 20254 16628 20482 16644
rect 21360 16706 21588 16794
rect 21360 16644 21450 16706
rect 21518 16644 21588 16706
rect 21360 16636 21588 16644
rect 22128 16698 22356 16794
rect 22128 16636 22208 16698
rect 22276 16636 22356 16698
rect 22128 16626 22356 16636
rect 23018 16700 23246 16794
rect 23018 16638 23098 16700
rect 23166 16638 23246 16700
rect 23018 16622 23246 16638
rect 16333 16184 16547 16199
rect 16333 16122 16410 16184
rect 16478 16122 16547 16184
rect 16333 16027 16547 16122
rect 17127 16174 17341 16185
rect 17127 16112 17196 16174
rect 17264 16112 17341 16174
rect 17127 16027 17341 16112
rect 17993 16174 18207 16191
rect 17993 16112 18076 16174
rect 18144 16112 18207 16174
rect 17993 16027 18207 16112
rect 18589 16174 18803 16189
rect 18589 16112 18666 16174
rect 18734 16112 18803 16174
rect 16197 16018 18300 16027
rect 16197 16017 18510 16018
rect 18589 16017 18803 16112
rect 19383 16164 19597 16175
rect 19383 16102 19452 16164
rect 19520 16102 19597 16164
rect 19383 16017 19597 16102
rect 20249 16164 20463 16181
rect 20249 16102 20332 16164
rect 20400 16102 20463 16164
rect 20249 16017 20463 16102
rect 21353 16168 21567 16183
rect 21353 16106 21430 16168
rect 21498 16106 21567 16168
rect 21353 16017 21567 16106
rect 16197 16011 21567 16017
rect 22147 16158 22361 16169
rect 22147 16096 22216 16158
rect 22284 16096 22361 16158
rect 22147 16011 22361 16096
rect 23013 16158 23227 16175
rect 23013 16096 23096 16158
rect 23164 16096 23227 16158
rect 23013 16027 23227 16096
rect 23657 16027 23871 17718
rect 22627 16011 23871 16027
rect 16197 16010 21710 16011
rect 21790 16010 21966 16011
rect 16197 16006 21966 16010
rect 22094 16006 23871 16011
rect 16197 15896 23871 16006
rect 16197 15813 23874 15896
rect 18292 15803 23874 15813
rect 20597 15797 23874 15803
rect 23270 15794 23874 15797
rect 15198 15178 24536 15406
rect 24310 15150 24536 15178
rect 24310 14870 24538 15150
rect 24310 14810 24400 14870
rect 24462 14810 24538 14870
rect 24310 14790 24538 14810
rect 26956 14766 27174 14788
rect 26956 14646 27000 14766
rect 27122 14646 27174 14766
rect 26956 14604 27174 14646
rect 27512 14492 27730 14510
rect 27512 14372 27550 14492
rect 27682 14372 27730 14492
rect 27512 14336 27730 14372
rect 12704 14226 12782 14288
rect 12850 14226 12938 14288
rect 12704 14192 12938 14226
rect 23852 14318 24212 14334
rect 23852 14258 23992 14318
rect 24054 14258 24212 14318
rect 23852 14128 24212 14258
rect 23852 13946 24204 14128
rect 12214 13742 12612 13756
rect 12214 13680 12522 13742
rect 12590 13680 12612 13742
rect 12214 13660 12612 13680
rect 15110 13726 24204 13946
rect 12214 13398 12418 13660
rect 10814 13382 11550 13394
rect 10206 12920 10964 12932
rect 10206 12860 10862 12920
rect 10930 12860 10964 12920
rect 10206 12858 10964 12860
rect 9792 12848 10964 12858
rect 9792 12782 9856 12848
rect 9928 12836 10964 12848
rect 9928 12782 10450 12836
rect 9792 12770 10450 12782
rect 8902 12646 9818 12662
rect 8902 12580 9500 12646
rect 9574 12580 9818 12646
rect 8902 12570 9818 12580
rect 8902 11844 9146 12570
rect 10206 12114 10450 12770
rect 11455 12458 11550 13382
rect 11958 13382 12418 13398
rect 11958 13320 12002 13382
rect 12070 13320 12418 13382
rect 11958 13302 12418 13320
rect 11059 12436 11550 12458
rect 11059 12374 11146 12436
rect 11214 12374 11550 12436
rect 11059 12363 11550 12374
rect 9716 12104 10450 12114
rect 9716 12038 9772 12104
rect 9846 12038 10450 12104
rect 9716 12026 10450 12038
rect 10206 11910 10450 12026
rect 10206 11896 10966 11910
rect 8902 11824 9704 11844
rect 8902 11760 9426 11824
rect 9506 11760 9704 11824
rect 8902 11752 9704 11760
rect 10206 11834 10868 11896
rect 10936 11834 10966 11896
rect 10206 11814 10966 11834
rect 8902 11094 9146 11752
rect 10206 11298 10450 11814
rect 9802 11282 10450 11298
rect 9802 11218 9860 11282
rect 9940 11218 10450 11282
rect 9802 11204 10450 11218
rect 8902 11078 9770 11094
rect 8902 11014 9492 11078
rect 9572 11014 9770 11078
rect 8902 11002 9770 11014
rect 8902 11000 9146 11002
rect 10206 10558 10450 11204
rect 9718 10544 10450 10558
rect 9718 10480 9770 10544
rect 9850 10480 10450 10544
rect 9718 10452 10450 10480
rect 10206 9944 10450 10452
rect 12214 9944 12418 13302
rect 15110 13586 24208 13726
rect 10206 9922 10540 9944
rect 12214 9922 12508 9944
rect 13258 9922 13626 9926
rect 8392 9890 14696 9922
rect 15110 9890 15470 13586
rect 8392 9886 15470 9890
rect 8312 9882 15470 9886
rect 800 9724 15470 9882
rect 800 9562 994 9724
rect 1146 9562 15470 9724
rect 800 9530 15470 9562
rect 800 9376 13253 9530
rect 6108 6638 6646 6736
rect 6108 6580 6226 6638
rect 6282 6580 6646 6638
rect 6108 6556 6646 6580
rect 372 6088 6274 6108
rect 372 6074 6170 6088
rect 372 5986 392 6074
rect 498 6030 6170 6074
rect 6226 6030 6274 6088
rect 498 5986 6274 6030
rect 372 5954 6274 5986
rect 6466 5814 6646 6556
rect 9652 6050 18838 6222
rect 9652 6042 11818 6050
rect 9652 5814 9832 6042
rect 802 5774 9844 5814
rect 802 5670 936 5774
rect 1052 5670 9844 5774
rect 802 5634 9844 5670
rect 2512 5578 2692 5634
rect 4378 5620 4558 5634
rect 2512 5520 2564 5578
rect 2620 5520 2692 5578
rect 2512 5506 2692 5520
rect 4628 5574 4808 5634
rect 6104 5620 6284 5634
rect 6572 5602 6766 5634
rect 8010 5620 8190 5634
rect 6572 5574 6762 5602
rect 4628 5570 4810 5574
rect 4628 5512 4686 5570
rect 4742 5512 4810 5570
rect 4628 5492 4810 5512
rect 6570 5570 6762 5574
rect 6570 5512 6638 5570
rect 6694 5512 6762 5570
rect 6570 5492 6762 5512
rect 8584 5576 8762 5634
rect 8584 5518 8640 5576
rect 8696 5574 8762 5576
rect 8696 5518 8764 5574
rect 8584 5498 8764 5518
rect 4628 5478 4808 5492
rect 6570 5488 6750 5492
rect 10128 5120 10308 6042
rect 10708 6000 10888 6042
rect 10708 5936 10774 6000
rect 10832 5936 10888 6000
rect 10708 5924 10888 5936
rect 12736 5986 12922 6050
rect 12736 5928 12796 5986
rect 12852 5928 12922 5986
rect 12736 5922 12922 5928
rect 12740 5908 12920 5922
rect 10972 5452 12936 5480
rect 10972 5394 11214 5452
rect 11270 5440 12936 5452
rect 11270 5394 12800 5440
rect 10972 5382 12800 5394
rect 12856 5382 12936 5440
rect 10972 5300 12936 5382
rect 10128 5062 10188 5120
rect 10244 5062 10308 5120
rect 2520 5040 2700 5048
rect 2520 4982 2584 5040
rect 2640 4982 2700 5040
rect 2520 4850 2700 4982
rect 4628 5024 4808 5048
rect 4628 4966 4690 5024
rect 4746 4966 4808 5024
rect 4380 4850 4560 4858
rect 4628 4850 4808 4966
rect 6580 5024 6760 5048
rect 6580 4966 6642 5024
rect 6698 4966 6760 5024
rect 6580 4948 6760 4966
rect 6092 4850 6272 4858
rect 6574 4850 6760 4948
rect 8582 5030 8762 5054
rect 10128 5046 10308 5062
rect 8582 4972 8644 5030
rect 8700 4972 8762 5030
rect 8002 4852 8182 4858
rect 8582 4852 8762 4972
rect 7674 4850 9835 4852
rect 198 4814 9835 4850
rect 198 4710 330 4814
rect 446 4710 9835 4814
rect 198 4670 9835 4710
rect 9652 4496 9832 4670
rect 10732 4580 10912 4598
rect 10732 4522 10788 4580
rect 10844 4522 10912 4580
rect 9652 4376 9834 4496
rect 10732 4376 10912 4522
rect 11576 4376 11756 5300
rect 13626 5174 13798 6050
rect 14696 5994 14882 6050
rect 14696 5952 14754 5994
rect 14698 5936 14754 5952
rect 14810 5952 14882 5994
rect 16690 6000 16876 6050
rect 17510 6042 18838 6050
rect 16690 5958 16748 6000
rect 14810 5936 14878 5952
rect 14698 5916 14878 5936
rect 16692 5942 16748 5958
rect 16804 5958 16876 6000
rect 16804 5942 16872 5958
rect 16692 5922 16872 5942
rect 14688 5454 16890 5480
rect 14688 5448 16752 5454
rect 14688 5390 14758 5448
rect 14814 5396 16752 5448
rect 16808 5396 16890 5454
rect 14814 5390 16890 5396
rect 14688 5308 16890 5390
rect 12976 5124 15154 5174
rect 12976 5080 15156 5124
rect 12976 5022 13032 5080
rect 13088 5074 15156 5080
rect 13088 5022 15034 5074
rect 12976 5016 15034 5022
rect 15090 5072 15156 5074
rect 15090 5016 15158 5072
rect 12976 5002 15158 5016
rect 14978 4996 15158 5002
rect 12974 4534 13154 4558
rect 12974 4476 13036 4534
rect 13092 4476 13154 4534
rect 9652 4368 11818 4376
rect 12974 4368 13154 4476
rect 14976 4528 15156 4552
rect 14976 4470 15038 4528
rect 15094 4470 15156 4528
rect 14976 4368 15156 4470
rect 15878 4368 16050 5308
rect 17648 5168 17828 6042
rect 18658 5428 18838 6042
rect 18658 5364 18726 5428
rect 18784 5364 18838 5428
rect 18658 5354 18838 5364
rect 17002 5106 17828 5168
rect 17000 5056 17828 5106
rect 17000 4998 17056 5056
rect 17112 4998 17828 5056
rect 17000 4988 17828 4998
rect 17000 4978 17180 4988
rect 18662 4880 18842 4888
rect 18662 4816 18720 4880
rect 18778 4816 18842 4880
rect 9652 4352 16050 4368
rect 16998 4510 17178 4534
rect 16998 4452 17060 4510
rect 17116 4452 17178 4510
rect 16998 4368 17178 4452
rect 18662 4376 18842 4816
rect 17510 4368 18840 4376
rect 16998 4352 18840 4368
rect 9652 4328 18840 4352
rect 9656 4196 18840 4328
rect 6082 3382 6656 3408
rect 6082 3320 6194 3382
rect 6254 3320 6656 3382
rect 6082 3228 6656 3320
rect 294 2828 6298 2858
rect 294 2808 6176 2828
rect 294 2714 384 2808
rect 484 2766 6176 2808
rect 6236 2766 6298 2828
rect 484 2714 6298 2766
rect 294 2664 6298 2714
rect 6476 2554 6656 3228
rect 794 2518 16633 2554
rect 794 2410 936 2518
rect 1068 2410 16633 2518
rect 794 2380 16633 2410
rect 794 2374 3426 2380
rect 3626 2374 5476 2380
rect 5676 2376 16633 2380
rect 2540 2318 2720 2374
rect 2540 2260 2604 2318
rect 2660 2260 2720 2318
rect 2540 2244 2720 2260
rect 4536 2314 4716 2374
rect 4536 2256 4592 2314
rect 4648 2256 4716 2314
rect 4536 2236 4716 2256
rect 6476 2314 6668 2376
rect 6476 2256 6544 2314
rect 6600 2256 6668 2314
rect 6476 2236 6668 2256
rect 8490 2320 8670 2376
rect 8490 2262 8546 2320
rect 8602 2262 8670 2320
rect 8490 2242 8670 2262
rect 10430 2320 10622 2376
rect 10430 2262 10498 2320
rect 10554 2262 10622 2320
rect 10430 2242 10622 2262
rect 12434 2320 12614 2376
rect 12434 2262 12490 2320
rect 12546 2262 12614 2320
rect 12434 2242 12614 2262
rect 14374 2320 14566 2376
rect 14374 2262 14442 2320
rect 14498 2262 14566 2320
rect 14374 2242 14566 2262
rect 16438 2320 16630 2376
rect 16438 2262 16506 2320
rect 16562 2262 16630 2320
rect 16438 2242 16630 2262
rect 10430 2238 10610 2242
rect 14374 2238 14554 2242
rect 16438 2238 16618 2242
rect 6476 2232 6656 2236
rect 2542 1778 2722 1790
rect 2542 1720 2604 1778
rect 2660 1720 2722 1778
rect 2542 1590 2722 1720
rect 4534 1768 4714 1792
rect 4534 1710 4596 1768
rect 4652 1710 4714 1768
rect 4534 1590 4714 1710
rect 6486 1768 6666 1792
rect 6486 1710 6548 1768
rect 6604 1710 6666 1768
rect 6486 1692 6666 1710
rect 6480 1590 6666 1692
rect 8488 1774 8668 1798
rect 8488 1716 8550 1774
rect 8606 1716 8668 1774
rect 8488 1596 8668 1716
rect 10440 1774 10620 1798
rect 10440 1716 10502 1774
rect 10558 1716 10620 1774
rect 10440 1698 10620 1716
rect 10434 1596 10620 1698
rect 12432 1774 12612 1798
rect 12432 1716 12494 1774
rect 12550 1716 12612 1774
rect 12432 1596 12612 1716
rect 14384 1774 14564 1798
rect 14384 1716 14446 1774
rect 14502 1716 14564 1774
rect 16448 1774 16628 1798
rect 16448 1716 16510 1774
rect 16566 1716 16628 1774
rect 14384 1698 14564 1716
rect 14378 1596 14564 1698
rect 16442 1686 16628 1716
rect 16442 1656 16626 1686
rect 7580 1592 9430 1596
rect 9630 1592 11402 1596
rect 11524 1592 13374 1596
rect 13574 1592 15346 1596
rect 7456 1590 15346 1592
rect 210 1586 3426 1590
rect 3626 1586 5476 1590
rect 5676 1588 15630 1590
rect 16446 1588 16626 1656
rect 5676 1586 16626 1588
rect 210 1548 16626 1586
rect 210 1438 336 1548
rect 456 1438 16626 1548
rect 210 1410 16626 1438
<< via3 >>
rect 18768 43898 18962 44096
rect 300 24092 488 24272
rect 978 21970 1166 22150
rect 996 17780 1066 17848
rect 322 16942 474 17104
rect 27000 14646 27122 14766
rect 27550 14372 27682 14492
rect 994 9562 1146 9724
rect 392 5986 498 6074
rect 936 5670 1052 5774
rect 330 4710 446 4814
rect 384 2714 484 2808
rect 936 2410 1068 2518
rect 336 1438 456 1548
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 44952 12818 45152
rect 13310 44952 13370 45152
rect 13862 44952 13922 45152
rect 14414 44952 14474 45152
rect 14966 44952 15026 45152
rect 15518 44952 15578 45152
rect 16070 44952 16130 45152
rect 16622 44952 16682 45152
rect 17174 44952 17234 45152
rect 17726 44952 17786 45152
rect 18278 44952 18338 45152
rect 18830 44168 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 200 24272 600 44152
rect 200 24092 300 24272
rect 488 24092 600 24272
rect 200 17104 600 24092
rect 200 16942 322 17104
rect 474 16942 600 17104
rect 200 6074 600 16942
rect 200 5986 392 6074
rect 498 5986 600 6074
rect 200 4814 600 5986
rect 200 4710 330 4814
rect 446 4710 600 4814
rect 200 2808 600 4710
rect 200 2714 384 2808
rect 484 2714 600 2808
rect 200 1548 600 2714
rect 200 1438 336 1548
rect 456 1438 600 1548
rect 200 1000 600 1438
rect 800 22150 1200 44152
rect 18590 44096 19130 44168
rect 18590 43898 18768 44096
rect 18962 43898 19130 44096
rect 18590 43830 19130 43898
rect 800 21970 978 22150
rect 1166 21970 1200 22150
rect 800 17848 1200 21970
rect 800 17780 996 17848
rect 1066 17780 1200 17848
rect 800 9724 1200 17780
rect 27110 14788 27170 45152
rect 26956 14766 27174 14788
rect 26956 14646 27000 14766
rect 27122 14646 27174 14766
rect 26956 14604 27174 14646
rect 27662 14510 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 27512 14492 27730 14510
rect 27512 14372 27550 14492
rect 27682 14372 27730 14492
rect 27512 14336 27730 14372
rect 800 9562 994 9724
rect 1146 9562 1200 9724
rect 800 5774 1200 9562
rect 800 5670 936 5774
rect 1052 5670 1200 5774
rect 800 2518 1200 5670
rect 800 2410 936 2518
rect 1068 2410 1200 2518
rect 800 1000 1200 2410
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
rlabel metal1 s 9916 23328 11664 23424 1 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 9916 22784 11664 22880 1 VGND
port 3 nsew ground bidirectional abutment
rlabel comment s 9916 22832 9916 22832 4 dfxbp_1
flabel nwell s 9962 23376 9962 23376 0 FreeSans 200 0 0 0 VPB
flabel nwell s 9945 23359 9979 23393 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 9962 22832 9962 22832 0 FreeSans 200 0 0 0 VNB
flabel pwell s 9945 22815 9979 22849 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel locali s 11306 22917 11340 22951 0 FreeSans 400 0 0 0 Q
port 7 nsew signal output
flabel locali s 9945 23053 9979 23087 0 FreeSans 400 0 0 0 CLK
port 1 nsew clock input
flabel locali s 10205 23053 10239 23087 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 11601 23136 11635 23170 0 FreeSans 400 0 0 0 Q_N
port 8 nsew signal output
flabel metal1 s 9945 23359 9979 23393 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 9945 22815 9979 22849 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 11664 23328 11756 23424 1 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 11664 22784 11756 22880 1 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 11664 22832 11664 22832 4 tapvpwrvgnd_1
flabel metal1 s 11685 22814 11736 22852 0 FreeSans 200 0 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 11686 23356 11739 23385 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 16096 23324 16188 23420 1 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 16096 22780 16188 22876 1 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 16096 22828 16096 22828 4 tapvpwrvgnd_1
flabel metal1 s 16117 22810 16168 22848 0 FreeSans 200 0 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 16118 23352 16171 23381 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 14348 23324 16096 23420 1 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 14348 22780 16096 22876 1 VGND
port 3 nsew ground bidirectional abutment
rlabel comment s 14348 22828 14348 22828 4 dfxbp_1
flabel nwell s 14394 23372 14394 23372 0 FreeSans 200 0 0 0 VPB
flabel nwell s 14377 23355 14411 23389 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 14394 22828 14394 22828 0 FreeSans 200 0 0 0 VNB
flabel pwell s 14377 22811 14411 22845 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel locali s 15738 22913 15772 22947 0 FreeSans 400 0 0 0 Q
port 7 nsew signal output
flabel locali s 14377 23049 14411 23083 0 FreeSans 400 0 0 0 CLK
port 1 nsew clock input
flabel locali s 14637 23049 14671 23083 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 16033 23132 16067 23166 0 FreeSans 400 0 0 0 Q_N
port 8 nsew signal output
flabel metal1 s 14377 23355 14411 23389 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 14377 22811 14411 22845 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 12102 23320 13850 23416 1 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 12102 22776 13850 22872 1 VGND
port 3 nsew ground bidirectional abutment
rlabel comment s 12102 22824 12102 22824 4 dfxbp_1
flabel nwell s 12148 23368 12148 23368 0 FreeSans 200 0 0 0 VPB
flabel nwell s 12131 23351 12165 23385 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 12148 22824 12148 22824 0 FreeSans 200 0 0 0 VNB
flabel pwell s 12131 22807 12165 22841 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel locali s 13492 22909 13526 22943 0 FreeSans 400 0 0 0 Q
port 7 nsew signal output
flabel locali s 12131 23045 12165 23079 0 FreeSans 400 0 0 0 CLK
port 1 nsew clock input
flabel locali s 12391 23045 12425 23079 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 13787 23128 13821 23162 0 FreeSans 400 0 0 0 Q_N
port 8 nsew signal output
flabel metal1 s 12131 23351 12165 23385 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 12131 22807 12165 22841 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 13850 23320 13942 23416 1 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 13850 22776 13942 22872 1 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 13850 22824 13850 22824 4 tapvpwrvgnd_1
flabel metal1 s 13871 22806 13922 22844 0 FreeSans 200 0 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 13872 23348 13925 23377 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 18400 23352 18453 23381 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 18399 22810 18450 22848 0 FreeSans 200 0 0 0 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 18378 22828 18378 22828 4 tapvpwrvgnd_1
rlabel metal1 s 18378 22780 18470 22876 1 VGND
port 1 nsew ground bidirectional abutment
rlabel metal1 s 18378 23324 18470 23420 1 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 16659 22811 16693 22845 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 16659 23355 16693 23389 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel locali s 18315 23132 18349 23166 0 FreeSans 400 0 0 0 Q_N
port 8 nsew signal output
flabel locali s 16919 23049 16953 23083 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 16659 23049 16693 23083 0 FreeSans 400 0 0 0 CLK
port 1 nsew clock input
flabel locali s 18020 22913 18054 22947 0 FreeSans 400 0 0 0 Q
port 7 nsew signal output
flabel pwell s 16659 22811 16693 22845 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel pwell s 16676 22828 16676 22828 0 FreeSans 200 0 0 0 VNB
flabel nwell s 16659 23355 16693 23389 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel nwell s 16676 23372 16676 23372 0 FreeSans 200 0 0 0 VPB
rlabel comment s 16630 22828 16630 22828 4 dfxbp_1
rlabel metal1 s 16630 22780 18378 22876 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 16630 23324 18378 23420 1 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 9440 23352 9493 23381 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_73.VPWR
flabel metal1 9439 22810 9490 22848 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_73.VGND
rlabel comment 9418 22828 9418 22828 4 sky130_fd_sc_hd__tapvpwrvgnd_1_73.tapvpwrvgnd_1
rlabel metal1 9418 22780 9510 22876 1 sky130_fd_sc_hd__tapvpwrvgnd_1_73.VGND
rlabel metal1 9418 23324 9510 23420 1 sky130_fd_sc_hd__tapvpwrvgnd_1_73.VPWR
flabel metal1 7699 22811 7733 22845 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0.VGND
flabel metal1 7699 23355 7733 23389 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0.VPWR
flabel locali 9355 23132 9389 23166 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_0.Q_N
flabel locali 7959 23049 7993 23083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0.D
flabel locali 7699 23049 7733 23083 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_0.CLK
flabel locali 9060 22913 9094 22947 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_0.Q
flabel pwell 7699 22811 7733 22845 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0.VNB
flabel pwell 7716 22828 7716 22828 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0.VNB
flabel nwell 7699 23355 7733 23389 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0.VPB
flabel nwell 7716 23372 7716 23372 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_0.VPB
rlabel comment 7670 22828 7670 22828 4 sky130_fd_sc_hd__dfxbp_1_0.dfxbp_1
rlabel metal1 7670 22780 9418 22876 1 sky130_fd_sc_hd__dfxbp_1_0.VGND
rlabel metal1 7670 23324 9418 23420 1 sky130_fd_sc_hd__dfxbp_1_0.VPWR
flabel metal1 12131 22807 12165 22841 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_2.VGND
flabel metal1 12131 23351 12165 23385 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_2.VPWR
flabel locali 13787 23128 13821 23162 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_2.Q_N
flabel locali 12391 23045 12425 23079 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_2.D
flabel locali 12131 23045 12165 23079 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_2.CLK
flabel locali 13492 22909 13526 22943 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_2.Q
flabel pwell 12131 22807 12165 22841 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_2.VNB
flabel pwell 12148 22824 12148 22824 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_2.VNB
flabel nwell 12131 23351 12165 23385 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_2.VPB
flabel nwell 12148 23368 12148 23368 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_2.VPB
rlabel comment 12102 22824 12102 22824 4 sky130_fd_sc_hd__dfxbp_1_2.dfxbp_1
rlabel metal1 12102 22776 13850 22872 1 sky130_fd_sc_hd__dfxbp_1_2.VGND
rlabel metal1 12102 23320 13850 23416 1 sky130_fd_sc_hd__dfxbp_1_2.VPWR
flabel metal1 9945 22815 9979 22849 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1.VGND
flabel metal1 9945 23359 9979 23393 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1.VPWR
flabel locali 11601 23136 11635 23170 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_1.Q_N
flabel locali 10205 23053 10239 23087 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1.D
flabel locali 9945 23053 9979 23087 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_1.CLK
flabel locali 11306 22917 11340 22951 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_1.Q
flabel pwell 9945 22815 9979 22849 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1.VNB
flabel pwell 9962 22832 9962 22832 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1.VNB
flabel nwell 9945 23359 9979 23393 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1.VPB
flabel nwell 9962 23376 9962 23376 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_1.VPB
rlabel comment 9916 22832 9916 22832 4 sky130_fd_sc_hd__dfxbp_1_1.dfxbp_1
rlabel metal1 9916 22784 11664 22880 1 sky130_fd_sc_hd__dfxbp_1_1.VGND
rlabel metal1 9916 23328 11664 23424 1 sky130_fd_sc_hd__dfxbp_1_1.VPWR
flabel metal1 11686 23356 11739 23385 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_74.VPWR
flabel metal1 11685 22814 11736 22852 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_74.VGND
rlabel comment 11664 22832 11664 22832 4 sky130_fd_sc_hd__tapvpwrvgnd_1_74.tapvpwrvgnd_1
rlabel metal1 11664 22784 11756 22880 1 sky130_fd_sc_hd__tapvpwrvgnd_1_74.VGND
rlabel metal1 11664 23328 11756 23424 1 sky130_fd_sc_hd__tapvpwrvgnd_1_74.VPWR
flabel metal1 16659 22811 16693 22845 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_4.VGND
flabel metal1 16659 23355 16693 23389 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_4.VPWR
flabel locali 18315 23132 18349 23166 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_4.Q_N
flabel locali 16919 23049 16953 23083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_4.D
flabel locali 16659 23049 16693 23083 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_4.CLK
flabel locali 18020 22913 18054 22947 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_4.Q
flabel pwell 16659 22811 16693 22845 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_4.VNB
flabel pwell 16676 22828 16676 22828 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_4.VNB
flabel nwell 16659 23355 16693 23389 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_4.VPB
flabel nwell 16676 23372 16676 23372 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_4.VPB
rlabel comment 16630 22828 16630 22828 4 sky130_fd_sc_hd__dfxbp_1_4.dfxbp_1
rlabel metal1 16630 22780 18378 22876 1 sky130_fd_sc_hd__dfxbp_1_4.VGND
rlabel metal1 16630 23324 18378 23420 1 sky130_fd_sc_hd__dfxbp_1_4.VPWR
flabel metal1 16118 23352 16171 23381 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_76.VPWR
flabel metal1 16117 22810 16168 22848 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_76.VGND
rlabel comment 16096 22828 16096 22828 4 sky130_fd_sc_hd__tapvpwrvgnd_1_76.tapvpwrvgnd_1
rlabel metal1 16096 22780 16188 22876 1 sky130_fd_sc_hd__tapvpwrvgnd_1_76.VGND
rlabel metal1 16096 23324 16188 23420 1 sky130_fd_sc_hd__tapvpwrvgnd_1_76.VPWR
flabel metal1 14377 22811 14411 22845 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_3.VGND
flabel metal1 14377 23355 14411 23389 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_3.VPWR
flabel locali 16033 23132 16067 23166 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_3.Q_N
flabel locali 14637 23049 14671 23083 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_3.D
flabel locali 14377 23049 14411 23083 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_3.CLK
flabel locali 15738 22913 15772 22947 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_3.Q
flabel pwell 14377 22811 14411 22845 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_3.VNB
flabel pwell 14394 22828 14394 22828 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_3.VNB
flabel nwell 14377 23355 14411 23389 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_3.VPB
flabel nwell 14394 23372 14394 23372 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_3.VPB
rlabel comment 14348 22828 14348 22828 4 sky130_fd_sc_hd__dfxbp_1_3.dfxbp_1
rlabel metal1 14348 22780 16096 22876 1 sky130_fd_sc_hd__dfxbp_1_3.VGND
rlabel metal1 14348 23324 16096 23420 1 sky130_fd_sc_hd__dfxbp_1_3.VPWR
flabel metal1 13872 23348 13925 23377 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_75.VPWR
flabel metal1 13871 22806 13922 22844 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_75.VGND
rlabel comment 13850 22824 13850 22824 4 sky130_fd_sc_hd__tapvpwrvgnd_1_75.tapvpwrvgnd_1
rlabel metal1 13850 22776 13942 22872 1 sky130_fd_sc_hd__tapvpwrvgnd_1_75.VGND
rlabel metal1 13850 23320 13942 23416 1 sky130_fd_sc_hd__tapvpwrvgnd_1_75.VPWR
flabel metal1 18400 23352 18453 23381 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_77.VPWR
flabel metal1 18399 22810 18450 22848 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_77.VGND
rlabel comment 18378 22828 18378 22828 4 sky130_fd_sc_hd__tapvpwrvgnd_1_77.tapvpwrvgnd_1
rlabel metal1 18378 22780 18470 22876 1 sky130_fd_sc_hd__tapvpwrvgnd_1_77.VGND
rlabel metal1 18378 23324 18470 23420 1 sky130_fd_sc_hd__tapvpwrvgnd_1_77.VPWR
rlabel metal1 18548 43418 18644 43510 7 sky130_fd_sc_hd__tapvpwrvgnd_1_89.VPWR
rlabel metal1 19092 43418 19188 43510 7 sky130_fd_sc_hd__tapvpwrvgnd_1_89.VGND
rlabel comment 19140 43418 19140 43418 2 sky130_fd_sc_hd__tapvpwrvgnd_1_89.tapvpwrvgnd_1
flabel metal1 19120 43439 19158 43490 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_89.VGND
flabel metal1 18587 43440 18616 43493 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_89.VPWR
rlabel metal1 18532 41432 18628 41524 7 sky130_fd_sc_hd__tapvpwrvgnd_1_88.VPWR
rlabel metal1 19076 41432 19172 41524 7 sky130_fd_sc_hd__tapvpwrvgnd_1_88.VGND
rlabel comment 19124 41432 19124 41432 2 sky130_fd_sc_hd__tapvpwrvgnd_1_88.tapvpwrvgnd_1
flabel metal1 19104 41453 19142 41504 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_88.VGND
flabel metal1 18571 41454 18600 41507 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_88.VPWR
rlabel metal1 18540 39636 18636 39728 7 sky130_fd_sc_hd__tapvpwrvgnd_1_87.VPWR
rlabel metal1 19084 39636 19180 39728 7 sky130_fd_sc_hd__tapvpwrvgnd_1_87.VGND
rlabel comment 19132 39636 19132 39636 2 sky130_fd_sc_hd__tapvpwrvgnd_1_87.tapvpwrvgnd_1
flabel metal1 19112 39657 19150 39708 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_87.VGND
flabel metal1 18579 39658 18608 39711 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_87.VPWR
rlabel metal1 18548 41948 18644 43420 7 sky130_fd_sc_hd__inv_16_0.VPWR
rlabel metal1 19092 41948 19188 43420 7 sky130_fd_sc_hd__inv_16_0.VGND
rlabel comment 19140 41948 19140 41948 2 sky130_fd_sc_hd__inv_16_0.inv_16
flabel metal1 18579 41977 18613 42011 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_16_0.VPWR
flabel metal1 19123 41977 19157 42011 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_16_0.VGND
flabel pwell 19123 41977 19157 42011 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_16_0.VNB
flabel nwell 18579 41977 18613 42011 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_16_0.VPB
flabel locali 18885 42805 18919 42839 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_16_0.A
flabel locali 18885 42713 18919 42747 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_16_0.A
flabel locali 18885 42345 18919 42379 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_16_0.A
flabel locali 18885 41977 18919 42011 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_16_0.A
flabel locali 18953 43265 18987 43299 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_16_0.Y
flabel locali 18885 43265 18919 43299 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_16_0.Y
rlabel metal1 18532 40236 18628 41432 7 sky130_fd_sc_hd__inv_12_0.VPWR
rlabel metal1 19076 40236 19172 41432 7 sky130_fd_sc_hd__inv_12_0.VGND
rlabel comment 19124 40236 19124 40236 2 sky130_fd_sc_hd__inv_12_0.inv_12
flabel metal1 18563 40265 18597 40299 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_12_0.VPWR
flabel metal1 19107 40265 19141 40299 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_12_0.VGND
flabel nwell 18563 40265 18597 40299 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_12_0.VPB
flabel pwell 19107 40265 19141 40299 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_12_0.VNB
flabel locali 18869 41237 18903 41271 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_12_0.A
flabel locali 18869 41153 18903 41187 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_12_0.A
flabel locali 18869 41077 18903 41111 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_12_0.A
flabel locali 18869 40985 18903 41019 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_12_0.A
flabel locali 18869 40265 18903 40299 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_12_0.Y
flabel locali 18869 41369 18903 41403 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_12_0.Y
flabel locali 18869 40909 18903 40943 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_12_0.A
flabel locali 18869 40817 18903 40851 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_12_0.A
flabel locali 18869 40725 18903 40759 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_12_0.A
flabel locali 18869 40633 18903 40667 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_12_0.A
flabel locali 18869 40541 18903 40575 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_12_0.A
flabel locali 18869 40449 18903 40483 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_12_0.A
rlabel metal1 18540 38808 18636 39636 7 sky130_fd_sc_hd__inv_8_0.VPWR
rlabel metal1 19084 38808 19180 39636 7 sky130_fd_sc_hd__inv_8_0.VGND
rlabel comment 19132 38808 19132 38808 2 sky130_fd_sc_hd__inv_8_0.inv_8
flabel metal1 18571 38837 18605 38871 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_8_0.VPWR
flabel metal1 19115 38837 19149 38871 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_8_0.VGND
flabel nwell 18571 38837 18605 38871 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_8_0.VPB
flabel pwell 19115 38837 19149 38871 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_8_0.VNB
flabel locali 18877 38837 18911 38871 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_8_0.Y
flabel locali 18877 39573 18911 39607 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_8_0.Y
flabel locali 18877 39481 18911 39515 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_8_0.A
flabel locali 18877 39389 18911 39423 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_8_0.A
flabel locali 18877 39297 18911 39331 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_8_0.A
flabel locali 18877 39205 18911 39239 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_8_0.A
flabel locali 18877 39113 18911 39147 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_8_0.A
flabel locali 18877 39021 18911 39055 0 FreeSans 250 0 0 0 sky130_fd_sc_hd__inv_8_0.A
rlabel metal1 18554 38374 18650 38466 7 sky130_fd_sc_hd__tapvpwrvgnd_1_86.VPWR
rlabel metal1 19098 38374 19194 38466 7 sky130_fd_sc_hd__tapvpwrvgnd_1_86.VGND
rlabel comment 19146 38374 19146 38374 2 sky130_fd_sc_hd__tapvpwrvgnd_1_86.tapvpwrvgnd_1
flabel metal1 19126 38395 19164 38446 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_86.VGND
flabel metal1 18593 38396 18622 38449 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_86.VPWR
rlabel metal1 18566 36764 18662 37224 7 sky130_fd_sc_hd__inv_4_0.VPWR
rlabel metal1 19110 36764 19206 37224 7 sky130_fd_sc_hd__inv_4_0.VGND
rlabel comment 19158 36764 19158 36764 2 sky130_fd_sc_hd__inv_4_0.inv_4
flabel metal1 19141 36793 19175 36827 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_0.VGND
flabel metal1 18597 36793 18631 36827 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_0.VPWR
flabel pwell 19141 36793 19175 36827 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_0.VNB
flabel nwell 18597 36793 18631 36827 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_4_0.VPB
flabel locali 18903 37069 18937 37103 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0.A
flabel locali 18903 36977 18937 37011 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0.A
flabel locali 18903 36885 18937 36919 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0.A
flabel locali 18903 36793 18937 36827 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0.A
flabel locali 18835 37161 18869 37195 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0.Y
flabel locali 18903 37161 18937 37195 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0.Y
flabel locali 18971 37161 19005 37195 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_4_0.Y
rlabel metal1 18554 37730 18650 38374 7 sky130_fd_sc_hd__inv_6_0.VPWR
rlabel metal1 19098 37730 19194 38374 7 sky130_fd_sc_hd__inv_6_0.VGND
rlabel comment 19146 37730 19146 37730 2 sky130_fd_sc_hd__inv_6_0.inv_6
flabel metal1 19129 37759 19163 37793 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_6_0.VGND
flabel metal1 18585 37759 18619 37793 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_6_0.VPWR
flabel pwell 19129 37759 19163 37793 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_6_0.VNB
flabel nwell 18585 37759 18619 37793 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_6_0.VPB
flabel locali 18891 38211 18925 38245 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_6_0.A
flabel locali 18891 38119 18925 38153 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_6_0.A
flabel locali 18891 38027 18925 38061 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_6_0.A
flabel locali 18891 37759 18925 37793 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_6_0.A
flabel locali 18823 38303 18857 38337 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_6_0.Y
flabel locali 18891 38303 18925 38337 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_6_0.Y
flabel locali 18959 38303 18993 38337 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_6_0.Y
rlabel metal1 18574 36336 18670 36428 7 sky130_fd_sc_hd__tapvpwrvgnd_1_84.VPWR
rlabel metal1 19118 36336 19214 36428 7 sky130_fd_sc_hd__tapvpwrvgnd_1_84.VGND
rlabel comment 19166 36336 19166 36336 2 sky130_fd_sc_hd__tapvpwrvgnd_1_84.tapvpwrvgnd_1
flabel metal1 19146 36357 19184 36408 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_84.VGND
flabel metal1 18613 36358 18642 36411 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_84.VPWR
rlabel metal1 18566 37220 18662 37312 7 sky130_fd_sc_hd__tapvpwrvgnd_1_85.VPWR
rlabel metal1 19110 37220 19206 37312 7 sky130_fd_sc_hd__tapvpwrvgnd_1_85.VGND
rlabel comment 19158 37220 19158 37220 2 sky130_fd_sc_hd__tapvpwrvgnd_1_85.tapvpwrvgnd_1
flabel metal1 19138 37241 19176 37292 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_85.VGND
flabel metal1 18605 37242 18634 37295 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_85.VPWR
rlabel metal1 18574 36060 18670 36336 7 sky130_fd_sc_hd__inv_2_0.VPWR
rlabel metal1 19118 36060 19214 36336 7 sky130_fd_sc_hd__inv_2_0.VGND
rlabel comment 19166 36060 19166 36060 2 sky130_fd_sc_hd__inv_2_0.inv_2
flabel metal1 19149 36089 19183 36123 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_2_0.VGND
flabel metal1 18605 36089 18639 36123 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_2_0.VPWR
flabel pwell 19149 36089 19183 36123 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_2_0.VNB
flabel nwell 18605 36089 18639 36123 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__inv_2_0.VPB
flabel locali 18911 36181 18945 36215 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_2_0.Y
flabel locali 18843 36181 18877 36215 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_2_0.Y
flabel locali 18979 36181 19013 36215 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_2_0.Y
flabel locali 18911 36089 18945 36123 0 FreeSans 340 0 0 0 sky130_fd_sc_hd__inv_2_0.A
rlabel metal1 18598 34948 18694 35040 7 sky130_fd_sc_hd__tapvpwrvgnd_1_82.VPWR
rlabel metal1 19142 34948 19238 35040 7 sky130_fd_sc_hd__tapvpwrvgnd_1_82.VGND
rlabel comment 19190 34948 19190 34948 2 sky130_fd_sc_hd__tapvpwrvgnd_1_82.tapvpwrvgnd_1
flabel metal1 19170 34969 19208 35020 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_82.VGND
flabel metal1 18637 34970 18666 35023 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_82.VPWR
rlabel metal1 18598 32666 18694 32758 7 sky130_fd_sc_hd__tapvpwrvgnd_1_80.VPWR
rlabel metal1 19142 32666 19238 32758 7 sky130_fd_sc_hd__tapvpwrvgnd_1_80.VGND
rlabel comment 19190 32666 19190 32666 2 sky130_fd_sc_hd__tapvpwrvgnd_1_80.tapvpwrvgnd_1
flabel metal1 19170 32687 19208 32738 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_80.VGND
flabel metal1 18637 32688 18666 32741 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_80.VPWR
rlabel metal1 18598 33200 18694 34948 7 sky130_fd_sc_hd__dfxbp_1_8.VPWR
rlabel metal1 19142 33200 19238 34948 7 sky130_fd_sc_hd__dfxbp_1_8.VGND
rlabel comment 19190 33200 19190 33200 2 sky130_fd_sc_hd__dfxbp_1_8.dfxbp_1
flabel nwell 18646 33246 18646 33246 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_8.VPB
flabel nwell 18629 33229 18663 33263 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_8.VPB
flabel pwell 19190 33246 19190 33246 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_8.VNB
flabel pwell 19173 33229 19207 33263 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_8.VNB
flabel locali 19071 34590 19105 34624 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_8.Q
flabel locali 18935 33229 18969 33263 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_8.CLK
flabel locali 18935 33489 18969 33523 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_8.D
flabel locali 18852 34885 18886 34919 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_8.Q_N
flabel metal1 18629 33229 18663 33263 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_8.VPWR
flabel metal1 19173 33229 19207 33263 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_8.VGND
rlabel metal1 18602 30420 18698 30512 7 sky130_fd_sc_hd__tapvpwrvgnd_1_81.VPWR
rlabel metal1 19146 30420 19242 30512 7 sky130_fd_sc_hd__tapvpwrvgnd_1_81.VGND
rlabel comment 19194 30420 19194 30420 2 sky130_fd_sc_hd__tapvpwrvgnd_1_81.tapvpwrvgnd_1
flabel metal1 19174 30441 19212 30492 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_81.VGND
flabel metal1 18641 30442 18670 30495 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_81.VPWR
rlabel metal1 18598 30918 18694 32666 7 sky130_fd_sc_hd__dfxbp_1_9.VPWR
rlabel metal1 19142 30918 19238 32666 7 sky130_fd_sc_hd__dfxbp_1_9.VGND
rlabel comment 19190 30918 19190 30918 2 sky130_fd_sc_hd__dfxbp_1_9.dfxbp_1
flabel nwell 18646 30964 18646 30964 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_9.VPB
flabel nwell 18629 30947 18663 30981 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_9.VPB
flabel pwell 19190 30964 19190 30964 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_9.VNB
flabel pwell 19173 30947 19207 30981 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_9.VNB
flabel locali 19071 32308 19105 32342 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_9.Q
flabel locali 18935 30947 18969 30981 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_9.CLK
flabel locali 18935 31207 18969 31241 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_9.D
flabel locali 18852 32603 18886 32637 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_9.Q_N
flabel metal1 18629 30947 18663 30981 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_9.VPWR
flabel metal1 19173 30947 19207 30981 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_9.VGND
rlabel metal1 18594 28234 18690 28326 7 sky130_fd_sc_hd__tapvpwrvgnd_1_79.VPWR
rlabel metal1 19138 28234 19234 28326 7 sky130_fd_sc_hd__tapvpwrvgnd_1_79.VGND
rlabel comment 19186 28234 19186 28234 2 sky130_fd_sc_hd__tapvpwrvgnd_1_79.tapvpwrvgnd_1
flabel metal1 19166 28255 19204 28306 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_79.VGND
flabel metal1 18633 28256 18662 28309 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_79.VPWR
rlabel metal1 18602 28672 18698 30420 7 sky130_fd_sc_hd__dfxbp_1_6.VPWR
rlabel metal1 19146 28672 19242 30420 7 sky130_fd_sc_hd__dfxbp_1_6.VGND
rlabel comment 19194 28672 19194 28672 2 sky130_fd_sc_hd__dfxbp_1_6.dfxbp_1
flabel nwell 18650 28718 18650 28718 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_6.VPB
flabel nwell 18633 28701 18667 28735 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_6.VPB
flabel pwell 19194 28718 19194 28718 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_6.VNB
flabel pwell 19177 28701 19211 28735 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_6.VNB
flabel locali 19075 30062 19109 30096 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_6.Q
flabel locali 18939 28701 18973 28735 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_6.CLK
flabel locali 18939 28961 18973 28995 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_6.D
flabel locali 18856 30357 18890 30391 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_6.Q_N
flabel metal1 18633 28701 18667 28735 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_6.VPWR
flabel metal1 19177 28701 19211 28735 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_6.VGND
rlabel metal1 18594 26486 18690 28234 7 sky130_fd_sc_hd__dfxbp_1_7.VPWR
rlabel metal1 19138 26486 19234 28234 7 sky130_fd_sc_hd__dfxbp_1_7.VGND
rlabel comment 19186 26486 19186 26486 2 sky130_fd_sc_hd__dfxbp_1_7.dfxbp_1
flabel nwell 18642 26532 18642 26532 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_7.VPB
flabel nwell 18625 26515 18659 26549 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_7.VPB
flabel pwell 19186 26532 19186 26532 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_7.VNB
flabel pwell 19169 26515 19203 26549 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_7.VNB
flabel locali 19067 27876 19101 27910 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_7.Q
flabel locali 18931 26515 18965 26549 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_7.CLK
flabel locali 18931 26775 18965 26809 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_7.D
flabel locali 18848 28171 18882 28205 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_7.Q_N
flabel metal1 18625 26515 18659 26549 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_7.VPWR
flabel metal1 19169 26515 19203 26549 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_7.VGND
rlabel metal1 18598 25988 18694 26080 7 sky130_fd_sc_hd__tapvpwrvgnd_1_78.VPWR
rlabel metal1 19142 25988 19238 26080 7 sky130_fd_sc_hd__tapvpwrvgnd_1_78.VGND
rlabel comment 19190 25988 19190 25988 2 sky130_fd_sc_hd__tapvpwrvgnd_1_78.tapvpwrvgnd_1
flabel metal1 19170 26009 19208 26060 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_78.VGND
flabel metal1 18637 26010 18666 26063 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__tapvpwrvgnd_1_78.VPWR
rlabel metal1 18598 24240 18694 25988 7 sky130_fd_sc_hd__dfxbp_1_5.VPWR
rlabel metal1 19142 24240 19238 25988 7 sky130_fd_sc_hd__dfxbp_1_5.VGND
rlabel comment 19190 24240 19190 24240 2 sky130_fd_sc_hd__dfxbp_1_5.dfxbp_1
flabel nwell 18646 24286 18646 24286 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_5.VPB
flabel nwell 18629 24269 18663 24303 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_5.VPB
flabel pwell 19190 24286 19190 24286 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_5.VNB
flabel pwell 19173 24269 19207 24303 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_5.VNB
flabel locali 19071 25630 19105 25664 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_5.Q
flabel locali 18935 24269 18969 24303 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_5.CLK
flabel locali 18935 24529 18969 24563 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_5.D
flabel locali 18852 25925 18886 25959 0 FreeSans 400 0 0 0 sky130_fd_sc_hd__dfxbp_1_5.Q_N
flabel metal1 18629 24269 18663 24303 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_5.VPWR
flabel metal1 19173 24269 19207 24303 0 FreeSans 200 0 0 0 sky130_fd_sc_hd__dfxbp_1_5.VGND
rlabel metal1 s 18598 34948 18694 35040 7 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 19142 34948 19238 35040 7 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 19190 34948 19190 34948 2 tapvpwrvgnd_1
flabel metal1 s 19170 34969 19208 35020 0 FreeSans 200 270 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 18637 34970 18666 35023 0 FreeSans 200 270 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 18602 30420 18698 30512 7 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 19146 30420 19242 30512 7 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 19194 30420 19194 30420 2 tapvpwrvgnd_1
flabel metal1 s 19174 30441 19212 30492 0 FreeSans 200 270 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 18641 30442 18670 30495 0 FreeSans 200 270 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 18598 30918 18694 32666 7 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 19142 30918 19238 32666 7 VGND
port 3 nsew ground bidirectional abutment
rlabel comment s 19190 30918 19190 30918 2 dfxbp_1
flabel nwell s 18646 30964 18646 30964 0 FreeSans 200 270 0 0 VPB
flabel nwell s 18629 30947 18663 30981 0 FreeSans 200 270 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 19190 30964 19190 30964 0 FreeSans 200 270 0 0 VNB
flabel pwell s 19173 30947 19207 30981 0 FreeSans 200 270 0 0 VNB
port 4 nsew ground bidirectional
flabel locali s 19071 32308 19105 32342 0 FreeSans 400 270 0 0 Q
port 7 nsew signal output
flabel locali s 18935 30947 18969 30981 0 FreeSans 400 270 0 0 CLK
port 1 nsew clock input
flabel locali s 18935 31207 18969 31241 0 FreeSans 200 270 0 0 D
port 2 nsew signal input
flabel locali s 18852 32603 18886 32637 0 FreeSans 400 270 0 0 Q_N
port 8 nsew signal output
flabel metal1 s 18629 30947 18663 30981 0 FreeSans 200 270 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 19173 30947 19207 30981 0 FreeSans 200 270 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 18598 32666 18694 32758 7 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 19142 32666 19238 32758 7 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 19190 32666 19190 32666 2 tapvpwrvgnd_1
flabel metal1 s 19170 32687 19208 32738 0 FreeSans 200 270 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 18637 32688 18666 32741 0 FreeSans 200 270 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 18598 33200 18694 34948 7 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 19142 33200 19238 34948 7 VGND
port 3 nsew ground bidirectional abutment
rlabel comment s 19190 33200 19190 33200 2 dfxbp_1
flabel nwell s 18646 33246 18646 33246 0 FreeSans 200 270 0 0 VPB
flabel nwell s 18629 33229 18663 33263 0 FreeSans 200 270 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 19190 33246 19190 33246 0 FreeSans 200 270 0 0 VNB
flabel pwell s 19173 33229 19207 33263 0 FreeSans 200 270 0 0 VNB
port 4 nsew ground bidirectional
flabel locali s 19071 34590 19105 34624 0 FreeSans 400 270 0 0 Q
port 7 nsew signal output
flabel locali s 18935 33229 18969 33263 0 FreeSans 400 270 0 0 CLK
port 1 nsew clock input
flabel locali s 18935 33489 18969 33523 0 FreeSans 200 270 0 0 D
port 2 nsew signal input
flabel locali s 18852 34885 18886 34919 0 FreeSans 400 270 0 0 Q_N
port 8 nsew signal output
flabel metal1 s 18629 33229 18663 33263 0 FreeSans 200 270 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 19173 33229 19207 33263 0 FreeSans 200 270 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 18594 28234 18690 28326 7 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 19138 28234 19234 28326 7 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 19186 28234 19186 28234 2 tapvpwrvgnd_1
flabel metal1 s 19166 28255 19204 28306 0 FreeSans 200 270 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 18633 28256 18662 28309 0 FreeSans 200 270 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 18594 26486 18690 28234 7 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 19138 26486 19234 28234 7 VGND
port 3 nsew ground bidirectional abutment
rlabel comment s 19186 26486 19186 26486 2 dfxbp_1
flabel nwell s 18642 26532 18642 26532 0 FreeSans 200 270 0 0 VPB
flabel nwell s 18625 26515 18659 26549 0 FreeSans 200 270 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 19186 26532 19186 26532 0 FreeSans 200 270 0 0 VNB
flabel pwell s 19169 26515 19203 26549 0 FreeSans 200 270 0 0 VNB
port 4 nsew ground bidirectional
flabel locali s 19067 27876 19101 27910 0 FreeSans 400 270 0 0 Q
port 7 nsew signal output
flabel locali s 18931 26515 18965 26549 0 FreeSans 400 270 0 0 CLK
port 1 nsew clock input
flabel locali s 18931 26775 18965 26809 0 FreeSans 200 270 0 0 D
port 2 nsew signal input
flabel locali s 18848 28171 18882 28205 0 FreeSans 400 270 0 0 Q_N
port 8 nsew signal output
flabel metal1 s 18625 26515 18659 26549 0 FreeSans 200 270 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 19169 26515 19203 26549 0 FreeSans 200 270 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 18602 28672 18698 30420 7 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 19146 28672 19242 30420 7 VGND
port 3 nsew ground bidirectional abutment
rlabel comment s 19194 28672 19194 28672 2 dfxbp_1
flabel nwell s 18650 28718 18650 28718 0 FreeSans 200 270 0 0 VPB
flabel nwell s 18633 28701 18667 28735 0 FreeSans 200 270 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 19194 28718 19194 28718 0 FreeSans 200 270 0 0 VNB
flabel pwell s 19177 28701 19211 28735 0 FreeSans 200 270 0 0 VNB
port 4 nsew ground bidirectional
flabel locali s 19075 30062 19109 30096 0 FreeSans 400 270 0 0 Q
port 7 nsew signal output
flabel locali s 18939 28701 18973 28735 0 FreeSans 400 270 0 0 CLK
port 1 nsew clock input
flabel locali s 18939 28961 18973 28995 0 FreeSans 200 270 0 0 D
port 2 nsew signal input
flabel locali s 18856 30357 18890 30391 0 FreeSans 400 270 0 0 Q_N
port 8 nsew signal output
flabel metal1 s 18633 28701 18667 28735 0 FreeSans 200 270 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 19177 28701 19211 28735 0 FreeSans 200 270 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 18598 24240 18694 25988 7 VPWR
port 6 nsew power bidirectional abutment
rlabel metal1 s 19142 24240 19238 25988 7 VGND
port 3 nsew ground bidirectional abutment
rlabel comment s 19190 24240 19190 24240 2 dfxbp_1
flabel nwell s 18646 24286 18646 24286 0 FreeSans 200 270 0 0 VPB
flabel nwell s 18629 24269 18663 24303 0 FreeSans 200 270 0 0 VPB
port 5 nsew power bidirectional
flabel pwell s 19190 24286 19190 24286 0 FreeSans 200 270 0 0 VNB
flabel pwell s 19173 24269 19207 24303 0 FreeSans 200 270 0 0 VNB
port 4 nsew ground bidirectional
flabel locali s 19071 25630 19105 25664 0 FreeSans 400 270 0 0 Q
port 7 nsew signal output
flabel locali s 18935 24269 18969 24303 0 FreeSans 400 270 0 0 CLK
port 1 nsew clock input
flabel locali s 18935 24529 18969 24563 0 FreeSans 200 270 0 0 D
port 2 nsew signal input
flabel locali s 18852 25925 18886 25959 0 FreeSans 400 270 0 0 Q_N
port 8 nsew signal output
flabel metal1 s 18629 24269 18663 24303 0 FreeSans 200 270 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel metal1 s 19173 24269 19207 24303 0 FreeSans 200 270 0 0 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 18598 25988 18694 26080 7 VPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 19142 25988 19238 26080 7 VGND
port 1 nsew ground bidirectional abutment
rlabel comment s 19190 25988 19190 25988 2 tapvpwrvgnd_1
flabel metal1 s 19170 26009 19208 26060 0 FreeSans 200 270 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 18637 26010 18666 26063 0 FreeSans 200 270 0 0 VPWR
port 2 nsew power bidirectional abutment
<< properties >>
string MASKHINTS_NSDM 1716 1782 1808 2009 3786 1778 3878 2005 1746 5042 1838 5269 3880 5034 3972 5261 5994 2834 6086 3061 5742 1778 5834 2005 7740 1784 7832 2011 5830 5034 5922 5261 6378 6094 6470 6321 7832 5040 7924 5267 9696 1784 9788 2011 11684 1784 11776 2011 12228 4544 12320 4771 11518 4588 11610 4815 9928 5462 10020 5689 11988 5450 12080 5677 13638 1784 13730 2011 15700 1784 15792 2011 14228 4538 14320 4765 16252 4520 16344 4747 13946 5458 14038 5685 15942 5464 16034 5691 19130 4890 19222 5117 4486 14013 4578 14240 4378 13089 4470 13316 4478 12345 4570 12572 4388 11525 4480 11752 4486 10781 4578 11008 9352 10785 9444 11012 9244 13093 9336 13320 9342 12349 9434 12576 9254 11529 9346 11756 9350 14017 9442 14244 8274 13985 8366 14212 7250 13627 7342 13854 5732 14001 5824 14228 5856 13159 5948 13386 5852 12139 5944 12366 12118 13631 12210 13858 13140 13989 13232 14216 10598 14005 10690 14232 10722 13163 10814 13390 10718 12143 10810 12370 4376 16321 4468 16548 4476 15577 4568 15804 4386 14757 4478 14984 6210 14967 6302 15194 7252 15467 7344 15694 9252 14761 9344 14988 9342 15581 9434 15808 9242 16325 9334 16552 9690 17288 9782 17515 12118 15471 12210 15698 11076 14971 11168 15198 16246 16429 16338 16656 16267 17178 16359 17405 17133 17180 17225 17407 17378 16419 17470 16646 17886 16421 17978 16648 18864 16419 18956 16646 19634 16409 19726 16636 20500 16411 20592 16638 17911 17170 18003 17397 19027 17172 19119 17399 20663 17164 20755 17391 19893 17174 19985 17401 21616 16413 21708 16640 22394 16403 22486 16630 23260 16405 23352 16632 22149 17164 22241 17391 21641 17162 21733 17389 23281 17154 23373 17381 25416 14567 25508 14794 9418 23107 9510 23334 11664 23111 11756 23338 16096 23107 16188 23334 13850 23103 13942 23330 18684 25988 18911 26080 18378 23107 18470 23334 18680 28234 18907 28326 18688 30420 18915 30512 18684 32666 18911 32758 18684 34948 18911 35040 18652 37220 18879 37312 18660 36336 18887 36428 18640 38374 18867 38466 18626 39636 18853 39728 18618 41432 18845 41524 18634 43418 18861 43510
string MASKHINTS_PSDM 1716 2093 1808 2250 3786 2089 3878 2246 1746 5353 1838 5510 3880 5345 3972 5502 5994 3145 6086 3302 5742 2089 5834 2246 7740 2095 7832 2252 5830 5345 5922 5502 6378 6405 6470 6562 7832 5351 7924 5508 9696 2095 9788 2252 11684 2095 11776 2252 12228 4855 12320 5012 11518 4899 11610 5056 9928 5773 10020 5930 11988 5761 12080 5918 13638 2095 13730 2252 15700 2095 15792 2252 14228 4849 14320 5006 16252 4831 16344 4988 13946 5769 14038 5926 15942 5775 16034 5932 19130 5201 19222 5358 4486 13772 4578 13929 4378 12848 4470 13005 4478 12104 4570 12261 4388 11284 4480 11441 4486 10540 4578 10697 9352 10544 9444 10701 9244 12852 9336 13009 9342 12108 9434 12265 9254 11288 9346 11445 9350 13776 9442 13933 8274 13744 8366 13901 7250 13386 7342 13543 5732 13760 5824 13917 5856 12918 5948 13075 5852 11898 5944 12055 12118 13390 12210 13547 13140 13748 13232 13905 10598 13764 10690 13921 10722 12922 10814 13079 10718 11902 10810 12059 4376 16080 4468 16237 4476 15336 4568 15493 4386 14516 4478 14673 6210 14726 6302 14883 7252 15226 7344 15383 9252 14520 9344 14677 9342 15340 9434 15497 9242 16084 9334 16241 9690 17599 9782 17756 12118 15230 12210 15387 11076 14730 11168 14887 16246 16188 16338 16345 16267 17489 16359 17646 17133 17491 17225 17648 17378 16178 17470 16335 17886 16180 17978 16337 18864 16178 18956 16335 19634 16168 19726 16325 20500 16170 20592 16327 17911 17481 18003 17638 19027 17483 19119 17640 20663 17475 20755 17632 19893 17485 19985 17642 21616 16172 21708 16329 22394 16162 22486 16319 23260 16164 23352 16321 22149 17475 22241 17632 21641 17473 21733 17630 23281 17465 23373 17622 25416 14326 25508 14483 9418 22866 9510 23023 11664 22870 11756 23027 16096 22866 16188 23023 13850 22862 13942 23019 18995 25988 19152 26080 18378 22866 18470 23023 18991 28234 19148 28326 18999 30420 19156 30512 18995 32666 19152 32758 18995 34948 19152 35040 18963 37220 19120 37312 18971 36336 19128 36428 18951 38374 19108 38466 18937 39636 19094 39728 18929 41432 19086 41524 18945 43418 19102 43510
<< end >>
